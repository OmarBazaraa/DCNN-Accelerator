//
// Verilog description for cell main, 
// Wed May  2 09:48:26 2018
//
// LeonardoSpectrum Level 3, 2017a.2 
//


module main ( CLK, RST, Start, FilterSize, Stride, Instr, Done ) ;

    input CLK ;
    input RST ;
    input Start ;
    input FilterSize ;
    input Stride ;
    input Instr ;
    output Done ;

    wire FirstCycle, MemWR, MemAddr_17, MemAddr_16, MemAddr_15, MemAddr_14, 
         MemAddr_13, MemAddr_12, MemAddr_11, MemAddr_10, MemAddr_9, MemAddr_8, 
         MemAddr_7, MemAddr_6, MemAddr_5, MemAddr_4, MemAddr_3, MemAddr_2, 
         MemAddr_1, MemAddr_0, MemDin_7, MemDin_6, MemDin_5, MemDin_4, MemDin_3, 
         MemDin_2, MemDin_1, MemDin_0, MemDout_39, MemDout_38, MemDout_37, 
         MemDout_36, MemDout_35, MemDout_34, MemDout_33, MemDout_32, MemDout_31, 
         MemDout_30, MemDout_29, MemDout_28, MemDout_27, MemDout_26, MemDout_25, 
         MemDout_24, MemDout_23, MemDout_22, MemDout_21, MemDout_20, MemDout_19, 
         MemDout_18, MemDout_17, MemDout_16, MemDout_15, MemDout_14, MemDout_13, 
         MemDout_12, MemDout_11, MemDout_10, MemDout_9, MemDout_8, MemDout_7, 
         MemDout_6, MemDout_5, MemDout_4, MemDout_3, MemDout_2, MemDout_1, 
         MemDout_0, CacheRST, CacheFilterWR, CacheWindowWR, CacheFilter_0__0__7, 
         CacheFilter_0__0__6, CacheFilter_0__0__5, CacheFilter_0__0__4, 
         CacheFilter_0__0__3, CacheFilter_0__0__2, CacheFilter_0__0__1, 
         CacheFilter_0__0__0, CacheFilter_0__1__7, CacheFilter_0__1__6, 
         CacheFilter_0__1__5, CacheFilter_0__1__4, CacheFilter_0__1__3, 
         CacheFilter_0__1__2, CacheFilter_0__1__1, CacheFilter_0__1__0, 
         CacheFilter_0__2__7, CacheFilter_0__2__6, CacheFilter_0__2__5, 
         CacheFilter_0__2__4, CacheFilter_0__2__3, CacheFilter_0__2__2, 
         CacheFilter_0__2__1, CacheFilter_0__2__0, CacheFilter_0__3__7, 
         CacheFilter_0__3__6, CacheFilter_0__3__5, CacheFilter_0__3__4, 
         CacheFilter_0__3__3, CacheFilter_0__3__2, CacheFilter_0__3__1, 
         CacheFilter_0__3__0, CacheFilter_0__4__7, CacheFilter_0__4__6, 
         CacheFilter_0__4__5, CacheFilter_0__4__4, CacheFilter_0__4__3, 
         CacheFilter_0__4__2, CacheFilter_0__4__1, CacheFilter_0__4__0, 
         CacheFilter_1__0__7, CacheFilter_1__0__6, CacheFilter_1__0__5, 
         CacheFilter_1__0__4, CacheFilter_1__0__3, CacheFilter_1__0__2, 
         CacheFilter_1__0__1, CacheFilter_1__0__0, CacheFilter_1__1__7, 
         CacheFilter_1__1__6, CacheFilter_1__1__5, CacheFilter_1__1__4, 
         CacheFilter_1__1__3, CacheFilter_1__1__2, CacheFilter_1__1__1, 
         CacheFilter_1__1__0, CacheFilter_1__2__7, CacheFilter_1__2__6, 
         CacheFilter_1__2__5, CacheFilter_1__2__4, CacheFilter_1__2__3, 
         CacheFilter_1__2__2, CacheFilter_1__2__1, CacheFilter_1__2__0, 
         CacheFilter_1__3__7, CacheFilter_1__3__6, CacheFilter_1__3__5, 
         CacheFilter_1__3__4, CacheFilter_1__3__3, CacheFilter_1__3__2, 
         CacheFilter_1__3__1, CacheFilter_1__3__0, CacheFilter_1__4__7, 
         CacheFilter_1__4__6, CacheFilter_1__4__5, CacheFilter_1__4__4, 
         CacheFilter_1__4__3, CacheFilter_1__4__2, CacheFilter_1__4__1, 
         CacheFilter_1__4__0, CacheFilter_2__0__7, CacheFilter_2__0__6, 
         CacheFilter_2__0__5, CacheFilter_2__0__4, CacheFilter_2__0__3, 
         CacheFilter_2__0__2, CacheFilter_2__0__1, CacheFilter_2__0__0, 
         CacheFilter_2__1__7, CacheFilter_2__1__6, CacheFilter_2__1__5, 
         CacheFilter_2__1__4, CacheFilter_2__1__3, CacheFilter_2__1__2, 
         CacheFilter_2__1__1, CacheFilter_2__1__0, CacheFilter_2__2__7, 
         CacheFilter_2__2__6, CacheFilter_2__2__5, CacheFilter_2__2__4, 
         CacheFilter_2__2__3, CacheFilter_2__2__2, CacheFilter_2__2__1, 
         CacheFilter_2__2__0, CacheFilter_2__3__7, CacheFilter_2__3__6, 
         CacheFilter_2__3__5, CacheFilter_2__3__4, CacheFilter_2__3__3, 
         CacheFilter_2__3__2, CacheFilter_2__3__1, CacheFilter_2__3__0, 
         CacheFilter_2__4__7, CacheFilter_2__4__6, CacheFilter_2__4__5, 
         CacheFilter_2__4__4, CacheFilter_2__4__3, CacheFilter_2__4__2, 
         CacheFilter_2__4__1, CacheFilter_2__4__0, CacheFilter_3__0__7, 
         CacheFilter_3__0__6, CacheFilter_3__0__5, CacheFilter_3__0__4, 
         CacheFilter_3__0__3, CacheFilter_3__0__2, CacheFilter_3__0__1, 
         CacheFilter_3__0__0, CacheFilter_3__1__7, CacheFilter_3__1__6, 
         CacheFilter_3__1__5, CacheFilter_3__1__4, CacheFilter_3__1__3, 
         CacheFilter_3__1__2, CacheFilter_3__1__1, CacheFilter_3__1__0, 
         CacheFilter_3__2__7, CacheFilter_3__2__6, CacheFilter_3__2__5, 
         CacheFilter_3__2__4, CacheFilter_3__2__3, CacheFilter_3__2__2, 
         CacheFilter_3__2__1, CacheFilter_3__2__0, CacheFilter_3__3__7, 
         CacheFilter_3__3__6, CacheFilter_3__3__5, CacheFilter_3__3__4, 
         CacheFilter_3__3__3, CacheFilter_3__3__2, CacheFilter_3__3__1, 
         CacheFilter_3__3__0, CacheFilter_3__4__7, CacheFilter_3__4__6, 
         CacheFilter_3__4__5, CacheFilter_3__4__4, CacheFilter_3__4__3, 
         CacheFilter_3__4__2, CacheFilter_3__4__1, CacheFilter_3__4__0, 
         CacheFilter_4__0__7, CacheFilter_4__0__6, CacheFilter_4__0__5, 
         CacheFilter_4__0__4, CacheFilter_4__0__3, CacheFilter_4__0__2, 
         CacheFilter_4__0__1, CacheFilter_4__0__0, CacheFilter_4__1__7, 
         CacheFilter_4__1__6, CacheFilter_4__1__5, CacheFilter_4__1__4, 
         CacheFilter_4__1__3, CacheFilter_4__1__2, CacheFilter_4__1__1, 
         CacheFilter_4__1__0, CacheFilter_4__2__7, CacheFilter_4__2__6, 
         CacheFilter_4__2__5, CacheFilter_4__2__4, CacheFilter_4__2__3, 
         CacheFilter_4__2__2, CacheFilter_4__2__1, CacheFilter_4__2__0, 
         CacheFilter_4__3__7, CacheFilter_4__3__6, CacheFilter_4__3__5, 
         CacheFilter_4__3__4, CacheFilter_4__3__3, CacheFilter_4__3__2, 
         CacheFilter_4__3__1, CacheFilter_4__3__0, CacheFilter_4__4__7, 
         CacheFilter_4__4__6, CacheFilter_4__4__5, CacheFilter_4__4__4, 
         CacheFilter_4__4__3, CacheFilter_4__4__2, CacheFilter_4__4__1, 
         CacheFilter_4__4__0, CacheWindow_0__0__7, CacheWindow_0__0__6, 
         CacheWindow_0__0__5, CacheWindow_0__0__4, CacheWindow_0__0__3, 
         CacheWindow_0__0__2, CacheWindow_0__0__1, CacheWindow_0__0__0, 
         CacheWindow_0__1__7, CacheWindow_0__1__6, CacheWindow_0__1__5, 
         CacheWindow_0__1__4, CacheWindow_0__1__3, CacheWindow_0__1__2, 
         CacheWindow_0__1__1, CacheWindow_0__1__0, CacheWindow_0__2__7, 
         CacheWindow_0__2__6, CacheWindow_0__2__5, CacheWindow_0__2__4, 
         CacheWindow_0__2__3, CacheWindow_0__2__2, CacheWindow_0__2__1, 
         CacheWindow_0__2__0, CacheWindow_0__3__7, CacheWindow_0__3__6, 
         CacheWindow_0__3__5, CacheWindow_0__3__4, CacheWindow_0__3__3, 
         CacheWindow_0__3__2, CacheWindow_0__3__1, CacheWindow_0__3__0, 
         CacheWindow_0__4__7, CacheWindow_0__4__6, CacheWindow_0__4__5, 
         CacheWindow_0__4__4, CacheWindow_0__4__3, CacheWindow_0__4__2, 
         CacheWindow_0__4__1, CacheWindow_0__4__0, CacheWindow_1__0__7, 
         CacheWindow_1__0__6, CacheWindow_1__0__5, CacheWindow_1__0__4, 
         CacheWindow_1__0__3, CacheWindow_1__0__2, CacheWindow_1__0__1, 
         CacheWindow_1__0__0, CacheWindow_1__1__7, CacheWindow_1__1__6, 
         CacheWindow_1__1__5, CacheWindow_1__1__4, CacheWindow_1__1__3, 
         CacheWindow_1__1__2, CacheWindow_1__1__1, CacheWindow_1__1__0, 
         CacheWindow_1__2__7, CacheWindow_1__2__6, CacheWindow_1__2__5, 
         CacheWindow_1__2__4, CacheWindow_1__2__3, CacheWindow_1__2__2, 
         CacheWindow_1__2__1, CacheWindow_1__2__0, CacheWindow_1__3__7, 
         CacheWindow_1__3__6, CacheWindow_1__3__5, CacheWindow_1__3__4, 
         CacheWindow_1__3__3, CacheWindow_1__3__2, CacheWindow_1__3__1, 
         CacheWindow_1__3__0, CacheWindow_1__4__7, CacheWindow_1__4__6, 
         CacheWindow_1__4__5, CacheWindow_1__4__4, CacheWindow_1__4__3, 
         CacheWindow_1__4__2, CacheWindow_1__4__1, CacheWindow_1__4__0, 
         CacheWindow_2__0__7, CacheWindow_2__0__6, CacheWindow_2__0__5, 
         CacheWindow_2__0__4, CacheWindow_2__0__3, CacheWindow_2__0__2, 
         CacheWindow_2__0__1, CacheWindow_2__0__0, CacheWindow_2__1__7, 
         CacheWindow_2__1__6, CacheWindow_2__1__5, CacheWindow_2__1__4, 
         CacheWindow_2__1__3, CacheWindow_2__1__2, CacheWindow_2__1__1, 
         CacheWindow_2__1__0, CacheWindow_2__2__7, CacheWindow_2__2__6, 
         CacheWindow_2__2__5, CacheWindow_2__2__4, CacheWindow_2__2__3, 
         CacheWindow_2__2__2, CacheWindow_2__2__1, CacheWindow_2__2__0, 
         CacheWindow_2__3__7, CacheWindow_2__3__6, CacheWindow_2__3__5, 
         CacheWindow_2__3__4, CacheWindow_2__3__3, CacheWindow_2__3__2, 
         CacheWindow_2__3__1, CacheWindow_2__3__0, CacheWindow_2__4__7, 
         CacheWindow_2__4__6, CacheWindow_2__4__5, CacheWindow_2__4__4, 
         CacheWindow_2__4__3, CacheWindow_2__4__2, CacheWindow_2__4__1, 
         CacheWindow_2__4__0, CacheWindow_3__0__7, CacheWindow_3__0__6, 
         CacheWindow_3__0__5, CacheWindow_3__0__4, CacheWindow_3__0__3, 
         CacheWindow_3__0__2, CacheWindow_3__0__1, CacheWindow_3__0__0, 
         CacheWindow_3__1__7, CacheWindow_3__1__6, CacheWindow_3__1__5, 
         CacheWindow_3__1__4, CacheWindow_3__1__3, CacheWindow_3__1__2, 
         CacheWindow_3__1__1, CacheWindow_3__1__0, CacheWindow_3__2__7, 
         CacheWindow_3__2__6, CacheWindow_3__2__5, CacheWindow_3__2__4, 
         CacheWindow_3__2__3, CacheWindow_3__2__2, CacheWindow_3__2__1, 
         CacheWindow_3__2__0, CacheWindow_3__3__7, CacheWindow_3__3__6, 
         CacheWindow_3__3__5, CacheWindow_3__3__4, CacheWindow_3__3__3, 
         CacheWindow_3__3__2, CacheWindow_3__3__1, CacheWindow_3__3__0, 
         CacheWindow_3__4__7, CacheWindow_3__4__6, CacheWindow_3__4__5, 
         CacheWindow_3__4__4, CacheWindow_3__4__3, CacheWindow_3__4__2, 
         CacheWindow_3__4__1, CacheWindow_3__4__0, CacheWindow_4__0__7, 
         CacheWindow_4__0__6, CacheWindow_4__0__5, CacheWindow_4__0__4, 
         CacheWindow_4__0__3, CacheWindow_4__0__2, CacheWindow_4__0__1, 
         CacheWindow_4__0__0, CacheWindow_4__1__7, CacheWindow_4__1__6, 
         CacheWindow_4__1__5, CacheWindow_4__1__4, CacheWindow_4__1__3, 
         CacheWindow_4__1__2, CacheWindow_4__1__1, CacheWindow_4__1__0, 
         CacheWindow_4__2__7, CacheWindow_4__2__6, CacheWindow_4__2__5, 
         CacheWindow_4__2__4, CacheWindow_4__2__3, CacheWindow_4__2__2, 
         CacheWindow_4__2__1, CacheWindow_4__2__0, CacheWindow_4__3__7, 
         CacheWindow_4__3__6, CacheWindow_4__3__5, CacheWindow_4__3__4, 
         CacheWindow_4__3__3, CacheWindow_4__3__2, CacheWindow_4__3__1, 
         CacheWindow_4__3__0, CacheWindow_4__4__7, CacheWindow_4__4__6, 
         CacheWindow_4__4__5, CacheWindow_4__4__4, CacheWindow_4__4__3, 
         CacheWindow_4__4__2, CacheWindow_4__4__1, CacheWindow_4__4__0, 
         AccStartCalc, AccFinishCalc, AccResult_7, AccResult_6, AccResult_5, 
         AccResult_4, AccResult_3, AccResult_2, AccResult_1, AccResult_0, GND0;
    wire [0:0] \$dummy ;




    controller CONTROLLER (.CLK (CLK), .RST (RST), .Start (Start), .FilterSize (
               FilterSize), .Stride (Stride), .Instr (Instr), .CalcFinished (
               AccFinishCalc), .Calc (AccStartCalc), .MemRD (\$dummy [0]), .MemWR (
               MemWR), .MemAddr ({MemAddr_17,MemAddr_16,MemAddr_15,MemAddr_14,
               MemAddr_13,MemAddr_12,MemAddr_11,MemAddr_10,MemAddr_9,MemAddr_8,
               MemAddr_7,MemAddr_6,MemAddr_5,MemAddr_4,MemAddr_3,MemAddr_2,
               MemAddr_1,MemAddr_0}), .CacheFilterWR (CacheFilterWR), .CacheWindowWR (
               CacheWindowWR), .FirstCycle (FirstCycle), .Done (Done)) ;
    accelerator ACCELERATOR (.CLK (CLK), .RST (RST), .Start (AccStartCalc), .FilterSize (
                FilterSize), .Instr (Instr), .FilterDin_0__0__7 (
                CacheFilter_0__0__7), .FilterDin_0__0__6 (CacheFilter_0__0__6), 
                .FilterDin_0__0__5 (CacheFilter_0__0__5), .FilterDin_0__0__4 (
                CacheFilter_0__0__4), .FilterDin_0__0__3 (CacheFilter_0__0__3), 
                .FilterDin_0__0__2 (CacheFilter_0__0__2), .FilterDin_0__0__1 (
                CacheFilter_0__0__1), .FilterDin_0__0__0 (CacheFilter_0__0__0), 
                .FilterDin_0__1__7 (CacheFilter_0__1__7), .FilterDin_0__1__6 (
                CacheFilter_0__1__6), .FilterDin_0__1__5 (CacheFilter_0__1__5), 
                .FilterDin_0__1__4 (CacheFilter_0__1__4), .FilterDin_0__1__3 (
                CacheFilter_0__1__3), .FilterDin_0__1__2 (CacheFilter_0__1__2), 
                .FilterDin_0__1__1 (CacheFilter_0__1__1), .FilterDin_0__1__0 (
                CacheFilter_0__1__0), .FilterDin_0__2__7 (CacheFilter_0__2__7), 
                .FilterDin_0__2__6 (CacheFilter_0__2__6), .FilterDin_0__2__5 (
                CacheFilter_0__2__5), .FilterDin_0__2__4 (CacheFilter_0__2__4), 
                .FilterDin_0__2__3 (CacheFilter_0__2__3), .FilterDin_0__2__2 (
                CacheFilter_0__2__2), .FilterDin_0__2__1 (CacheFilter_0__2__1), 
                .FilterDin_0__2__0 (CacheFilter_0__2__0), .FilterDin_0__3__7 (
                CacheFilter_0__3__7), .FilterDin_0__3__6 (CacheFilter_0__3__6), 
                .FilterDin_0__3__5 (CacheFilter_0__3__5), .FilterDin_0__3__4 (
                CacheFilter_0__3__4), .FilterDin_0__3__3 (CacheFilter_0__3__3), 
                .FilterDin_0__3__2 (CacheFilter_0__3__2), .FilterDin_0__3__1 (
                CacheFilter_0__3__1), .FilterDin_0__3__0 (CacheFilter_0__3__0), 
                .FilterDin_0__4__7 (CacheFilter_0__4__7), .FilterDin_0__4__6 (
                CacheFilter_0__4__6), .FilterDin_0__4__5 (CacheFilter_0__4__5), 
                .FilterDin_0__4__4 (CacheFilter_0__4__4), .FilterDin_0__4__3 (
                CacheFilter_0__4__3), .FilterDin_0__4__2 (CacheFilter_0__4__2), 
                .FilterDin_0__4__1 (CacheFilter_0__4__1), .FilterDin_0__4__0 (
                CacheFilter_0__4__0), .FilterDin_1__0__7 (CacheFilter_1__0__7), 
                .FilterDin_1__0__6 (CacheFilter_1__0__6), .FilterDin_1__0__5 (
                CacheFilter_1__0__5), .FilterDin_1__0__4 (CacheFilter_1__0__4), 
                .FilterDin_1__0__3 (CacheFilter_1__0__3), .FilterDin_1__0__2 (
                CacheFilter_1__0__2), .FilterDin_1__0__1 (CacheFilter_1__0__1), 
                .FilterDin_1__0__0 (CacheFilter_1__0__0), .FilterDin_1__1__7 (
                CacheFilter_1__1__7), .FilterDin_1__1__6 (CacheFilter_1__1__6), 
                .FilterDin_1__1__5 (CacheFilter_1__1__5), .FilterDin_1__1__4 (
                CacheFilter_1__1__4), .FilterDin_1__1__3 (CacheFilter_1__1__3), 
                .FilterDin_1__1__2 (CacheFilter_1__1__2), .FilterDin_1__1__1 (
                CacheFilter_1__1__1), .FilterDin_1__1__0 (CacheFilter_1__1__0), 
                .FilterDin_1__2__7 (CacheFilter_1__2__7), .FilterDin_1__2__6 (
                CacheFilter_1__2__6), .FilterDin_1__2__5 (CacheFilter_1__2__5), 
                .FilterDin_1__2__4 (CacheFilter_1__2__4), .FilterDin_1__2__3 (
                CacheFilter_1__2__3), .FilterDin_1__2__2 (CacheFilter_1__2__2), 
                .FilterDin_1__2__1 (CacheFilter_1__2__1), .FilterDin_1__2__0 (
                CacheFilter_1__2__0), .FilterDin_1__3__7 (CacheFilter_1__3__7), 
                .FilterDin_1__3__6 (CacheFilter_1__3__6), .FilterDin_1__3__5 (
                CacheFilter_1__3__5), .FilterDin_1__3__4 (CacheFilter_1__3__4), 
                .FilterDin_1__3__3 (CacheFilter_1__3__3), .FilterDin_1__3__2 (
                CacheFilter_1__3__2), .FilterDin_1__3__1 (CacheFilter_1__3__1), 
                .FilterDin_1__3__0 (CacheFilter_1__3__0), .FilterDin_1__4__7 (
                CacheFilter_1__4__7), .FilterDin_1__4__6 (CacheFilter_1__4__6), 
                .FilterDin_1__4__5 (CacheFilter_1__4__5), .FilterDin_1__4__4 (
                CacheFilter_1__4__4), .FilterDin_1__4__3 (CacheFilter_1__4__3), 
                .FilterDin_1__4__2 (CacheFilter_1__4__2), .FilterDin_1__4__1 (
                CacheFilter_1__4__1), .FilterDin_1__4__0 (CacheFilter_1__4__0), 
                .FilterDin_2__0__7 (CacheFilter_2__0__7), .FilterDin_2__0__6 (
                CacheFilter_2__0__6), .FilterDin_2__0__5 (CacheFilter_2__0__5), 
                .FilterDin_2__0__4 (CacheFilter_2__0__4), .FilterDin_2__0__3 (
                CacheFilter_2__0__3), .FilterDin_2__0__2 (CacheFilter_2__0__2), 
                .FilterDin_2__0__1 (CacheFilter_2__0__1), .FilterDin_2__0__0 (
                CacheFilter_2__0__0), .FilterDin_2__1__7 (CacheFilter_2__1__7), 
                .FilterDin_2__1__6 (CacheFilter_2__1__6), .FilterDin_2__1__5 (
                CacheFilter_2__1__5), .FilterDin_2__1__4 (CacheFilter_2__1__4), 
                .FilterDin_2__1__3 (CacheFilter_2__1__3), .FilterDin_2__1__2 (
                CacheFilter_2__1__2), .FilterDin_2__1__1 (CacheFilter_2__1__1), 
                .FilterDin_2__1__0 (CacheFilter_2__1__0), .FilterDin_2__2__7 (
                CacheFilter_2__2__7), .FilterDin_2__2__6 (CacheFilter_2__2__6), 
                .FilterDin_2__2__5 (CacheFilter_2__2__5), .FilterDin_2__2__4 (
                CacheFilter_2__2__4), .FilterDin_2__2__3 (CacheFilter_2__2__3), 
                .FilterDin_2__2__2 (CacheFilter_2__2__2), .FilterDin_2__2__1 (
                CacheFilter_2__2__1), .FilterDin_2__2__0 (CacheFilter_2__2__0), 
                .FilterDin_2__3__7 (CacheFilter_2__3__7), .FilterDin_2__3__6 (
                CacheFilter_2__3__6), .FilterDin_2__3__5 (CacheFilter_2__3__5), 
                .FilterDin_2__3__4 (CacheFilter_2__3__4), .FilterDin_2__3__3 (
                CacheFilter_2__3__3), .FilterDin_2__3__2 (CacheFilter_2__3__2), 
                .FilterDin_2__3__1 (CacheFilter_2__3__1), .FilterDin_2__3__0 (
                CacheFilter_2__3__0), .FilterDin_2__4__7 (CacheFilter_2__4__7), 
                .FilterDin_2__4__6 (CacheFilter_2__4__6), .FilterDin_2__4__5 (
                CacheFilter_2__4__5), .FilterDin_2__4__4 (CacheFilter_2__4__4), 
                .FilterDin_2__4__3 (CacheFilter_2__4__3), .FilterDin_2__4__2 (
                CacheFilter_2__4__2), .FilterDin_2__4__1 (CacheFilter_2__4__1), 
                .FilterDin_2__4__0 (CacheFilter_2__4__0), .FilterDin_3__0__7 (
                CacheFilter_3__0__7), .FilterDin_3__0__6 (CacheFilter_3__0__6), 
                .FilterDin_3__0__5 (CacheFilter_3__0__5), .FilterDin_3__0__4 (
                CacheFilter_3__0__4), .FilterDin_3__0__3 (CacheFilter_3__0__3), 
                .FilterDin_3__0__2 (CacheFilter_3__0__2), .FilterDin_3__0__1 (
                CacheFilter_3__0__1), .FilterDin_3__0__0 (CacheFilter_3__0__0), 
                .FilterDin_3__1__7 (CacheFilter_3__1__7), .FilterDin_3__1__6 (
                CacheFilter_3__1__6), .FilterDin_3__1__5 (CacheFilter_3__1__5), 
                .FilterDin_3__1__4 (CacheFilter_3__1__4), .FilterDin_3__1__3 (
                CacheFilter_3__1__3), .FilterDin_3__1__2 (CacheFilter_3__1__2), 
                .FilterDin_3__1__1 (CacheFilter_3__1__1), .FilterDin_3__1__0 (
                CacheFilter_3__1__0), .FilterDin_3__2__7 (CacheFilter_3__2__7), 
                .FilterDin_3__2__6 (CacheFilter_3__2__6), .FilterDin_3__2__5 (
                CacheFilter_3__2__5), .FilterDin_3__2__4 (CacheFilter_3__2__4), 
                .FilterDin_3__2__3 (CacheFilter_3__2__3), .FilterDin_3__2__2 (
                CacheFilter_3__2__2), .FilterDin_3__2__1 (CacheFilter_3__2__1), 
                .FilterDin_3__2__0 (CacheFilter_3__2__0), .FilterDin_3__3__7 (
                CacheFilter_3__3__7), .FilterDin_3__3__6 (CacheFilter_3__3__6), 
                .FilterDin_3__3__5 (CacheFilter_3__3__5), .FilterDin_3__3__4 (
                CacheFilter_3__3__4), .FilterDin_3__3__3 (CacheFilter_3__3__3), 
                .FilterDin_3__3__2 (CacheFilter_3__3__2), .FilterDin_3__3__1 (
                CacheFilter_3__3__1), .FilterDin_3__3__0 (CacheFilter_3__3__0), 
                .FilterDin_3__4__7 (CacheFilter_3__4__7), .FilterDin_3__4__6 (
                CacheFilter_3__4__6), .FilterDin_3__4__5 (CacheFilter_3__4__5), 
                .FilterDin_3__4__4 (CacheFilter_3__4__4), .FilterDin_3__4__3 (
                CacheFilter_3__4__3), .FilterDin_3__4__2 (CacheFilter_3__4__2), 
                .FilterDin_3__4__1 (CacheFilter_3__4__1), .FilterDin_3__4__0 (
                CacheFilter_3__4__0), .FilterDin_4__0__7 (CacheFilter_4__0__7), 
                .FilterDin_4__0__6 (CacheFilter_4__0__6), .FilterDin_4__0__5 (
                CacheFilter_4__0__5), .FilterDin_4__0__4 (CacheFilter_4__0__4), 
                .FilterDin_4__0__3 (CacheFilter_4__0__3), .FilterDin_4__0__2 (
                CacheFilter_4__0__2), .FilterDin_4__0__1 (CacheFilter_4__0__1), 
                .FilterDin_4__0__0 (CacheFilter_4__0__0), .FilterDin_4__1__7 (
                CacheFilter_4__1__7), .FilterDin_4__1__6 (CacheFilter_4__1__6), 
                .FilterDin_4__1__5 (CacheFilter_4__1__5), .FilterDin_4__1__4 (
                CacheFilter_4__1__4), .FilterDin_4__1__3 (CacheFilter_4__1__3), 
                .FilterDin_4__1__2 (CacheFilter_4__1__2), .FilterDin_4__1__1 (
                CacheFilter_4__1__1), .FilterDin_4__1__0 (CacheFilter_4__1__0), 
                .FilterDin_4__2__7 (CacheFilter_4__2__7), .FilterDin_4__2__6 (
                CacheFilter_4__2__6), .FilterDin_4__2__5 (CacheFilter_4__2__5), 
                .FilterDin_4__2__4 (CacheFilter_4__2__4), .FilterDin_4__2__3 (
                CacheFilter_4__2__3), .FilterDin_4__2__2 (CacheFilter_4__2__2), 
                .FilterDin_4__2__1 (CacheFilter_4__2__1), .FilterDin_4__2__0 (
                CacheFilter_4__2__0), .FilterDin_4__3__7 (CacheFilter_4__3__7), 
                .FilterDin_4__3__6 (CacheFilter_4__3__6), .FilterDin_4__3__5 (
                CacheFilter_4__3__5), .FilterDin_4__3__4 (CacheFilter_4__3__4), 
                .FilterDin_4__3__3 (CacheFilter_4__3__3), .FilterDin_4__3__2 (
                CacheFilter_4__3__2), .FilterDin_4__3__1 (CacheFilter_4__3__1), 
                .FilterDin_4__3__0 (CacheFilter_4__3__0), .FilterDin_4__4__7 (
                CacheFilter_4__4__7), .FilterDin_4__4__6 (CacheFilter_4__4__6), 
                .FilterDin_4__4__5 (CacheFilter_4__4__5), .FilterDin_4__4__4 (
                CacheFilter_4__4__4), .FilterDin_4__4__3 (CacheFilter_4__4__3), 
                .FilterDin_4__4__2 (CacheFilter_4__4__2), .FilterDin_4__4__1 (
                CacheFilter_4__4__1), .FilterDin_4__4__0 (CacheFilter_4__4__0), 
                .WindowDin_0__0__7 (CacheWindow_0__0__7), .WindowDin_0__0__6 (
                CacheWindow_0__0__6), .WindowDin_0__0__5 (CacheWindow_0__0__5), 
                .WindowDin_0__0__4 (CacheWindow_0__0__4), .WindowDin_0__0__3 (
                CacheWindow_0__0__3), .WindowDin_0__0__2 (CacheWindow_0__0__2), 
                .WindowDin_0__0__1 (CacheWindow_0__0__1), .WindowDin_0__0__0 (
                CacheWindow_0__0__0), .WindowDin_0__1__7 (CacheWindow_0__1__7), 
                .WindowDin_0__1__6 (CacheWindow_0__1__6), .WindowDin_0__1__5 (
                CacheWindow_0__1__5), .WindowDin_0__1__4 (CacheWindow_0__1__4), 
                .WindowDin_0__1__3 (CacheWindow_0__1__3), .WindowDin_0__1__2 (
                CacheWindow_0__1__2), .WindowDin_0__1__1 (CacheWindow_0__1__1), 
                .WindowDin_0__1__0 (CacheWindow_0__1__0), .WindowDin_0__2__7 (
                CacheWindow_0__2__7), .WindowDin_0__2__6 (CacheWindow_0__2__6), 
                .WindowDin_0__2__5 (CacheWindow_0__2__5), .WindowDin_0__2__4 (
                CacheWindow_0__2__4), .WindowDin_0__2__3 (CacheWindow_0__2__3), 
                .WindowDin_0__2__2 (CacheWindow_0__2__2), .WindowDin_0__2__1 (
                CacheWindow_0__2__1), .WindowDin_0__2__0 (CacheWindow_0__2__0), 
                .WindowDin_0__3__7 (CacheWindow_0__3__7), .WindowDin_0__3__6 (
                CacheWindow_0__3__6), .WindowDin_0__3__5 (CacheWindow_0__3__5), 
                .WindowDin_0__3__4 (CacheWindow_0__3__4), .WindowDin_0__3__3 (
                CacheWindow_0__3__3), .WindowDin_0__3__2 (CacheWindow_0__3__2), 
                .WindowDin_0__3__1 (CacheWindow_0__3__1), .WindowDin_0__3__0 (
                CacheWindow_0__3__0), .WindowDin_0__4__7 (CacheWindow_0__4__7), 
                .WindowDin_0__4__6 (CacheWindow_0__4__6), .WindowDin_0__4__5 (
                CacheWindow_0__4__5), .WindowDin_0__4__4 (CacheWindow_0__4__4), 
                .WindowDin_0__4__3 (CacheWindow_0__4__3), .WindowDin_0__4__2 (
                CacheWindow_0__4__2), .WindowDin_0__4__1 (CacheWindow_0__4__1), 
                .WindowDin_0__4__0 (CacheWindow_0__4__0), .WindowDin_1__0__7 (
                CacheWindow_1__0__7), .WindowDin_1__0__6 (CacheWindow_1__0__6), 
                .WindowDin_1__0__5 (CacheWindow_1__0__5), .WindowDin_1__0__4 (
                CacheWindow_1__0__4), .WindowDin_1__0__3 (CacheWindow_1__0__3), 
                .WindowDin_1__0__2 (CacheWindow_1__0__2), .WindowDin_1__0__1 (
                CacheWindow_1__0__1), .WindowDin_1__0__0 (CacheWindow_1__0__0), 
                .WindowDin_1__1__7 (CacheWindow_1__1__7), .WindowDin_1__1__6 (
                CacheWindow_1__1__6), .WindowDin_1__1__5 (CacheWindow_1__1__5), 
                .WindowDin_1__1__4 (CacheWindow_1__1__4), .WindowDin_1__1__3 (
                CacheWindow_1__1__3), .WindowDin_1__1__2 (CacheWindow_1__1__2), 
                .WindowDin_1__1__1 (CacheWindow_1__1__1), .WindowDin_1__1__0 (
                CacheWindow_1__1__0), .WindowDin_1__2__7 (CacheWindow_1__2__7), 
                .WindowDin_1__2__6 (CacheWindow_1__2__6), .WindowDin_1__2__5 (
                CacheWindow_1__2__5), .WindowDin_1__2__4 (CacheWindow_1__2__4), 
                .WindowDin_1__2__3 (CacheWindow_1__2__3), .WindowDin_1__2__2 (
                CacheWindow_1__2__2), .WindowDin_1__2__1 (CacheWindow_1__2__1), 
                .WindowDin_1__2__0 (CacheWindow_1__2__0), .WindowDin_1__3__7 (
                CacheWindow_1__3__7), .WindowDin_1__3__6 (CacheWindow_1__3__6), 
                .WindowDin_1__3__5 (CacheWindow_1__3__5), .WindowDin_1__3__4 (
                CacheWindow_1__3__4), .WindowDin_1__3__3 (CacheWindow_1__3__3), 
                .WindowDin_1__3__2 (CacheWindow_1__3__2), .WindowDin_1__3__1 (
                CacheWindow_1__3__1), .WindowDin_1__3__0 (CacheWindow_1__3__0), 
                .WindowDin_1__4__7 (CacheWindow_1__4__7), .WindowDin_1__4__6 (
                CacheWindow_1__4__6), .WindowDin_1__4__5 (CacheWindow_1__4__5), 
                .WindowDin_1__4__4 (CacheWindow_1__4__4), .WindowDin_1__4__3 (
                CacheWindow_1__4__3), .WindowDin_1__4__2 (CacheWindow_1__4__2), 
                .WindowDin_1__4__1 (CacheWindow_1__4__1), .WindowDin_1__4__0 (
                CacheWindow_1__4__0), .WindowDin_2__0__7 (CacheWindow_2__0__7), 
                .WindowDin_2__0__6 (CacheWindow_2__0__6), .WindowDin_2__0__5 (
                CacheWindow_2__0__5), .WindowDin_2__0__4 (CacheWindow_2__0__4), 
                .WindowDin_2__0__3 (CacheWindow_2__0__3), .WindowDin_2__0__2 (
                CacheWindow_2__0__2), .WindowDin_2__0__1 (CacheWindow_2__0__1), 
                .WindowDin_2__0__0 (CacheWindow_2__0__0), .WindowDin_2__1__7 (
                CacheWindow_2__1__7), .WindowDin_2__1__6 (CacheWindow_2__1__6), 
                .WindowDin_2__1__5 (CacheWindow_2__1__5), .WindowDin_2__1__4 (
                CacheWindow_2__1__4), .WindowDin_2__1__3 (CacheWindow_2__1__3), 
                .WindowDin_2__1__2 (CacheWindow_2__1__2), .WindowDin_2__1__1 (
                CacheWindow_2__1__1), .WindowDin_2__1__0 (CacheWindow_2__1__0), 
                .WindowDin_2__2__7 (CacheWindow_2__2__7), .WindowDin_2__2__6 (
                CacheWindow_2__2__6), .WindowDin_2__2__5 (CacheWindow_2__2__5), 
                .WindowDin_2__2__4 (CacheWindow_2__2__4), .WindowDin_2__2__3 (
                CacheWindow_2__2__3), .WindowDin_2__2__2 (CacheWindow_2__2__2), 
                .WindowDin_2__2__1 (CacheWindow_2__2__1), .WindowDin_2__2__0 (
                CacheWindow_2__2__0), .WindowDin_2__3__7 (CacheWindow_2__3__7), 
                .WindowDin_2__3__6 (CacheWindow_2__3__6), .WindowDin_2__3__5 (
                CacheWindow_2__3__5), .WindowDin_2__3__4 (CacheWindow_2__3__4), 
                .WindowDin_2__3__3 (CacheWindow_2__3__3), .WindowDin_2__3__2 (
                CacheWindow_2__3__2), .WindowDin_2__3__1 (CacheWindow_2__3__1), 
                .WindowDin_2__3__0 (CacheWindow_2__3__0), .WindowDin_2__4__7 (
                CacheWindow_2__4__7), .WindowDin_2__4__6 (CacheWindow_2__4__6), 
                .WindowDin_2__4__5 (CacheWindow_2__4__5), .WindowDin_2__4__4 (
                CacheWindow_2__4__4), .WindowDin_2__4__3 (CacheWindow_2__4__3), 
                .WindowDin_2__4__2 (CacheWindow_2__4__2), .WindowDin_2__4__1 (
                CacheWindow_2__4__1), .WindowDin_2__4__0 (CacheWindow_2__4__0), 
                .WindowDin_3__0__7 (CacheWindow_3__0__7), .WindowDin_3__0__6 (
                CacheWindow_3__0__6), .WindowDin_3__0__5 (CacheWindow_3__0__5), 
                .WindowDin_3__0__4 (CacheWindow_3__0__4), .WindowDin_3__0__3 (
                CacheWindow_3__0__3), .WindowDin_3__0__2 (CacheWindow_3__0__2), 
                .WindowDin_3__0__1 (CacheWindow_3__0__1), .WindowDin_3__0__0 (
                CacheWindow_3__0__0), .WindowDin_3__1__7 (CacheWindow_3__1__7), 
                .WindowDin_3__1__6 (CacheWindow_3__1__6), .WindowDin_3__1__5 (
                CacheWindow_3__1__5), .WindowDin_3__1__4 (CacheWindow_3__1__4), 
                .WindowDin_3__1__3 (CacheWindow_3__1__3), .WindowDin_3__1__2 (
                CacheWindow_3__1__2), .WindowDin_3__1__1 (CacheWindow_3__1__1), 
                .WindowDin_3__1__0 (CacheWindow_3__1__0), .WindowDin_3__2__7 (
                CacheWindow_3__2__7), .WindowDin_3__2__6 (CacheWindow_3__2__6), 
                .WindowDin_3__2__5 (CacheWindow_3__2__5), .WindowDin_3__2__4 (
                CacheWindow_3__2__4), .WindowDin_3__2__3 (CacheWindow_3__2__3), 
                .WindowDin_3__2__2 (CacheWindow_3__2__2), .WindowDin_3__2__1 (
                CacheWindow_3__2__1), .WindowDin_3__2__0 (CacheWindow_3__2__0), 
                .WindowDin_3__3__7 (CacheWindow_3__3__7), .WindowDin_3__3__6 (
                CacheWindow_3__3__6), .WindowDin_3__3__5 (CacheWindow_3__3__5), 
                .WindowDin_3__3__4 (CacheWindow_3__3__4), .WindowDin_3__3__3 (
                CacheWindow_3__3__3), .WindowDin_3__3__2 (CacheWindow_3__3__2), 
                .WindowDin_3__3__1 (CacheWindow_3__3__1), .WindowDin_3__3__0 (
                CacheWindow_3__3__0), .WindowDin_3__4__7 (CacheWindow_3__4__7), 
                .WindowDin_3__4__6 (CacheWindow_3__4__6), .WindowDin_3__4__5 (
                CacheWindow_3__4__5), .WindowDin_3__4__4 (CacheWindow_3__4__4), 
                .WindowDin_3__4__3 (CacheWindow_3__4__3), .WindowDin_3__4__2 (
                CacheWindow_3__4__2), .WindowDin_3__4__1 (CacheWindow_3__4__1), 
                .WindowDin_3__4__0 (CacheWindow_3__4__0), .WindowDin_4__0__7 (
                CacheWindow_4__0__7), .WindowDin_4__0__6 (CacheWindow_4__0__6), 
                .WindowDin_4__0__5 (CacheWindow_4__0__5), .WindowDin_4__0__4 (
                CacheWindow_4__0__4), .WindowDin_4__0__3 (CacheWindow_4__0__3), 
                .WindowDin_4__0__2 (CacheWindow_4__0__2), .WindowDin_4__0__1 (
                CacheWindow_4__0__1), .WindowDin_4__0__0 (CacheWindow_4__0__0), 
                .WindowDin_4__1__7 (CacheWindow_4__1__7), .WindowDin_4__1__6 (
                CacheWindow_4__1__6), .WindowDin_4__1__5 (CacheWindow_4__1__5), 
                .WindowDin_4__1__4 (CacheWindow_4__1__4), .WindowDin_4__1__3 (
                CacheWindow_4__1__3), .WindowDin_4__1__2 (CacheWindow_4__1__2), 
                .WindowDin_4__1__1 (CacheWindow_4__1__1), .WindowDin_4__1__0 (
                CacheWindow_4__1__0), .WindowDin_4__2__7 (CacheWindow_4__2__7), 
                .WindowDin_4__2__6 (CacheWindow_4__2__6), .WindowDin_4__2__5 (
                CacheWindow_4__2__5), .WindowDin_4__2__4 (CacheWindow_4__2__4), 
                .WindowDin_4__2__3 (CacheWindow_4__2__3), .WindowDin_4__2__2 (
                CacheWindow_4__2__2), .WindowDin_4__2__1 (CacheWindow_4__2__1), 
                .WindowDin_4__2__0 (CacheWindow_4__2__0), .WindowDin_4__3__7 (
                CacheWindow_4__3__7), .WindowDin_4__3__6 (CacheWindow_4__3__6), 
                .WindowDin_4__3__5 (CacheWindow_4__3__5), .WindowDin_4__3__4 (
                CacheWindow_4__3__4), .WindowDin_4__3__3 (CacheWindow_4__3__3), 
                .WindowDin_4__3__2 (CacheWindow_4__3__2), .WindowDin_4__3__1 (
                CacheWindow_4__3__1), .WindowDin_4__3__0 (CacheWindow_4__3__0), 
                .WindowDin_4__4__7 (CacheWindow_4__4__7), .WindowDin_4__4__6 (
                CacheWindow_4__4__6), .WindowDin_4__4__5 (CacheWindow_4__4__5), 
                .WindowDin_4__4__4 (CacheWindow_4__4__4), .WindowDin_4__4__3 (
                CacheWindow_4__4__3), .WindowDin_4__4__2 (CacheWindow_4__4__2), 
                .WindowDin_4__4__1 (CacheWindow_4__4__1), .WindowDin_4__4__0 (
                CacheWindow_4__4__0), .Done (AccFinishCalc), .Result ({
                AccResult_7,AccResult_6,AccResult_5,AccResult_4,AccResult_3,
                AccResult_2,AccResult_1,AccResult_0})) ;
    RAM_8_18 RAM (.CLK (CLK), .WR (MemWR), .Address ({MemAddr_17,MemAddr_16,
             MemAddr_15,MemAddr_14,MemAddr_13,MemAddr_12,MemAddr_11,MemAddr_10,
             MemAddr_9,MemAddr_8,MemAddr_7,MemAddr_6,MemAddr_5,MemAddr_4,
             MemAddr_3,MemAddr_2,MemAddr_1,MemAddr_0}), .Din ({MemDin_7,MemDin_6
             ,MemDin_5,MemDin_4,MemDin_3,MemDin_2,MemDin_1,MemDin_0}), .Dout ({
             MemDout_39,MemDout_38,MemDout_37,MemDout_36,MemDout_35,MemDout_34,
             MemDout_33,MemDout_32,MemDout_31,MemDout_30,MemDout_29,MemDout_28,
             MemDout_27,MemDout_26,MemDout_25,MemDout_24,MemDout_23,MemDout_22,
             MemDout_21,MemDout_20,MemDout_19,MemDout_18,MemDout_17,MemDout_16,
             MemDout_15,MemDout_14,MemDout_13,MemDout_12,MemDout_11,MemDout_10,
             MemDout_9,MemDout_8,MemDout_7,MemDout_6,MemDout_5,MemDout_4,
             MemDout_3,MemDout_2,MemDout_1,MemDout_0})) ;
    or (CacheRST, RST, FirstCycle) ;
    cache CACHE (.CLK (CLK), .RST (CacheRST), .FilterSize (FilterSize), .FilterWR (
          CacheFilterWR), .WindowWR (CacheWindowWR), .Din ({MemDout_39,
          MemDout_38,MemDout_37,MemDout_36,MemDout_35,MemDout_34,MemDout_33,
          MemDout_32,MemDout_31,MemDout_30,MemDout_29,MemDout_28,MemDout_27,
          MemDout_26,MemDout_25,MemDout_24,MemDout_23,MemDout_22,MemDout_21,
          MemDout_20,MemDout_19,MemDout_18,MemDout_17,MemDout_16,MemDout_15,
          MemDout_14,MemDout_13,MemDout_12,MemDout_11,MemDout_10,MemDout_9,
          MemDout_8,MemDout_7,MemDout_6,MemDout_5,MemDout_4,MemDout_3,MemDout_2,
          MemDout_1,MemDout_0}), .FilterDout_0__0__7 (CacheFilter_0__0__7), .FilterDout_0__0__6 (
          CacheFilter_0__0__6), .FilterDout_0__0__5 (CacheFilter_0__0__5), .FilterDout_0__0__4 (
          CacheFilter_0__0__4), .FilterDout_0__0__3 (CacheFilter_0__0__3), .FilterDout_0__0__2 (
          CacheFilter_0__0__2), .FilterDout_0__0__1 (CacheFilter_0__0__1), .FilterDout_0__0__0 (
          CacheFilter_0__0__0), .FilterDout_0__1__7 (CacheFilter_0__1__7), .FilterDout_0__1__6 (
          CacheFilter_0__1__6), .FilterDout_0__1__5 (CacheFilter_0__1__5), .FilterDout_0__1__4 (
          CacheFilter_0__1__4), .FilterDout_0__1__3 (CacheFilter_0__1__3), .FilterDout_0__1__2 (
          CacheFilter_0__1__2), .FilterDout_0__1__1 (CacheFilter_0__1__1), .FilterDout_0__1__0 (
          CacheFilter_0__1__0), .FilterDout_0__2__7 (CacheFilter_0__2__7), .FilterDout_0__2__6 (
          CacheFilter_0__2__6), .FilterDout_0__2__5 (CacheFilter_0__2__5), .FilterDout_0__2__4 (
          CacheFilter_0__2__4), .FilterDout_0__2__3 (CacheFilter_0__2__3), .FilterDout_0__2__2 (
          CacheFilter_0__2__2), .FilterDout_0__2__1 (CacheFilter_0__2__1), .FilterDout_0__2__0 (
          CacheFilter_0__2__0), .FilterDout_0__3__7 (CacheFilter_0__3__7), .FilterDout_0__3__6 (
          CacheFilter_0__3__6), .FilterDout_0__3__5 (CacheFilter_0__3__5), .FilterDout_0__3__4 (
          CacheFilter_0__3__4), .FilterDout_0__3__3 (CacheFilter_0__3__3), .FilterDout_0__3__2 (
          CacheFilter_0__3__2), .FilterDout_0__3__1 (CacheFilter_0__3__1), .FilterDout_0__3__0 (
          CacheFilter_0__3__0), .FilterDout_0__4__7 (CacheFilter_0__4__7), .FilterDout_0__4__6 (
          CacheFilter_0__4__6), .FilterDout_0__4__5 (CacheFilter_0__4__5), .FilterDout_0__4__4 (
          CacheFilter_0__4__4), .FilterDout_0__4__3 (CacheFilter_0__4__3), .FilterDout_0__4__2 (
          CacheFilter_0__4__2), .FilterDout_0__4__1 (CacheFilter_0__4__1), .FilterDout_0__4__0 (
          CacheFilter_0__4__0), .FilterDout_1__0__7 (CacheFilter_1__0__7), .FilterDout_1__0__6 (
          CacheFilter_1__0__6), .FilterDout_1__0__5 (CacheFilter_1__0__5), .FilterDout_1__0__4 (
          CacheFilter_1__0__4), .FilterDout_1__0__3 (CacheFilter_1__0__3), .FilterDout_1__0__2 (
          CacheFilter_1__0__2), .FilterDout_1__0__1 (CacheFilter_1__0__1), .FilterDout_1__0__0 (
          CacheFilter_1__0__0), .FilterDout_1__1__7 (CacheFilter_1__1__7), .FilterDout_1__1__6 (
          CacheFilter_1__1__6), .FilterDout_1__1__5 (CacheFilter_1__1__5), .FilterDout_1__1__4 (
          CacheFilter_1__1__4), .FilterDout_1__1__3 (CacheFilter_1__1__3), .FilterDout_1__1__2 (
          CacheFilter_1__1__2), .FilterDout_1__1__1 (CacheFilter_1__1__1), .FilterDout_1__1__0 (
          CacheFilter_1__1__0), .FilterDout_1__2__7 (CacheFilter_1__2__7), .FilterDout_1__2__6 (
          CacheFilter_1__2__6), .FilterDout_1__2__5 (CacheFilter_1__2__5), .FilterDout_1__2__4 (
          CacheFilter_1__2__4), .FilterDout_1__2__3 (CacheFilter_1__2__3), .FilterDout_1__2__2 (
          CacheFilter_1__2__2), .FilterDout_1__2__1 (CacheFilter_1__2__1), .FilterDout_1__2__0 (
          CacheFilter_1__2__0), .FilterDout_1__3__7 (CacheFilter_1__3__7), .FilterDout_1__3__6 (
          CacheFilter_1__3__6), .FilterDout_1__3__5 (CacheFilter_1__3__5), .FilterDout_1__3__4 (
          CacheFilter_1__3__4), .FilterDout_1__3__3 (CacheFilter_1__3__3), .FilterDout_1__3__2 (
          CacheFilter_1__3__2), .FilterDout_1__3__1 (CacheFilter_1__3__1), .FilterDout_1__3__0 (
          CacheFilter_1__3__0), .FilterDout_1__4__7 (CacheFilter_1__4__7), .FilterDout_1__4__6 (
          CacheFilter_1__4__6), .FilterDout_1__4__5 (CacheFilter_1__4__5), .FilterDout_1__4__4 (
          CacheFilter_1__4__4), .FilterDout_1__4__3 (CacheFilter_1__4__3), .FilterDout_1__4__2 (
          CacheFilter_1__4__2), .FilterDout_1__4__1 (CacheFilter_1__4__1), .FilterDout_1__4__0 (
          CacheFilter_1__4__0), .FilterDout_2__0__7 (CacheFilter_2__0__7), .FilterDout_2__0__6 (
          CacheFilter_2__0__6), .FilterDout_2__0__5 (CacheFilter_2__0__5), .FilterDout_2__0__4 (
          CacheFilter_2__0__4), .FilterDout_2__0__3 (CacheFilter_2__0__3), .FilterDout_2__0__2 (
          CacheFilter_2__0__2), .FilterDout_2__0__1 (CacheFilter_2__0__1), .FilterDout_2__0__0 (
          CacheFilter_2__0__0), .FilterDout_2__1__7 (CacheFilter_2__1__7), .FilterDout_2__1__6 (
          CacheFilter_2__1__6), .FilterDout_2__1__5 (CacheFilter_2__1__5), .FilterDout_2__1__4 (
          CacheFilter_2__1__4), .FilterDout_2__1__3 (CacheFilter_2__1__3), .FilterDout_2__1__2 (
          CacheFilter_2__1__2), .FilterDout_2__1__1 (CacheFilter_2__1__1), .FilterDout_2__1__0 (
          CacheFilter_2__1__0), .FilterDout_2__2__7 (CacheFilter_2__2__7), .FilterDout_2__2__6 (
          CacheFilter_2__2__6), .FilterDout_2__2__5 (CacheFilter_2__2__5), .FilterDout_2__2__4 (
          CacheFilter_2__2__4), .FilterDout_2__2__3 (CacheFilter_2__2__3), .FilterDout_2__2__2 (
          CacheFilter_2__2__2), .FilterDout_2__2__1 (CacheFilter_2__2__1), .FilterDout_2__2__0 (
          CacheFilter_2__2__0), .FilterDout_2__3__7 (CacheFilter_2__3__7), .FilterDout_2__3__6 (
          CacheFilter_2__3__6), .FilterDout_2__3__5 (CacheFilter_2__3__5), .FilterDout_2__3__4 (
          CacheFilter_2__3__4), .FilterDout_2__3__3 (CacheFilter_2__3__3), .FilterDout_2__3__2 (
          CacheFilter_2__3__2), .FilterDout_2__3__1 (CacheFilter_2__3__1), .FilterDout_2__3__0 (
          CacheFilter_2__3__0), .FilterDout_2__4__7 (CacheFilter_2__4__7), .FilterDout_2__4__6 (
          CacheFilter_2__4__6), .FilterDout_2__4__5 (CacheFilter_2__4__5), .FilterDout_2__4__4 (
          CacheFilter_2__4__4), .FilterDout_2__4__3 (CacheFilter_2__4__3), .FilterDout_2__4__2 (
          CacheFilter_2__4__2), .FilterDout_2__4__1 (CacheFilter_2__4__1), .FilterDout_2__4__0 (
          CacheFilter_2__4__0), .FilterDout_3__0__7 (CacheFilter_3__0__7), .FilterDout_3__0__6 (
          CacheFilter_3__0__6), .FilterDout_3__0__5 (CacheFilter_3__0__5), .FilterDout_3__0__4 (
          CacheFilter_3__0__4), .FilterDout_3__0__3 (CacheFilter_3__0__3), .FilterDout_3__0__2 (
          CacheFilter_3__0__2), .FilterDout_3__0__1 (CacheFilter_3__0__1), .FilterDout_3__0__0 (
          CacheFilter_3__0__0), .FilterDout_3__1__7 (CacheFilter_3__1__7), .FilterDout_3__1__6 (
          CacheFilter_3__1__6), .FilterDout_3__1__5 (CacheFilter_3__1__5), .FilterDout_3__1__4 (
          CacheFilter_3__1__4), .FilterDout_3__1__3 (CacheFilter_3__1__3), .FilterDout_3__1__2 (
          CacheFilter_3__1__2), .FilterDout_3__1__1 (CacheFilter_3__1__1), .FilterDout_3__1__0 (
          CacheFilter_3__1__0), .FilterDout_3__2__7 (CacheFilter_3__2__7), .FilterDout_3__2__6 (
          CacheFilter_3__2__6), .FilterDout_3__2__5 (CacheFilter_3__2__5), .FilterDout_3__2__4 (
          CacheFilter_3__2__4), .FilterDout_3__2__3 (CacheFilter_3__2__3), .FilterDout_3__2__2 (
          CacheFilter_3__2__2), .FilterDout_3__2__1 (CacheFilter_3__2__1), .FilterDout_3__2__0 (
          CacheFilter_3__2__0), .FilterDout_3__3__7 (CacheFilter_3__3__7), .FilterDout_3__3__6 (
          CacheFilter_3__3__6), .FilterDout_3__3__5 (CacheFilter_3__3__5), .FilterDout_3__3__4 (
          CacheFilter_3__3__4), .FilterDout_3__3__3 (CacheFilter_3__3__3), .FilterDout_3__3__2 (
          CacheFilter_3__3__2), .FilterDout_3__3__1 (CacheFilter_3__3__1), .FilterDout_3__3__0 (
          CacheFilter_3__3__0), .FilterDout_3__4__7 (CacheFilter_3__4__7), .FilterDout_3__4__6 (
          CacheFilter_3__4__6), .FilterDout_3__4__5 (CacheFilter_3__4__5), .FilterDout_3__4__4 (
          CacheFilter_3__4__4), .FilterDout_3__4__3 (CacheFilter_3__4__3), .FilterDout_3__4__2 (
          CacheFilter_3__4__2), .FilterDout_3__4__1 (CacheFilter_3__4__1), .FilterDout_3__4__0 (
          CacheFilter_3__4__0), .FilterDout_4__0__7 (CacheFilter_4__0__7), .FilterDout_4__0__6 (
          CacheFilter_4__0__6), .FilterDout_4__0__5 (CacheFilter_4__0__5), .FilterDout_4__0__4 (
          CacheFilter_4__0__4), .FilterDout_4__0__3 (CacheFilter_4__0__3), .FilterDout_4__0__2 (
          CacheFilter_4__0__2), .FilterDout_4__0__1 (CacheFilter_4__0__1), .FilterDout_4__0__0 (
          CacheFilter_4__0__0), .FilterDout_4__1__7 (CacheFilter_4__1__7), .FilterDout_4__1__6 (
          CacheFilter_4__1__6), .FilterDout_4__1__5 (CacheFilter_4__1__5), .FilterDout_4__1__4 (
          CacheFilter_4__1__4), .FilterDout_4__1__3 (CacheFilter_4__1__3), .FilterDout_4__1__2 (
          CacheFilter_4__1__2), .FilterDout_4__1__1 (CacheFilter_4__1__1), .FilterDout_4__1__0 (
          CacheFilter_4__1__0), .FilterDout_4__2__7 (CacheFilter_4__2__7), .FilterDout_4__2__6 (
          CacheFilter_4__2__6), .FilterDout_4__2__5 (CacheFilter_4__2__5), .FilterDout_4__2__4 (
          CacheFilter_4__2__4), .FilterDout_4__2__3 (CacheFilter_4__2__3), .FilterDout_4__2__2 (
          CacheFilter_4__2__2), .FilterDout_4__2__1 (CacheFilter_4__2__1), .FilterDout_4__2__0 (
          CacheFilter_4__2__0), .FilterDout_4__3__7 (CacheFilter_4__3__7), .FilterDout_4__3__6 (
          CacheFilter_4__3__6), .FilterDout_4__3__5 (CacheFilter_4__3__5), .FilterDout_4__3__4 (
          CacheFilter_4__3__4), .FilterDout_4__3__3 (CacheFilter_4__3__3), .FilterDout_4__3__2 (
          CacheFilter_4__3__2), .FilterDout_4__3__1 (CacheFilter_4__3__1), .FilterDout_4__3__0 (
          CacheFilter_4__3__0), .FilterDout_4__4__7 (CacheFilter_4__4__7), .FilterDout_4__4__6 (
          CacheFilter_4__4__6), .FilterDout_4__4__5 (CacheFilter_4__4__5), .FilterDout_4__4__4 (
          CacheFilter_4__4__4), .FilterDout_4__4__3 (CacheFilter_4__4__3), .FilterDout_4__4__2 (
          CacheFilter_4__4__2), .FilterDout_4__4__1 (CacheFilter_4__4__1), .FilterDout_4__4__0 (
          CacheFilter_4__4__0), .WindowDout_0__0__7 (CacheWindow_0__0__7), .WindowDout_0__0__6 (
          CacheWindow_0__0__6), .WindowDout_0__0__5 (CacheWindow_0__0__5), .WindowDout_0__0__4 (
          CacheWindow_0__0__4), .WindowDout_0__0__3 (CacheWindow_0__0__3), .WindowDout_0__0__2 (
          CacheWindow_0__0__2), .WindowDout_0__0__1 (CacheWindow_0__0__1), .WindowDout_0__0__0 (
          CacheWindow_0__0__0), .WindowDout_0__1__7 (CacheWindow_0__1__7), .WindowDout_0__1__6 (
          CacheWindow_0__1__6), .WindowDout_0__1__5 (CacheWindow_0__1__5), .WindowDout_0__1__4 (
          CacheWindow_0__1__4), .WindowDout_0__1__3 (CacheWindow_0__1__3), .WindowDout_0__1__2 (
          CacheWindow_0__1__2), .WindowDout_0__1__1 (CacheWindow_0__1__1), .WindowDout_0__1__0 (
          CacheWindow_0__1__0), .WindowDout_0__2__7 (CacheWindow_0__2__7), .WindowDout_0__2__6 (
          CacheWindow_0__2__6), .WindowDout_0__2__5 (CacheWindow_0__2__5), .WindowDout_0__2__4 (
          CacheWindow_0__2__4), .WindowDout_0__2__3 (CacheWindow_0__2__3), .WindowDout_0__2__2 (
          CacheWindow_0__2__2), .WindowDout_0__2__1 (CacheWindow_0__2__1), .WindowDout_0__2__0 (
          CacheWindow_0__2__0), .WindowDout_0__3__7 (CacheWindow_0__3__7), .WindowDout_0__3__6 (
          CacheWindow_0__3__6), .WindowDout_0__3__5 (CacheWindow_0__3__5), .WindowDout_0__3__4 (
          CacheWindow_0__3__4), .WindowDout_0__3__3 (CacheWindow_0__3__3), .WindowDout_0__3__2 (
          CacheWindow_0__3__2), .WindowDout_0__3__1 (CacheWindow_0__3__1), .WindowDout_0__3__0 (
          CacheWindow_0__3__0), .WindowDout_0__4__7 (CacheWindow_0__4__7), .WindowDout_0__4__6 (
          CacheWindow_0__4__6), .WindowDout_0__4__5 (CacheWindow_0__4__5), .WindowDout_0__4__4 (
          CacheWindow_0__4__4), .WindowDout_0__4__3 (CacheWindow_0__4__3), .WindowDout_0__4__2 (
          CacheWindow_0__4__2), .WindowDout_0__4__1 (CacheWindow_0__4__1), .WindowDout_0__4__0 (
          CacheWindow_0__4__0), .WindowDout_1__0__7 (CacheWindow_1__0__7), .WindowDout_1__0__6 (
          CacheWindow_1__0__6), .WindowDout_1__0__5 (CacheWindow_1__0__5), .WindowDout_1__0__4 (
          CacheWindow_1__0__4), .WindowDout_1__0__3 (CacheWindow_1__0__3), .WindowDout_1__0__2 (
          CacheWindow_1__0__2), .WindowDout_1__0__1 (CacheWindow_1__0__1), .WindowDout_1__0__0 (
          CacheWindow_1__0__0), .WindowDout_1__1__7 (CacheWindow_1__1__7), .WindowDout_1__1__6 (
          CacheWindow_1__1__6), .WindowDout_1__1__5 (CacheWindow_1__1__5), .WindowDout_1__1__4 (
          CacheWindow_1__1__4), .WindowDout_1__1__3 (CacheWindow_1__1__3), .WindowDout_1__1__2 (
          CacheWindow_1__1__2), .WindowDout_1__1__1 (CacheWindow_1__1__1), .WindowDout_1__1__0 (
          CacheWindow_1__1__0), .WindowDout_1__2__7 (CacheWindow_1__2__7), .WindowDout_1__2__6 (
          CacheWindow_1__2__6), .WindowDout_1__2__5 (CacheWindow_1__2__5), .WindowDout_1__2__4 (
          CacheWindow_1__2__4), .WindowDout_1__2__3 (CacheWindow_1__2__3), .WindowDout_1__2__2 (
          CacheWindow_1__2__2), .WindowDout_1__2__1 (CacheWindow_1__2__1), .WindowDout_1__2__0 (
          CacheWindow_1__2__0), .WindowDout_1__3__7 (CacheWindow_1__3__7), .WindowDout_1__3__6 (
          CacheWindow_1__3__6), .WindowDout_1__3__5 (CacheWindow_1__3__5), .WindowDout_1__3__4 (
          CacheWindow_1__3__4), .WindowDout_1__3__3 (CacheWindow_1__3__3), .WindowDout_1__3__2 (
          CacheWindow_1__3__2), .WindowDout_1__3__1 (CacheWindow_1__3__1), .WindowDout_1__3__0 (
          CacheWindow_1__3__0), .WindowDout_1__4__7 (CacheWindow_1__4__7), .WindowDout_1__4__6 (
          CacheWindow_1__4__6), .WindowDout_1__4__5 (CacheWindow_1__4__5), .WindowDout_1__4__4 (
          CacheWindow_1__4__4), .WindowDout_1__4__3 (CacheWindow_1__4__3), .WindowDout_1__4__2 (
          CacheWindow_1__4__2), .WindowDout_1__4__1 (CacheWindow_1__4__1), .WindowDout_1__4__0 (
          CacheWindow_1__4__0), .WindowDout_2__0__7 (CacheWindow_2__0__7), .WindowDout_2__0__6 (
          CacheWindow_2__0__6), .WindowDout_2__0__5 (CacheWindow_2__0__5), .WindowDout_2__0__4 (
          CacheWindow_2__0__4), .WindowDout_2__0__3 (CacheWindow_2__0__3), .WindowDout_2__0__2 (
          CacheWindow_2__0__2), .WindowDout_2__0__1 (CacheWindow_2__0__1), .WindowDout_2__0__0 (
          CacheWindow_2__0__0), .WindowDout_2__1__7 (CacheWindow_2__1__7), .WindowDout_2__1__6 (
          CacheWindow_2__1__6), .WindowDout_2__1__5 (CacheWindow_2__1__5), .WindowDout_2__1__4 (
          CacheWindow_2__1__4), .WindowDout_2__1__3 (CacheWindow_2__1__3), .WindowDout_2__1__2 (
          CacheWindow_2__1__2), .WindowDout_2__1__1 (CacheWindow_2__1__1), .WindowDout_2__1__0 (
          CacheWindow_2__1__0), .WindowDout_2__2__7 (CacheWindow_2__2__7), .WindowDout_2__2__6 (
          CacheWindow_2__2__6), .WindowDout_2__2__5 (CacheWindow_2__2__5), .WindowDout_2__2__4 (
          CacheWindow_2__2__4), .WindowDout_2__2__3 (CacheWindow_2__2__3), .WindowDout_2__2__2 (
          CacheWindow_2__2__2), .WindowDout_2__2__1 (CacheWindow_2__2__1), .WindowDout_2__2__0 (
          CacheWindow_2__2__0), .WindowDout_2__3__7 (CacheWindow_2__3__7), .WindowDout_2__3__6 (
          CacheWindow_2__3__6), .WindowDout_2__3__5 (CacheWindow_2__3__5), .WindowDout_2__3__4 (
          CacheWindow_2__3__4), .WindowDout_2__3__3 (CacheWindow_2__3__3), .WindowDout_2__3__2 (
          CacheWindow_2__3__2), .WindowDout_2__3__1 (CacheWindow_2__3__1), .WindowDout_2__3__0 (
          CacheWindow_2__3__0), .WindowDout_2__4__7 (CacheWindow_2__4__7), .WindowDout_2__4__6 (
          CacheWindow_2__4__6), .WindowDout_2__4__5 (CacheWindow_2__4__5), .WindowDout_2__4__4 (
          CacheWindow_2__4__4), .WindowDout_2__4__3 (CacheWindow_2__4__3), .WindowDout_2__4__2 (
          CacheWindow_2__4__2), .WindowDout_2__4__1 (CacheWindow_2__4__1), .WindowDout_2__4__0 (
          CacheWindow_2__4__0), .WindowDout_3__0__7 (CacheWindow_3__0__7), .WindowDout_3__0__6 (
          CacheWindow_3__0__6), .WindowDout_3__0__5 (CacheWindow_3__0__5), .WindowDout_3__0__4 (
          CacheWindow_3__0__4), .WindowDout_3__0__3 (CacheWindow_3__0__3), .WindowDout_3__0__2 (
          CacheWindow_3__0__2), .WindowDout_3__0__1 (CacheWindow_3__0__1), .WindowDout_3__0__0 (
          CacheWindow_3__0__0), .WindowDout_3__1__7 (CacheWindow_3__1__7), .WindowDout_3__1__6 (
          CacheWindow_3__1__6), .WindowDout_3__1__5 (CacheWindow_3__1__5), .WindowDout_3__1__4 (
          CacheWindow_3__1__4), .WindowDout_3__1__3 (CacheWindow_3__1__3), .WindowDout_3__1__2 (
          CacheWindow_3__1__2), .WindowDout_3__1__1 (CacheWindow_3__1__1), .WindowDout_3__1__0 (
          CacheWindow_3__1__0), .WindowDout_3__2__7 (CacheWindow_3__2__7), .WindowDout_3__2__6 (
          CacheWindow_3__2__6), .WindowDout_3__2__5 (CacheWindow_3__2__5), .WindowDout_3__2__4 (
          CacheWindow_3__2__4), .WindowDout_3__2__3 (CacheWindow_3__2__3), .WindowDout_3__2__2 (
          CacheWindow_3__2__2), .WindowDout_3__2__1 (CacheWindow_3__2__1), .WindowDout_3__2__0 (
          CacheWindow_3__2__0), .WindowDout_3__3__7 (CacheWindow_3__3__7), .WindowDout_3__3__6 (
          CacheWindow_3__3__6), .WindowDout_3__3__5 (CacheWindow_3__3__5), .WindowDout_3__3__4 (
          CacheWindow_3__3__4), .WindowDout_3__3__3 (CacheWindow_3__3__3), .WindowDout_3__3__2 (
          CacheWindow_3__3__2), .WindowDout_3__3__1 (CacheWindow_3__3__1), .WindowDout_3__3__0 (
          CacheWindow_3__3__0), .WindowDout_3__4__7 (CacheWindow_3__4__7), .WindowDout_3__4__6 (
          CacheWindow_3__4__6), .WindowDout_3__4__5 (CacheWindow_3__4__5), .WindowDout_3__4__4 (
          CacheWindow_3__4__4), .WindowDout_3__4__3 (CacheWindow_3__4__3), .WindowDout_3__4__2 (
          CacheWindow_3__4__2), .WindowDout_3__4__1 (CacheWindow_3__4__1), .WindowDout_3__4__0 (
          CacheWindow_3__4__0), .WindowDout_4__0__7 (CacheWindow_4__0__7), .WindowDout_4__0__6 (
          CacheWindow_4__0__6), .WindowDout_4__0__5 (CacheWindow_4__0__5), .WindowDout_4__0__4 (
          CacheWindow_4__0__4), .WindowDout_4__0__3 (CacheWindow_4__0__3), .WindowDout_4__0__2 (
          CacheWindow_4__0__2), .WindowDout_4__0__1 (CacheWindow_4__0__1), .WindowDout_4__0__0 (
          CacheWindow_4__0__0), .WindowDout_4__1__7 (CacheWindow_4__1__7), .WindowDout_4__1__6 (
          CacheWindow_4__1__6), .WindowDout_4__1__5 (CacheWindow_4__1__5), .WindowDout_4__1__4 (
          CacheWindow_4__1__4), .WindowDout_4__1__3 (CacheWindow_4__1__3), .WindowDout_4__1__2 (
          CacheWindow_4__1__2), .WindowDout_4__1__1 (CacheWindow_4__1__1), .WindowDout_4__1__0 (
          CacheWindow_4__1__0), .WindowDout_4__2__7 (CacheWindow_4__2__7), .WindowDout_4__2__6 (
          CacheWindow_4__2__6), .WindowDout_4__2__5 (CacheWindow_4__2__5), .WindowDout_4__2__4 (
          CacheWindow_4__2__4), .WindowDout_4__2__3 (CacheWindow_4__2__3), .WindowDout_4__2__2 (
          CacheWindow_4__2__2), .WindowDout_4__2__1 (CacheWindow_4__2__1), .WindowDout_4__2__0 (
          CacheWindow_4__2__0), .WindowDout_4__3__7 (CacheWindow_4__3__7), .WindowDout_4__3__6 (
          CacheWindow_4__3__6), .WindowDout_4__3__5 (CacheWindow_4__3__5), .WindowDout_4__3__4 (
          CacheWindow_4__3__4), .WindowDout_4__3__3 (CacheWindow_4__3__3), .WindowDout_4__3__2 (
          CacheWindow_4__3__2), .WindowDout_4__3__1 (CacheWindow_4__3__1), .WindowDout_4__3__0 (
          CacheWindow_4__3__0), .WindowDout_4__4__7 (CacheWindow_4__4__7), .WindowDout_4__4__6 (
          CacheWindow_4__4__6), .WindowDout_4__4__5 (CacheWindow_4__4__5), .WindowDout_4__4__4 (
          CacheWindow_4__4__4), .WindowDout_4__4__3 (CacheWindow_4__4__3), .WindowDout_4__4__2 (
          CacheWindow_4__4__2), .WindowDout_4__4__1 (CacheWindow_4__4__1), .WindowDout_4__4__0 (
          CacheWindow_4__4__0), .ResultWR (GND0), .ResultDin ({AccResult_7,
          AccResult_6,AccResult_5,AccResult_4,AccResult_3,AccResult_2,
          AccResult_1,AccResult_0}), .ResultDout ({MemDin_7,MemDin_6,MemDin_5,
          MemDin_4,MemDin_3,MemDin_2,MemDin_1,MemDin_0})) ;
    assign GND0 = 0 ;
endmodule


module cache ( CLK, RST, FilterSize, FilterWR, WindowWR, Din, FilterDout_0__0__7, 
               FilterDout_0__0__6, FilterDout_0__0__5, FilterDout_0__0__4, 
               FilterDout_0__0__3, FilterDout_0__0__2, FilterDout_0__0__1, 
               FilterDout_0__0__0, FilterDout_0__1__7, FilterDout_0__1__6, 
               FilterDout_0__1__5, FilterDout_0__1__4, FilterDout_0__1__3, 
               FilterDout_0__1__2, FilterDout_0__1__1, FilterDout_0__1__0, 
               FilterDout_0__2__7, FilterDout_0__2__6, FilterDout_0__2__5, 
               FilterDout_0__2__4, FilterDout_0__2__3, FilterDout_0__2__2, 
               FilterDout_0__2__1, FilterDout_0__2__0, FilterDout_0__3__7, 
               FilterDout_0__3__6, FilterDout_0__3__5, FilterDout_0__3__4, 
               FilterDout_0__3__3, FilterDout_0__3__2, FilterDout_0__3__1, 
               FilterDout_0__3__0, FilterDout_0__4__7, FilterDout_0__4__6, 
               FilterDout_0__4__5, FilterDout_0__4__4, FilterDout_0__4__3, 
               FilterDout_0__4__2, FilterDout_0__4__1, FilterDout_0__4__0, 
               FilterDout_1__0__7, FilterDout_1__0__6, FilterDout_1__0__5, 
               FilterDout_1__0__4, FilterDout_1__0__3, FilterDout_1__0__2, 
               FilterDout_1__0__1, FilterDout_1__0__0, FilterDout_1__1__7, 
               FilterDout_1__1__6, FilterDout_1__1__5, FilterDout_1__1__4, 
               FilterDout_1__1__3, FilterDout_1__1__2, FilterDout_1__1__1, 
               FilterDout_1__1__0, FilterDout_1__2__7, FilterDout_1__2__6, 
               FilterDout_1__2__5, FilterDout_1__2__4, FilterDout_1__2__3, 
               FilterDout_1__2__2, FilterDout_1__2__1, FilterDout_1__2__0, 
               FilterDout_1__3__7, FilterDout_1__3__6, FilterDout_1__3__5, 
               FilterDout_1__3__4, FilterDout_1__3__3, FilterDout_1__3__2, 
               FilterDout_1__3__1, FilterDout_1__3__0, FilterDout_1__4__7, 
               FilterDout_1__4__6, FilterDout_1__4__5, FilterDout_1__4__4, 
               FilterDout_1__4__3, FilterDout_1__4__2, FilterDout_1__4__1, 
               FilterDout_1__4__0, FilterDout_2__0__7, FilterDout_2__0__6, 
               FilterDout_2__0__5, FilterDout_2__0__4, FilterDout_2__0__3, 
               FilterDout_2__0__2, FilterDout_2__0__1, FilterDout_2__0__0, 
               FilterDout_2__1__7, FilterDout_2__1__6, FilterDout_2__1__5, 
               FilterDout_2__1__4, FilterDout_2__1__3, FilterDout_2__1__2, 
               FilterDout_2__1__1, FilterDout_2__1__0, FilterDout_2__2__7, 
               FilterDout_2__2__6, FilterDout_2__2__5, FilterDout_2__2__4, 
               FilterDout_2__2__3, FilterDout_2__2__2, FilterDout_2__2__1, 
               FilterDout_2__2__0, FilterDout_2__3__7, FilterDout_2__3__6, 
               FilterDout_2__3__5, FilterDout_2__3__4, FilterDout_2__3__3, 
               FilterDout_2__3__2, FilterDout_2__3__1, FilterDout_2__3__0, 
               FilterDout_2__4__7, FilterDout_2__4__6, FilterDout_2__4__5, 
               FilterDout_2__4__4, FilterDout_2__4__3, FilterDout_2__4__2, 
               FilterDout_2__4__1, FilterDout_2__4__0, FilterDout_3__0__7, 
               FilterDout_3__0__6, FilterDout_3__0__5, FilterDout_3__0__4, 
               FilterDout_3__0__3, FilterDout_3__0__2, FilterDout_3__0__1, 
               FilterDout_3__0__0, FilterDout_3__1__7, FilterDout_3__1__6, 
               FilterDout_3__1__5, FilterDout_3__1__4, FilterDout_3__1__3, 
               FilterDout_3__1__2, FilterDout_3__1__1, FilterDout_3__1__0, 
               FilterDout_3__2__7, FilterDout_3__2__6, FilterDout_3__2__5, 
               FilterDout_3__2__4, FilterDout_3__2__3, FilterDout_3__2__2, 
               FilterDout_3__2__1, FilterDout_3__2__0, FilterDout_3__3__7, 
               FilterDout_3__3__6, FilterDout_3__3__5, FilterDout_3__3__4, 
               FilterDout_3__3__3, FilterDout_3__3__2, FilterDout_3__3__1, 
               FilterDout_3__3__0, FilterDout_3__4__7, FilterDout_3__4__6, 
               FilterDout_3__4__5, FilterDout_3__4__4, FilterDout_3__4__3, 
               FilterDout_3__4__2, FilterDout_3__4__1, FilterDout_3__4__0, 
               FilterDout_4__0__7, FilterDout_4__0__6, FilterDout_4__0__5, 
               FilterDout_4__0__4, FilterDout_4__0__3, FilterDout_4__0__2, 
               FilterDout_4__0__1, FilterDout_4__0__0, FilterDout_4__1__7, 
               FilterDout_4__1__6, FilterDout_4__1__5, FilterDout_4__1__4, 
               FilterDout_4__1__3, FilterDout_4__1__2, FilterDout_4__1__1, 
               FilterDout_4__1__0, FilterDout_4__2__7, FilterDout_4__2__6, 
               FilterDout_4__2__5, FilterDout_4__2__4, FilterDout_4__2__3, 
               FilterDout_4__2__2, FilterDout_4__2__1, FilterDout_4__2__0, 
               FilterDout_4__3__7, FilterDout_4__3__6, FilterDout_4__3__5, 
               FilterDout_4__3__4, FilterDout_4__3__3, FilterDout_4__3__2, 
               FilterDout_4__3__1, FilterDout_4__3__0, FilterDout_4__4__7, 
               FilterDout_4__4__6, FilterDout_4__4__5, FilterDout_4__4__4, 
               FilterDout_4__4__3, FilterDout_4__4__2, FilterDout_4__4__1, 
               FilterDout_4__4__0, WindowDout_0__0__7, WindowDout_0__0__6, 
               WindowDout_0__0__5, WindowDout_0__0__4, WindowDout_0__0__3, 
               WindowDout_0__0__2, WindowDout_0__0__1, WindowDout_0__0__0, 
               WindowDout_0__1__7, WindowDout_0__1__6, WindowDout_0__1__5, 
               WindowDout_0__1__4, WindowDout_0__1__3, WindowDout_0__1__2, 
               WindowDout_0__1__1, WindowDout_0__1__0, WindowDout_0__2__7, 
               WindowDout_0__2__6, WindowDout_0__2__5, WindowDout_0__2__4, 
               WindowDout_0__2__3, WindowDout_0__2__2, WindowDout_0__2__1, 
               WindowDout_0__2__0, WindowDout_0__3__7, WindowDout_0__3__6, 
               WindowDout_0__3__5, WindowDout_0__3__4, WindowDout_0__3__3, 
               WindowDout_0__3__2, WindowDout_0__3__1, WindowDout_0__3__0, 
               WindowDout_0__4__7, WindowDout_0__4__6, WindowDout_0__4__5, 
               WindowDout_0__4__4, WindowDout_0__4__3, WindowDout_0__4__2, 
               WindowDout_0__4__1, WindowDout_0__4__0, WindowDout_1__0__7, 
               WindowDout_1__0__6, WindowDout_1__0__5, WindowDout_1__0__4, 
               WindowDout_1__0__3, WindowDout_1__0__2, WindowDout_1__0__1, 
               WindowDout_1__0__0, WindowDout_1__1__7, WindowDout_1__1__6, 
               WindowDout_1__1__5, WindowDout_1__1__4, WindowDout_1__1__3, 
               WindowDout_1__1__2, WindowDout_1__1__1, WindowDout_1__1__0, 
               WindowDout_1__2__7, WindowDout_1__2__6, WindowDout_1__2__5, 
               WindowDout_1__2__4, WindowDout_1__2__3, WindowDout_1__2__2, 
               WindowDout_1__2__1, WindowDout_1__2__0, WindowDout_1__3__7, 
               WindowDout_1__3__6, WindowDout_1__3__5, WindowDout_1__3__4, 
               WindowDout_1__3__3, WindowDout_1__3__2, WindowDout_1__3__1, 
               WindowDout_1__3__0, WindowDout_1__4__7, WindowDout_1__4__6, 
               WindowDout_1__4__5, WindowDout_1__4__4, WindowDout_1__4__3, 
               WindowDout_1__4__2, WindowDout_1__4__1, WindowDout_1__4__0, 
               WindowDout_2__0__7, WindowDout_2__0__6, WindowDout_2__0__5, 
               WindowDout_2__0__4, WindowDout_2__0__3, WindowDout_2__0__2, 
               WindowDout_2__0__1, WindowDout_2__0__0, WindowDout_2__1__7, 
               WindowDout_2__1__6, WindowDout_2__1__5, WindowDout_2__1__4, 
               WindowDout_2__1__3, WindowDout_2__1__2, WindowDout_2__1__1, 
               WindowDout_2__1__0, WindowDout_2__2__7, WindowDout_2__2__6, 
               WindowDout_2__2__5, WindowDout_2__2__4, WindowDout_2__2__3, 
               WindowDout_2__2__2, WindowDout_2__2__1, WindowDout_2__2__0, 
               WindowDout_2__3__7, WindowDout_2__3__6, WindowDout_2__3__5, 
               WindowDout_2__3__4, WindowDout_2__3__3, WindowDout_2__3__2, 
               WindowDout_2__3__1, WindowDout_2__3__0, WindowDout_2__4__7, 
               WindowDout_2__4__6, WindowDout_2__4__5, WindowDout_2__4__4, 
               WindowDout_2__4__3, WindowDout_2__4__2, WindowDout_2__4__1, 
               WindowDout_2__4__0, WindowDout_3__0__7, WindowDout_3__0__6, 
               WindowDout_3__0__5, WindowDout_3__0__4, WindowDout_3__0__3, 
               WindowDout_3__0__2, WindowDout_3__0__1, WindowDout_3__0__0, 
               WindowDout_3__1__7, WindowDout_3__1__6, WindowDout_3__1__5, 
               WindowDout_3__1__4, WindowDout_3__1__3, WindowDout_3__1__2, 
               WindowDout_3__1__1, WindowDout_3__1__0, WindowDout_3__2__7, 
               WindowDout_3__2__6, WindowDout_3__2__5, WindowDout_3__2__4, 
               WindowDout_3__2__3, WindowDout_3__2__2, WindowDout_3__2__1, 
               WindowDout_3__2__0, WindowDout_3__3__7, WindowDout_3__3__6, 
               WindowDout_3__3__5, WindowDout_3__3__4, WindowDout_3__3__3, 
               WindowDout_3__3__2, WindowDout_3__3__1, WindowDout_3__3__0, 
               WindowDout_3__4__7, WindowDout_3__4__6, WindowDout_3__4__5, 
               WindowDout_3__4__4, WindowDout_3__4__3, WindowDout_3__4__2, 
               WindowDout_3__4__1, WindowDout_3__4__0, WindowDout_4__0__7, 
               WindowDout_4__0__6, WindowDout_4__0__5, WindowDout_4__0__4, 
               WindowDout_4__0__3, WindowDout_4__0__2, WindowDout_4__0__1, 
               WindowDout_4__0__0, WindowDout_4__1__7, WindowDout_4__1__6, 
               WindowDout_4__1__5, WindowDout_4__1__4, WindowDout_4__1__3, 
               WindowDout_4__1__2, WindowDout_4__1__1, WindowDout_4__1__0, 
               WindowDout_4__2__7, WindowDout_4__2__6, WindowDout_4__2__5, 
               WindowDout_4__2__4, WindowDout_4__2__3, WindowDout_4__2__2, 
               WindowDout_4__2__1, WindowDout_4__2__0, WindowDout_4__3__7, 
               WindowDout_4__3__6, WindowDout_4__3__5, WindowDout_4__3__4, 
               WindowDout_4__3__3, WindowDout_4__3__2, WindowDout_4__3__1, 
               WindowDout_4__3__0, WindowDout_4__4__7, WindowDout_4__4__6, 
               WindowDout_4__4__5, WindowDout_4__4__4, WindowDout_4__4__3, 
               WindowDout_4__4__2, WindowDout_4__4__1, WindowDout_4__4__0, 
               ResultWR, ResultDin, ResultDout ) ;

    input CLK ;
    input RST ;
    input FilterSize ;
    input FilterWR ;
    input WindowWR ;
    input [39:0]Din ;
    output FilterDout_0__0__7 ;
    output FilterDout_0__0__6 ;
    output FilterDout_0__0__5 ;
    output FilterDout_0__0__4 ;
    output FilterDout_0__0__3 ;
    output FilterDout_0__0__2 ;
    output FilterDout_0__0__1 ;
    output FilterDout_0__0__0 ;
    output FilterDout_0__1__7 ;
    output FilterDout_0__1__6 ;
    output FilterDout_0__1__5 ;
    output FilterDout_0__1__4 ;
    output FilterDout_0__1__3 ;
    output FilterDout_0__1__2 ;
    output FilterDout_0__1__1 ;
    output FilterDout_0__1__0 ;
    output FilterDout_0__2__7 ;
    output FilterDout_0__2__6 ;
    output FilterDout_0__2__5 ;
    output FilterDout_0__2__4 ;
    output FilterDout_0__2__3 ;
    output FilterDout_0__2__2 ;
    output FilterDout_0__2__1 ;
    output FilterDout_0__2__0 ;
    output FilterDout_0__3__7 ;
    output FilterDout_0__3__6 ;
    output FilterDout_0__3__5 ;
    output FilterDout_0__3__4 ;
    output FilterDout_0__3__3 ;
    output FilterDout_0__3__2 ;
    output FilterDout_0__3__1 ;
    output FilterDout_0__3__0 ;
    output FilterDout_0__4__7 ;
    output FilterDout_0__4__6 ;
    output FilterDout_0__4__5 ;
    output FilterDout_0__4__4 ;
    output FilterDout_0__4__3 ;
    output FilterDout_0__4__2 ;
    output FilterDout_0__4__1 ;
    output FilterDout_0__4__0 ;
    output FilterDout_1__0__7 ;
    output FilterDout_1__0__6 ;
    output FilterDout_1__0__5 ;
    output FilterDout_1__0__4 ;
    output FilterDout_1__0__3 ;
    output FilterDout_1__0__2 ;
    output FilterDout_1__0__1 ;
    output FilterDout_1__0__0 ;
    output FilterDout_1__1__7 ;
    output FilterDout_1__1__6 ;
    output FilterDout_1__1__5 ;
    output FilterDout_1__1__4 ;
    output FilterDout_1__1__3 ;
    output FilterDout_1__1__2 ;
    output FilterDout_1__1__1 ;
    output FilterDout_1__1__0 ;
    output FilterDout_1__2__7 ;
    output FilterDout_1__2__6 ;
    output FilterDout_1__2__5 ;
    output FilterDout_1__2__4 ;
    output FilterDout_1__2__3 ;
    output FilterDout_1__2__2 ;
    output FilterDout_1__2__1 ;
    output FilterDout_1__2__0 ;
    output FilterDout_1__3__7 ;
    output FilterDout_1__3__6 ;
    output FilterDout_1__3__5 ;
    output FilterDout_1__3__4 ;
    output FilterDout_1__3__3 ;
    output FilterDout_1__3__2 ;
    output FilterDout_1__3__1 ;
    output FilterDout_1__3__0 ;
    output FilterDout_1__4__7 ;
    output FilterDout_1__4__6 ;
    output FilterDout_1__4__5 ;
    output FilterDout_1__4__4 ;
    output FilterDout_1__4__3 ;
    output FilterDout_1__4__2 ;
    output FilterDout_1__4__1 ;
    output FilterDout_1__4__0 ;
    output FilterDout_2__0__7 ;
    output FilterDout_2__0__6 ;
    output FilterDout_2__0__5 ;
    output FilterDout_2__0__4 ;
    output FilterDout_2__0__3 ;
    output FilterDout_2__0__2 ;
    output FilterDout_2__0__1 ;
    output FilterDout_2__0__0 ;
    output FilterDout_2__1__7 ;
    output FilterDout_2__1__6 ;
    output FilterDout_2__1__5 ;
    output FilterDout_2__1__4 ;
    output FilterDout_2__1__3 ;
    output FilterDout_2__1__2 ;
    output FilterDout_2__1__1 ;
    output FilterDout_2__1__0 ;
    output FilterDout_2__2__7 ;
    output FilterDout_2__2__6 ;
    output FilterDout_2__2__5 ;
    output FilterDout_2__2__4 ;
    output FilterDout_2__2__3 ;
    output FilterDout_2__2__2 ;
    output FilterDout_2__2__1 ;
    output FilterDout_2__2__0 ;
    output FilterDout_2__3__7 ;
    output FilterDout_2__3__6 ;
    output FilterDout_2__3__5 ;
    output FilterDout_2__3__4 ;
    output FilterDout_2__3__3 ;
    output FilterDout_2__3__2 ;
    output FilterDout_2__3__1 ;
    output FilterDout_2__3__0 ;
    output FilterDout_2__4__7 ;
    output FilterDout_2__4__6 ;
    output FilterDout_2__4__5 ;
    output FilterDout_2__4__4 ;
    output FilterDout_2__4__3 ;
    output FilterDout_2__4__2 ;
    output FilterDout_2__4__1 ;
    output FilterDout_2__4__0 ;
    output FilterDout_3__0__7 ;
    output FilterDout_3__0__6 ;
    output FilterDout_3__0__5 ;
    output FilterDout_3__0__4 ;
    output FilterDout_3__0__3 ;
    output FilterDout_3__0__2 ;
    output FilterDout_3__0__1 ;
    output FilterDout_3__0__0 ;
    output FilterDout_3__1__7 ;
    output FilterDout_3__1__6 ;
    output FilterDout_3__1__5 ;
    output FilterDout_3__1__4 ;
    output FilterDout_3__1__3 ;
    output FilterDout_3__1__2 ;
    output FilterDout_3__1__1 ;
    output FilterDout_3__1__0 ;
    output FilterDout_3__2__7 ;
    output FilterDout_3__2__6 ;
    output FilterDout_3__2__5 ;
    output FilterDout_3__2__4 ;
    output FilterDout_3__2__3 ;
    output FilterDout_3__2__2 ;
    output FilterDout_3__2__1 ;
    output FilterDout_3__2__0 ;
    output FilterDout_3__3__7 ;
    output FilterDout_3__3__6 ;
    output FilterDout_3__3__5 ;
    output FilterDout_3__3__4 ;
    output FilterDout_3__3__3 ;
    output FilterDout_3__3__2 ;
    output FilterDout_3__3__1 ;
    output FilterDout_3__3__0 ;
    output FilterDout_3__4__7 ;
    output FilterDout_3__4__6 ;
    output FilterDout_3__4__5 ;
    output FilterDout_3__4__4 ;
    output FilterDout_3__4__3 ;
    output FilterDout_3__4__2 ;
    output FilterDout_3__4__1 ;
    output FilterDout_3__4__0 ;
    output FilterDout_4__0__7 ;
    output FilterDout_4__0__6 ;
    output FilterDout_4__0__5 ;
    output FilterDout_4__0__4 ;
    output FilterDout_4__0__3 ;
    output FilterDout_4__0__2 ;
    output FilterDout_4__0__1 ;
    output FilterDout_4__0__0 ;
    output FilterDout_4__1__7 ;
    output FilterDout_4__1__6 ;
    output FilterDout_4__1__5 ;
    output FilterDout_4__1__4 ;
    output FilterDout_4__1__3 ;
    output FilterDout_4__1__2 ;
    output FilterDout_4__1__1 ;
    output FilterDout_4__1__0 ;
    output FilterDout_4__2__7 ;
    output FilterDout_4__2__6 ;
    output FilterDout_4__2__5 ;
    output FilterDout_4__2__4 ;
    output FilterDout_4__2__3 ;
    output FilterDout_4__2__2 ;
    output FilterDout_4__2__1 ;
    output FilterDout_4__2__0 ;
    output FilterDout_4__3__7 ;
    output FilterDout_4__3__6 ;
    output FilterDout_4__3__5 ;
    output FilterDout_4__3__4 ;
    output FilterDout_4__3__3 ;
    output FilterDout_4__3__2 ;
    output FilterDout_4__3__1 ;
    output FilterDout_4__3__0 ;
    output FilterDout_4__4__7 ;
    output FilterDout_4__4__6 ;
    output FilterDout_4__4__5 ;
    output FilterDout_4__4__4 ;
    output FilterDout_4__4__3 ;
    output FilterDout_4__4__2 ;
    output FilterDout_4__4__1 ;
    output FilterDout_4__4__0 ;
    output WindowDout_0__0__7 ;
    output WindowDout_0__0__6 ;
    output WindowDout_0__0__5 ;
    output WindowDout_0__0__4 ;
    output WindowDout_0__0__3 ;
    output WindowDout_0__0__2 ;
    output WindowDout_0__0__1 ;
    output WindowDout_0__0__0 ;
    output WindowDout_0__1__7 ;
    output WindowDout_0__1__6 ;
    output WindowDout_0__1__5 ;
    output WindowDout_0__1__4 ;
    output WindowDout_0__1__3 ;
    output WindowDout_0__1__2 ;
    output WindowDout_0__1__1 ;
    output WindowDout_0__1__0 ;
    output WindowDout_0__2__7 ;
    output WindowDout_0__2__6 ;
    output WindowDout_0__2__5 ;
    output WindowDout_0__2__4 ;
    output WindowDout_0__2__3 ;
    output WindowDout_0__2__2 ;
    output WindowDout_0__2__1 ;
    output WindowDout_0__2__0 ;
    output WindowDout_0__3__7 ;
    output WindowDout_0__3__6 ;
    output WindowDout_0__3__5 ;
    output WindowDout_0__3__4 ;
    output WindowDout_0__3__3 ;
    output WindowDout_0__3__2 ;
    output WindowDout_0__3__1 ;
    output WindowDout_0__3__0 ;
    output WindowDout_0__4__7 ;
    output WindowDout_0__4__6 ;
    output WindowDout_0__4__5 ;
    output WindowDout_0__4__4 ;
    output WindowDout_0__4__3 ;
    output WindowDout_0__4__2 ;
    output WindowDout_0__4__1 ;
    output WindowDout_0__4__0 ;
    output WindowDout_1__0__7 ;
    output WindowDout_1__0__6 ;
    output WindowDout_1__0__5 ;
    output WindowDout_1__0__4 ;
    output WindowDout_1__0__3 ;
    output WindowDout_1__0__2 ;
    output WindowDout_1__0__1 ;
    output WindowDout_1__0__0 ;
    output WindowDout_1__1__7 ;
    output WindowDout_1__1__6 ;
    output WindowDout_1__1__5 ;
    output WindowDout_1__1__4 ;
    output WindowDout_1__1__3 ;
    output WindowDout_1__1__2 ;
    output WindowDout_1__1__1 ;
    output WindowDout_1__1__0 ;
    output WindowDout_1__2__7 ;
    output WindowDout_1__2__6 ;
    output WindowDout_1__2__5 ;
    output WindowDout_1__2__4 ;
    output WindowDout_1__2__3 ;
    output WindowDout_1__2__2 ;
    output WindowDout_1__2__1 ;
    output WindowDout_1__2__0 ;
    output WindowDout_1__3__7 ;
    output WindowDout_1__3__6 ;
    output WindowDout_1__3__5 ;
    output WindowDout_1__3__4 ;
    output WindowDout_1__3__3 ;
    output WindowDout_1__3__2 ;
    output WindowDout_1__3__1 ;
    output WindowDout_1__3__0 ;
    output WindowDout_1__4__7 ;
    output WindowDout_1__4__6 ;
    output WindowDout_1__4__5 ;
    output WindowDout_1__4__4 ;
    output WindowDout_1__4__3 ;
    output WindowDout_1__4__2 ;
    output WindowDout_1__4__1 ;
    output WindowDout_1__4__0 ;
    output WindowDout_2__0__7 ;
    output WindowDout_2__0__6 ;
    output WindowDout_2__0__5 ;
    output WindowDout_2__0__4 ;
    output WindowDout_2__0__3 ;
    output WindowDout_2__0__2 ;
    output WindowDout_2__0__1 ;
    output WindowDout_2__0__0 ;
    output WindowDout_2__1__7 ;
    output WindowDout_2__1__6 ;
    output WindowDout_2__1__5 ;
    output WindowDout_2__1__4 ;
    output WindowDout_2__1__3 ;
    output WindowDout_2__1__2 ;
    output WindowDout_2__1__1 ;
    output WindowDout_2__1__0 ;
    output WindowDout_2__2__7 ;
    output WindowDout_2__2__6 ;
    output WindowDout_2__2__5 ;
    output WindowDout_2__2__4 ;
    output WindowDout_2__2__3 ;
    output WindowDout_2__2__2 ;
    output WindowDout_2__2__1 ;
    output WindowDout_2__2__0 ;
    output WindowDout_2__3__7 ;
    output WindowDout_2__3__6 ;
    output WindowDout_2__3__5 ;
    output WindowDout_2__3__4 ;
    output WindowDout_2__3__3 ;
    output WindowDout_2__3__2 ;
    output WindowDout_2__3__1 ;
    output WindowDout_2__3__0 ;
    output WindowDout_2__4__7 ;
    output WindowDout_2__4__6 ;
    output WindowDout_2__4__5 ;
    output WindowDout_2__4__4 ;
    output WindowDout_2__4__3 ;
    output WindowDout_2__4__2 ;
    output WindowDout_2__4__1 ;
    output WindowDout_2__4__0 ;
    output WindowDout_3__0__7 ;
    output WindowDout_3__0__6 ;
    output WindowDout_3__0__5 ;
    output WindowDout_3__0__4 ;
    output WindowDout_3__0__3 ;
    output WindowDout_3__0__2 ;
    output WindowDout_3__0__1 ;
    output WindowDout_3__0__0 ;
    output WindowDout_3__1__7 ;
    output WindowDout_3__1__6 ;
    output WindowDout_3__1__5 ;
    output WindowDout_3__1__4 ;
    output WindowDout_3__1__3 ;
    output WindowDout_3__1__2 ;
    output WindowDout_3__1__1 ;
    output WindowDout_3__1__0 ;
    output WindowDout_3__2__7 ;
    output WindowDout_3__2__6 ;
    output WindowDout_3__2__5 ;
    output WindowDout_3__2__4 ;
    output WindowDout_3__2__3 ;
    output WindowDout_3__2__2 ;
    output WindowDout_3__2__1 ;
    output WindowDout_3__2__0 ;
    output WindowDout_3__3__7 ;
    output WindowDout_3__3__6 ;
    output WindowDout_3__3__5 ;
    output WindowDout_3__3__4 ;
    output WindowDout_3__3__3 ;
    output WindowDout_3__3__2 ;
    output WindowDout_3__3__1 ;
    output WindowDout_3__3__0 ;
    output WindowDout_3__4__7 ;
    output WindowDout_3__4__6 ;
    output WindowDout_3__4__5 ;
    output WindowDout_3__4__4 ;
    output WindowDout_3__4__3 ;
    output WindowDout_3__4__2 ;
    output WindowDout_3__4__1 ;
    output WindowDout_3__4__0 ;
    output WindowDout_4__0__7 ;
    output WindowDout_4__0__6 ;
    output WindowDout_4__0__5 ;
    output WindowDout_4__0__4 ;
    output WindowDout_4__0__3 ;
    output WindowDout_4__0__2 ;
    output WindowDout_4__0__1 ;
    output WindowDout_4__0__0 ;
    output WindowDout_4__1__7 ;
    output WindowDout_4__1__6 ;
    output WindowDout_4__1__5 ;
    output WindowDout_4__1__4 ;
    output WindowDout_4__1__3 ;
    output WindowDout_4__1__2 ;
    output WindowDout_4__1__1 ;
    output WindowDout_4__1__0 ;
    output WindowDout_4__2__7 ;
    output WindowDout_4__2__6 ;
    output WindowDout_4__2__5 ;
    output WindowDout_4__2__4 ;
    output WindowDout_4__2__3 ;
    output WindowDout_4__2__2 ;
    output WindowDout_4__2__1 ;
    output WindowDout_4__2__0 ;
    output WindowDout_4__3__7 ;
    output WindowDout_4__3__6 ;
    output WindowDout_4__3__5 ;
    output WindowDout_4__3__4 ;
    output WindowDout_4__3__3 ;
    output WindowDout_4__3__2 ;
    output WindowDout_4__3__1 ;
    output WindowDout_4__3__0 ;
    output WindowDout_4__4__7 ;
    output WindowDout_4__4__6 ;
    output WindowDout_4__4__5 ;
    output WindowDout_4__4__4 ;
    output WindowDout_4__4__3 ;
    output WindowDout_4__4__2 ;
    output WindowDout_4__4__1 ;
    output WindowDout_4__4__0 ;
    input ResultWR ;
    input [7:0]ResultDin ;
    output [7:0]ResultDout ;

    wire nx84, nx88, nx98, nx108, nx118, nx128, nx138, nx148, nx158, nx168, 
         nx220, nx230, nx240, nx250, nx260, nx270, nx280, nx290, nx1931, nx1941, 
         nx1951, nx1961, nx1971, nx1981, nx1991, nx2001, nx2011, nx2021, nx2031, 
         nx2041, nx2051, nx2061, nx2071, nx2081, nx2091, nx2101, nx2111, nx2121, 
         nx2131, nx2141, nx2151, nx2161, nx2171, nx2181, nx2191, nx2201, nx2211, 
         nx2221, nx2231, nx2241, nx2251, nx2261, nx2271, nx2281, nx2291, nx2301, 
         nx2311, nx2321, nx2331, nx2341, nx2351, nx2361, nx2371, nx2381, nx2391, 
         nx2401, nx2411, nx2421, nx2431, nx2441, nx2451, nx2461, nx2471, nx2481, 
         nx2491, nx2501, nx2511, nx2521, nx2531, nx2541, nx2551, nx2561, nx2571, 
         nx2581, nx2591, nx2601, nx2611, nx2621, nx2631, nx2641, nx2651, nx2661, 
         nx2671, nx2681, nx2691, nx2701, nx2711, nx2721, nx2731, nx2741, nx2751, 
         nx2761, nx2771, nx2781, nx2791, nx2801, nx2811, nx2821, nx2831, nx2841, 
         nx2851, nx2861, nx2871, nx2881, nx2891, nx2901, nx2911, nx2921, nx2931, 
         nx2941, nx2951, nx2961, nx2971, nx2981, nx2991, nx3001, nx3011, nx3021, 
         nx3031, nx3041, nx3051, nx3061, nx3071, nx3081, nx3091, nx3101, nx3111, 
         nx3121, nx3131, nx3141, nx3151, nx3161, nx3171, nx3181, nx3191, nx3201, 
         nx3211, nx3221, nx3231, nx3241, nx3251, nx3261, nx3271, nx3281, nx3291, 
         nx3301, nx3311, nx3321, nx3331, nx3341, nx3351, nx3361, nx3371, nx3381, 
         nx3391, nx3401, nx3411, nx3421, nx3431, nx3441, nx3451, nx3461, nx3471, 
         nx3481, nx3491, nx3501, nx3511, nx3521, nx3531, nx3541, nx3551, nx3561, 
         nx3571, nx3581, nx3591, nx3601, nx3611, nx3621, nx3631, nx3641, nx3651, 
         nx3661, nx3671, nx3681, nx3691, nx3701, nx3711, nx3721, nx3731, nx3741, 
         nx3751, nx3761, nx3771, nx3781, nx3791, nx3801, nx3811, nx3821, nx3831, 
         nx3841, nx3851, nx3861, nx3871, nx3881, nx3891, nx3901, nx3911, nx3921, 
         nx3931, nx3941, nx3951, nx3961, nx3971, nx3981, nx3991, nx4001, nx4011, 
         nx4021, nx4031, nx4041, nx4051, nx4061, nx4071, nx4081, nx4091, nx4101, 
         nx4111, nx4121, nx4131, nx4141, nx4151, nx4161, nx4171, nx4181, nx4191, 
         nx4201, nx4211, nx4221, nx4231, nx4241, nx4251, nx4261, nx4271, nx4281, 
         nx4291, nx4301, nx4311, nx4321, nx4331, nx4341, nx4351, nx4361, nx4371, 
         nx4381, nx4391, nx4401, nx4411, nx4421, nx4431, nx4441, nx4451, nx4461, 
         nx4471, nx4481, nx4491, nx4501, nx4511, nx4521, nx4531, nx4541, nx4551, 
         nx4561, nx4571, nx4581, nx4591, nx4601, nx4611, nx4621, nx4631, nx4641, 
         nx4651, nx4661, nx4671, nx4681, nx4691, nx4701, nx4711, nx4721, nx4731, 
         nx4741, nx4751, nx4761, nx4771, nx4781, nx4791, nx4801, nx4811, nx4821, 
         nx4831, nx4841, nx4851, nx4861, nx4871, nx4881, nx4891, nx4901, nx4911, 
         nx4921, nx4931, nx4941, nx4951, nx4961, nx4971, nx4981, nx4991, nx5001, 
         nx5011, nx5021, nx5031, nx5041, nx5051, nx5061, nx5071, nx5081, nx5091, 
         nx5101, nx5111, nx5121, nx5131, nx5141, nx5151, nx5161, nx5171, nx5181, 
         nx5191, nx5201, nx5211, nx5221, nx5231, nx5241, nx5251, nx5261, nx5271, 
         nx5281, nx5291, nx5301, nx5311, nx5321, nx5331, nx5341, nx5351, nx5361, 
         nx5371, nx5381, nx5391, nx5401, nx5411, nx5421, nx5431, nx5441, nx5451, 
         nx5461, nx5471, nx5481, nx5491, nx5501, nx5511, nx5521, nx5531, nx5541, 
         nx5551, nx5561, nx5571, nx5581, nx5591, nx5601, nx5611, nx5621, nx5631, 
         nx5641, nx5651, nx5661, nx5671, nx5681, nx5691, nx5701, nx5711, nx5721, 
         nx5731, nx5741, nx5751, nx5761, nx5771, nx5781, nx5791, nx5801, nx5811, 
         nx5821, nx5831, nx5841, nx5851, nx5861, nx5871, nx5881, nx5891, nx5901, 
         nx5911, nx5921, nx5931, nx5941, nx5951, nx5961, nx5971, nx5981, nx5991, 
         nx6001, nx6015, nx6042, nx6107, nx6181, nx6184, nx6188, nx6190, nx6194, 
         nx6196, nx6200, nx6202, nx6206, nx6208, nx6212, nx6214, nx6218, nx6220, 
         nx6224, nx6226, nx6230, nx6232, nx6236, nx6238, nx6242, nx6244, nx6248, 
         nx6250, nx6254, nx6256, nx6260, nx6262, nx6266, nx6268, nx6272, nx6274, 
         nx6350, nx6352, nx6356, nx6358, nx6362, nx6364, nx6368, nx6370, nx6374, 
         nx6376, nx6380, nx6382, nx6386, nx6388, nx6392, nx6394, nx6398, nx6400, 
         nx6404, nx6406, nx6410, nx6412, nx6416, nx6418, nx6422, nx6424, nx6428, 
         nx6430, nx6434, nx6436, nx6440, nx6442, nx6518, nx6520, nx6524, nx6526, 
         nx6530, nx6532, nx6536, nx6538, nx6542, nx6544, nx6548, nx6550, nx6554, 
         nx6556, nx6560, nx6562, nx6566, nx6568, nx6572, nx6574, nx6578, nx6580, 
         nx6584, nx6586, nx6590, nx6592, nx6596, nx6598, nx6602, nx6604, nx6608, 
         nx6610, nx6614, nx6616, nx6620, nx6622, nx6626, nx6628, nx6632, nx6634, 
         nx6638, nx6640, nx6644, nx6646, nx6650, nx6652, nx6656, nx6658, nx6662, 
         nx6664, nx6668, nx6670, nx6674, nx6676, nx6680, nx6682, nx6686, nx6688, 
         nx6692, nx6694, nx6698, nx6700, nx6704, nx6706, nx6710, nx6712, nx6716, 
         nx6718, nx6722, nx6724, nx6728, nx6730, nx6734, nx6736, nx6740, nx6742, 
         nx6746, nx6748, nx6752, nx6754, nx6758, nx6760, nx6764, nx6766, nx6770, 
         nx6772, nx6776, nx6778, nx6782, nx6784, nx6788, nx6790, nx6794, nx6796, 
         nx6800, nx6802, nx6806, nx6808, nx6812, nx6814, nx6818, nx6820, nx6824, 
         nx6826, nx6830, nx6832, nx6836, nx6838, nx6842, nx6844, nx6848, nx6850, 
         nx6854, nx6856, nx6860, nx6862, nx6866, nx6868, nx6872, nx6874, nx6878, 
         nx6880, nx6884, nx6886, nx6890, nx6892, nx6896, nx6898, nx6902, nx6904, 
         nx6908, nx6910, nx6914, nx6916, nx6920, nx6922, nx6926, nx6928, nx6932, 
         nx6934, nx6938, nx6940, nx6944, nx6946, nx6950, nx6952, nx6956, nx6958, 
         nx6962, nx6964, nx6968, nx6970, nx6974, nx6976, nx6980, nx6982, nx6986, 
         nx6988, nx6992, nx6994, nx6998, nx7048, nx7122, nx7125, nx7129, nx7131, 
         nx7135, nx7137, nx7141, nx7143, nx7147, nx7149, nx7153, nx7155, nx7159, 
         nx7161, nx7165, nx7167, nx7171, nx7173, nx7177, nx7179, nx7183, nx7185, 
         nx7189, nx7191, nx7195, nx7197, nx7201, nx7203, nx7207, nx7209, nx7213, 
         nx7215, nx7291, nx7293, nx7297, nx7299, nx7303, nx7305, nx7309, nx7311, 
         nx7315, nx7317, nx7321, nx7323, nx7327, nx7329, nx7333, nx7335, nx7339, 
         nx7341, nx7345, nx7347, nx7351, nx7353, nx7357, nx7359, nx7363, nx7365, 
         nx7369, nx7371, nx7375, nx7377, nx7381, nx7383, nx7459, nx7461, nx7465, 
         nx7467, nx7471, nx7473, nx7477, nx7479, nx7483, nx7485, nx7489, nx7491, 
         nx7495, nx7497, nx7501, nx7503, nx7507, nx7509, nx7513, nx7515, nx7519, 
         nx7521, nx7525, nx7527, nx7531, nx7533, nx7537, nx7539, nx7543, nx7545, 
         nx7549, nx7551, nx7555, nx7557, nx7561, nx7563, nx7567, nx7569, nx7573, 
         nx7575, nx7579, nx7581, nx7585, nx7587, nx7591, nx7593, nx7597, nx7599, 
         nx7603, nx7605, nx7609, nx7611, nx7615, nx7617, nx7621, nx7623, nx7627, 
         nx7629, nx7633, nx7635, nx7639, nx7641, nx7645, nx7647, nx7651, nx7653, 
         nx7657, nx7659, nx7663, nx7665, nx7669, nx7671, nx7675, nx7677, nx7681, 
         nx7683, nx7687, nx7689, nx7693, nx7695, nx7699, nx7701, nx7705, nx7707, 
         nx7711, nx7713, nx7717, nx7719, nx7723, nx7725, nx7729, nx7731, nx7735, 
         nx7737, nx7741, nx7743, nx7747, nx7749, nx7753, nx7755, nx7759, nx7761, 
         nx7765, nx7767, nx7771, nx7773, nx7777, nx7779, nx7783, nx7785, nx7789, 
         nx7791, nx7795, nx7797, nx7801, nx7803, nx7807, nx7809, nx7813, nx7815, 
         nx7819, nx7821, nx7825, nx7827, nx7831, nx7833, nx7837, nx7839, nx7843, 
         nx7845, nx7849, nx7851, nx7855, nx7857, nx7861, nx7863, nx7867, nx7869, 
         nx7873, nx7875, nx7879, nx7881, nx7885, nx7887, nx7891, nx7893, nx7897, 
         nx7899, nx7903, nx7905, nx7909, nx7911, nx7915, nx7917, nx7921, nx7923, 
         nx7927, nx7929, nx7933, nx7935, nx7942, nx7944, nx7946, nx7948, nx7950, 
         nx7952, nx7954, nx7956, nx7958, nx7960, nx7962, nx7964, nx7966, nx7968, 
         nx7970, nx7972, nx7974, nx7976, nx7978, nx7980, nx7982, nx7984, nx7986, 
         nx7988, nx7990, nx7992, nx7994, nx7996, nx7998, nx8000, nx8002, nx8004, 
         nx8006, nx8008, nx8010, nx8012, nx8014, nx8016, nx8018, nx8020, nx8022, 
         nx8024, nx8026, nx8028, nx8030, nx8032, nx8034, nx8036, nx8038, nx8040, 
         nx8042, nx8044, nx8046, nx8048, nx8050, nx8052, nx8054, nx8056, nx8058, 
         nx8060, nx8062, nx8064, nx8066, nx8068, nx8070, nx8072, nx8074, nx8076, 
         nx8078, nx8080, nx8082, nx8084, nx8086, nx8088, nx8090, nx8094, nx8096, 
         nx8098, nx8100, nx8106, nx8108, nx8110, nx8112, nx8124, nx8126, nx8128, 
         nx8130, nx8132, nx8134, nx8136, nx8138, nx8140, nx8142, nx8146, nx8148, 
         nx8150, nx8152, nx8154, nx8158, nx8160, nx8162, nx8164, nx8182, nx8184, 
         nx8186, nx8188, nx8190, nx8194, nx8196, nx8198, nx8200, nx8202, nx8204, 
         nx8206, nx8208, nx8210, nx8212, nx8214, nx8220, nx8222, nx8224, nx8226, 
         nx8228, nx8232, nx8234, nx8236, nx8238, nx8240, nx8242, nx8244, nx8246, 
         nx8248, nx8250, nx8252, nx8254, nx8256, nx8258, nx8260, nx8270, nx8272, 
         nx8274, nx8276, nx8278, nx8280, nx8282, nx8284, nx8286, nx8288, nx8290, 
         nx8292, nx8294, nx8296, nx8298, nx8300, nx8302, nx8304, nx8306, nx8308, 
         nx8310, nx8312, nx8314, nx8316, nx8318, nx8320, nx8322, nx8324, nx8326, 
         nx8328, nx8334, nx8336;
    wire [183:0] \$dummy ;




    dff RESULT_REG_reg_Dout_0 (.Q (ResultDout[0]), .QB (\$dummy [0]), .D (nx1931
        ), .CLK (CLK)) ;
    ao32 ix1932 (.Y (nx1931), .A0 (ResultDin[0]), .A1 (nx8070), .A2 (ResultWR), 
         .B0 (ResultDout[0]), .B1 (nx6015)) ;
    nor02_2x ix6016 (.Y (nx6015), .A0 (RST), .A1 (ResultWR)) ;
    dff RESULT_REG_reg_Dout_1 (.Q (ResultDout[1]), .QB (\$dummy [1]), .D (nx1941
        ), .CLK (CLK)) ;
    ao32 ix1942 (.Y (nx1941), .A0 (ResultDin[1]), .A1 (nx8070), .A2 (ResultWR), 
         .B0 (ResultDout[1]), .B1 (nx6015)) ;
    dff RESULT_REG_reg_Dout_2 (.Q (ResultDout[2]), .QB (\$dummy [2]), .D (nx1951
        ), .CLK (CLK)) ;
    ao32 ix1952 (.Y (nx1951), .A0 (ResultDin[2]), .A1 (nx8070), .A2 (ResultWR), 
         .B0 (ResultDout[2]), .B1 (nx6015)) ;
    dff RESULT_REG_reg_Dout_3 (.Q (ResultDout[3]), .QB (\$dummy [3]), .D (nx1961
        ), .CLK (CLK)) ;
    ao32 ix1962 (.Y (nx1961), .A0 (ResultDin[3]), .A1 (nx8070), .A2 (ResultWR), 
         .B0 (ResultDout[3]), .B1 (nx6015)) ;
    dff RESULT_REG_reg_Dout_4 (.Q (ResultDout[4]), .QB (\$dummy [4]), .D (nx1971
        ), .CLK (CLK)) ;
    ao32 ix1972 (.Y (nx1971), .A0 (ResultDin[4]), .A1 (nx8070), .A2 (ResultWR), 
         .B0 (ResultDout[4]), .B1 (nx6015)) ;
    dff RESULT_REG_reg_Dout_5 (.Q (ResultDout[5]), .QB (\$dummy [5]), .D (nx1981
        ), .CLK (CLK)) ;
    ao32 ix1982 (.Y (nx1981), .A0 (ResultDin[5]), .A1 (nx8070), .A2 (ResultWR), 
         .B0 (ResultDout[5]), .B1 (nx6015)) ;
    dff RESULT_REG_reg_Dout_6 (.Q (ResultDout[6]), .QB (\$dummy [6]), .D (nx1991
        ), .CLK (CLK)) ;
    ao32 ix1992 (.Y (nx1991), .A0 (ResultDin[6]), .A1 (nx8070), .A2 (ResultWR), 
         .B0 (ResultDout[6]), .B1 (nx6015)) ;
    dff RESULT_REG_reg_Dout_7 (.Q (ResultDout[7]), .QB (\$dummy [7]), .D (nx2001
        ), .CLK (CLK)) ;
    ao32 ix2002 (.Y (nx2001), .A0 (ResultDin[7]), .A1 (nx8072), .A2 (ResultWR), 
         .B0 (ResultDout[7]), .B1 (nx6015)) ;
    dff L0_4_L1_4_Wij_reg_Dout_0 (.Q (WindowDout_4__4__0), .QB (\$dummy [8]), .D (
        nx2011), .CLK (CLK)) ;
    nor02ii ix89 (.Y (nx88), .A0 (RST), .A1 (Din[32])) ;
    aoi21 ix6043 (.Y (nx6042), .A0 (WindowWR), .A1 (FilterSize), .B0 (RST)) ;
    dff L0_4_L1_4_Wij_reg_Dout_1 (.Q (WindowDout_4__4__1), .QB (\$dummy [9]), .D (
        nx2021), .CLK (CLK)) ;
    nor02ii ix99 (.Y (nx98), .A0 (RST), .A1 (Din[33])) ;
    dff L0_4_L1_4_Wij_reg_Dout_2 (.Q (WindowDout_4__4__2), .QB (\$dummy [10]), .D (
        nx2031), .CLK (CLK)) ;
    nor02ii ix109 (.Y (nx108), .A0 (RST), .A1 (Din[34])) ;
    dff L0_4_L1_4_Wij_reg_Dout_3 (.Q (WindowDout_4__4__3), .QB (\$dummy [11]), .D (
        nx2041), .CLK (CLK)) ;
    nor02ii ix119 (.Y (nx118), .A0 (RST), .A1 (Din[35])) ;
    dff L0_4_L1_4_Wij_reg_Dout_4 (.Q (WindowDout_4__4__4), .QB (\$dummy [12]), .D (
        nx2051), .CLK (CLK)) ;
    nor02ii ix129 (.Y (nx128), .A0 (RST), .A1 (Din[36])) ;
    dff L0_4_L1_4_Wij_reg_Dout_5 (.Q (WindowDout_4__4__5), .QB (\$dummy [13]), .D (
        nx2061), .CLK (CLK)) ;
    nor02ii ix139 (.Y (nx138), .A0 (RST), .A1 (Din[37])) ;
    dff L0_4_L1_4_Wij_reg_Dout_6 (.Q (WindowDout_4__4__6), .QB (\$dummy [14]), .D (
        nx2071), .CLK (CLK)) ;
    nor02ii ix149 (.Y (nx148), .A0 (RST), .A1 (Din[38])) ;
    dff L0_4_L1_4_Wij_reg_Dout_7 (.Q (WindowDout_4__4__7), .QB (\$dummy [15]), .D (
        nx2081), .CLK (CLK)) ;
    nor02ii ix159 (.Y (nx158), .A0 (RST), .A1 (Din[39])) ;
    dff L0_4_L1_3_Wij_reg_Dout_0 (.Q (WindowDout_4__3__0), .QB (\$dummy [16]), .D (
        nx2171), .CLK (CLK)) ;
    nor02ii ix221 (.Y (nx220), .A0 (RST), .A1 (Din[24])) ;
    dff L0_4_L1_3_Wij_reg_Dout_1 (.Q (WindowDout_4__3__1), .QB (\$dummy [17]), .D (
        nx2181), .CLK (CLK)) ;
    nor02ii ix231 (.Y (nx230), .A0 (RST), .A1 (Din[25])) ;
    dff L0_4_L1_3_Wij_reg_Dout_2 (.Q (WindowDout_4__3__2), .QB (\$dummy [18]), .D (
        nx2191), .CLK (CLK)) ;
    nor02ii ix241 (.Y (nx240), .A0 (RST), .A1 (Din[26])) ;
    dff L0_4_L1_3_Wij_reg_Dout_3 (.Q (WindowDout_4__3__3), .QB (\$dummy [19]), .D (
        nx2201), .CLK (CLK)) ;
    nor02ii ix251 (.Y (nx250), .A0 (RST), .A1 (Din[27])) ;
    dff L0_4_L1_3_Wij_reg_Dout_4 (.Q (WindowDout_4__3__4), .QB (\$dummy [20]), .D (
        nx2211), .CLK (CLK)) ;
    nor02ii ix261 (.Y (nx260), .A0 (RST), .A1 (Din[28])) ;
    dff L0_4_L1_3_Wij_reg_Dout_5 (.Q (WindowDout_4__3__5), .QB (\$dummy [21]), .D (
        nx2221), .CLK (CLK)) ;
    nor02ii ix271 (.Y (nx270), .A0 (RST), .A1 (Din[29])) ;
    dff L0_4_L1_3_Wij_reg_Dout_6 (.Q (WindowDout_4__3__6), .QB (\$dummy [22]), .D (
        nx2231), .CLK (CLK)) ;
    nor02ii ix281 (.Y (nx280), .A0 (RST), .A1 (Din[30])) ;
    dff L0_4_L1_3_Wij_reg_Dout_7 (.Q (WindowDout_4__3__7), .QB (\$dummy [23]), .D (
        nx2241), .CLK (CLK)) ;
    nor02ii ix291 (.Y (nx290), .A0 (RST), .A1 (Din[31])) ;
    dff L0_4_L1_2_Wij_reg_Dout_0 (.Q (WindowDout_4__2__0), .QB (\$dummy [24]), .D (
        nx2331), .CLK (CLK)) ;
    ao32 ix2332 (.Y (nx2331), .A0 (Din[16]), .A1 (nx8072), .A2 (WindowWR), .B0 (
         WindowDout_4__2__0), .B1 (nx8194)) ;
    nor02_2x ix6108 (.Y (nx6107), .A0 (WindowWR), .A1 (RST)) ;
    dff L0_4_L1_2_Wij_reg_Dout_1 (.Q (WindowDout_4__2__1), .QB (\$dummy [25]), .D (
        nx2341), .CLK (CLK)) ;
    ao32 ix2342 (.Y (nx2341), .A0 (Din[17]), .A1 (nx8072), .A2 (WindowWR), .B0 (
         WindowDout_4__2__1), .B1 (nx8194)) ;
    dff L0_4_L1_2_Wij_reg_Dout_2 (.Q (WindowDout_4__2__2), .QB (\$dummy [26]), .D (
        nx2351), .CLK (CLK)) ;
    ao32 ix2352 (.Y (nx2351), .A0 (Din[18]), .A1 (nx8072), .A2 (WindowWR), .B0 (
         WindowDout_4__2__2), .B1 (nx8194)) ;
    dff L0_4_L1_2_Wij_reg_Dout_3 (.Q (WindowDout_4__2__3), .QB (\$dummy [27]), .D (
        nx2361), .CLK (CLK)) ;
    ao32 ix2362 (.Y (nx2361), .A0 (Din[19]), .A1 (nx8072), .A2 (WindowWR), .B0 (
         WindowDout_4__2__3), .B1 (nx8194)) ;
    dff L0_4_L1_2_Wij_reg_Dout_4 (.Q (WindowDout_4__2__4), .QB (\$dummy [28]), .D (
        nx2371), .CLK (CLK)) ;
    ao32 ix2372 (.Y (nx2371), .A0 (Din[20]), .A1 (nx8072), .A2 (WindowWR), .B0 (
         WindowDout_4__2__4), .B1 (nx8194)) ;
    dff L0_4_L1_2_Wij_reg_Dout_5 (.Q (WindowDout_4__2__5), .QB (\$dummy [29]), .D (
        nx2381), .CLK (CLK)) ;
    ao32 ix2382 (.Y (nx2381), .A0 (Din[21]), .A1 (nx8072), .A2 (WindowWR), .B0 (
         WindowDout_4__2__5), .B1 (nx8194)) ;
    dff L0_4_L1_2_Wij_reg_Dout_6 (.Q (WindowDout_4__2__6), .QB (\$dummy [30]), .D (
        nx2391), .CLK (CLK)) ;
    ao32 ix2392 (.Y (nx2391), .A0 (Din[22]), .A1 (nx8074), .A2 (WindowWR), .B0 (
         WindowDout_4__2__6), .B1 (nx8194)) ;
    dff L0_4_L1_2_Wij_reg_Dout_7 (.Q (WindowDout_4__2__7), .QB (\$dummy [31]), .D (
        nx2401), .CLK (CLK)) ;
    ao32 ix2402 (.Y (nx2401), .A0 (Din[23]), .A1 (nx8074), .A2 (WindowWR), .B0 (
         WindowDout_4__2__7), .B1 (nx8196)) ;
    dff L0_4_L1_1_Wij_reg_Dout_0 (.Q (WindowDout_4__1__0), .QB (\$dummy [32]), .D (
        nx2491), .CLK (CLK)) ;
    ao32 ix2492 (.Y (nx2491), .A0 (Din[8]), .A1 (nx8074), .A2 (WindowWR), .B0 (
         WindowDout_4__1__0), .B1 (nx8196)) ;
    dff L0_4_L1_1_Wij_reg_Dout_1 (.Q (WindowDout_4__1__1), .QB (\$dummy [33]), .D (
        nx2501), .CLK (CLK)) ;
    ao32 ix2502 (.Y (nx2501), .A0 (Din[9]), .A1 (nx8074), .A2 (WindowWR), .B0 (
         WindowDout_4__1__1), .B1 (nx8196)) ;
    dff L0_4_L1_1_Wij_reg_Dout_2 (.Q (WindowDout_4__1__2), .QB (\$dummy [34]), .D (
        nx2511), .CLK (CLK)) ;
    ao32 ix2512 (.Y (nx2511), .A0 (Din[10]), .A1 (nx8074), .A2 (WindowWR), .B0 (
         WindowDout_4__1__2), .B1 (nx8196)) ;
    dff L0_4_L1_1_Wij_reg_Dout_3 (.Q (WindowDout_4__1__3), .QB (\$dummy [35]), .D (
        nx2521), .CLK (CLK)) ;
    ao32 ix2522 (.Y (nx2521), .A0 (Din[11]), .A1 (nx8074), .A2 (WindowWR), .B0 (
         WindowDout_4__1__3), .B1 (nx8196)) ;
    dff L0_4_L1_1_Wij_reg_Dout_4 (.Q (WindowDout_4__1__4), .QB (\$dummy [36]), .D (
        nx2531), .CLK (CLK)) ;
    ao32 ix2532 (.Y (nx2531), .A0 (Din[12]), .A1 (nx8074), .A2 (WindowWR), .B0 (
         WindowDout_4__1__4), .B1 (nx8196)) ;
    dff L0_4_L1_1_Wij_reg_Dout_5 (.Q (WindowDout_4__1__5), .QB (\$dummy [37]), .D (
        nx2541), .CLK (CLK)) ;
    ao32 ix2542 (.Y (nx2541), .A0 (Din[13]), .A1 (nx8076), .A2 (WindowWR), .B0 (
         WindowDout_4__1__5), .B1 (nx8196)) ;
    dff L0_4_L1_1_Wij_reg_Dout_6 (.Q (WindowDout_4__1__6), .QB (\$dummy [38]), .D (
        nx2551), .CLK (CLK)) ;
    ao32 ix2552 (.Y (nx2551), .A0 (Din[14]), .A1 (nx8076), .A2 (WindowWR), .B0 (
         WindowDout_4__1__6), .B1 (nx8198)) ;
    dff L0_4_L1_1_Wij_reg_Dout_7 (.Q (WindowDout_4__1__7), .QB (\$dummy [39]), .D (
        nx2561), .CLK (CLK)) ;
    ao32 ix2562 (.Y (nx2561), .A0 (Din[15]), .A1 (nx8076), .A2 (WindowWR), .B0 (
         WindowDout_4__1__7), .B1 (nx8198)) ;
    dff L0_4_L1_0_Wij_reg_Dout_0 (.Q (WindowDout_4__0__0), .QB (\$dummy [40]), .D (
        nx2651), .CLK (CLK)) ;
    ao32 ix2652 (.Y (nx2651), .A0 (Din[0]), .A1 (nx8076), .A2 (WindowWR), .B0 (
         WindowDout_4__0__0), .B1 (nx8198)) ;
    dff L0_4_L1_0_Wij_reg_Dout_1 (.Q (WindowDout_4__0__1), .QB (\$dummy [41]), .D (
        nx2661), .CLK (CLK)) ;
    ao32 ix2662 (.Y (nx2661), .A0 (Din[1]), .A1 (nx8076), .A2 (WindowWR), .B0 (
         WindowDout_4__0__1), .B1 (nx8198)) ;
    dff L0_4_L1_0_Wij_reg_Dout_2 (.Q (WindowDout_4__0__2), .QB (\$dummy [42]), .D (
        nx2671), .CLK (CLK)) ;
    ao32 ix2672 (.Y (nx2671), .A0 (Din[2]), .A1 (nx8076), .A2 (WindowWR), .B0 (
         WindowDout_4__0__2), .B1 (nx8198)) ;
    dff L0_4_L1_0_Wij_reg_Dout_3 (.Q (WindowDout_4__0__3), .QB (\$dummy [43]), .D (
        nx2681), .CLK (CLK)) ;
    ao32 ix2682 (.Y (nx2681), .A0 (Din[3]), .A1 (nx8076), .A2 (WindowWR), .B0 (
         WindowDout_4__0__3), .B1 (nx8198)) ;
    dff L0_4_L1_0_Wij_reg_Dout_4 (.Q (WindowDout_4__0__4), .QB (\$dummy [44]), .D (
        nx2691), .CLK (CLK)) ;
    ao32 ix2692 (.Y (nx2691), .A0 (Din[4]), .A1 (nx8078), .A2 (WindowWR), .B0 (
         WindowDout_4__0__4), .B1 (nx8198)) ;
    dff L0_4_L1_0_Wij_reg_Dout_5 (.Q (WindowDout_4__0__5), .QB (\$dummy [45]), .D (
        nx2701), .CLK (CLK)) ;
    ao32 ix2702 (.Y (nx2701), .A0 (Din[5]), .A1 (nx8078), .A2 (WindowWR), .B0 (
         WindowDout_4__0__5), .B1 (nx8200)) ;
    dff L0_4_L1_0_Wij_reg_Dout_6 (.Q (WindowDout_4__0__6), .QB (\$dummy [46]), .D (
        nx2711), .CLK (CLK)) ;
    ao32 ix2712 (.Y (nx2711), .A0 (Din[6]), .A1 (nx8078), .A2 (WindowWR), .B0 (
         WindowDout_4__0__6), .B1 (nx8200)) ;
    dff L0_4_L1_0_Wij_reg_Dout_7 (.Q (WindowDout_4__0__7), .QB (\$dummy [47]), .D (
        nx2721), .CLK (CLK)) ;
    ao32 ix2722 (.Y (nx2721), .A0 (Din[7]), .A1 (nx8078), .A2 (WindowWR), .B0 (
         WindowDout_4__0__7), .B1 (nx8200)) ;
    oai21 ix2812 (.Y (nx2811), .A0 (nx6181), .A1 (nx7942), .B0 (nx6184)) ;
    dff L0_3_L1_4_Wij_reg_Dout_0 (.Q (WindowDout_3__4__0), .QB (nx6181), .D (
        nx2811), .CLK (CLK)) ;
    nand03 ix6185 (.Y (nx6184), .A0 (nx8078), .A1 (WindowDout_4__4__0), .A2 (
           nx7942)) ;
    oai21 ix2822 (.Y (nx2821), .A0 (nx6188), .A1 (nx7942), .B0 (nx6190)) ;
    dff L0_3_L1_4_Wij_reg_Dout_1 (.Q (WindowDout_3__4__1), .QB (nx6188), .D (
        nx2821), .CLK (CLK)) ;
    nand03 ix6191 (.Y (nx6190), .A0 (nx8078), .A1 (WindowDout_4__4__1), .A2 (
           nx7942)) ;
    oai21 ix2832 (.Y (nx2831), .A0 (nx6194), .A1 (nx7942), .B0 (nx6196)) ;
    dff L0_3_L1_4_Wij_reg_Dout_2 (.Q (WindowDout_3__4__2), .QB (nx6194), .D (
        nx2831), .CLK (CLK)) ;
    nand03 ix6197 (.Y (nx6196), .A0 (nx8078), .A1 (WindowDout_4__4__2), .A2 (
           nx7942)) ;
    oai21 ix2842 (.Y (nx2841), .A0 (nx6200), .A1 (nx7942), .B0 (nx6202)) ;
    dff L0_3_L1_4_Wij_reg_Dout_3 (.Q (WindowDout_3__4__3), .QB (nx6200), .D (
        nx2841), .CLK (CLK)) ;
    nand03 ix6203 (.Y (nx6202), .A0 (nx8080), .A1 (WindowDout_4__4__3), .A2 (
           nx7944)) ;
    oai21 ix2852 (.Y (nx2851), .A0 (nx6206), .A1 (nx7944), .B0 (nx6208)) ;
    dff L0_3_L1_4_Wij_reg_Dout_4 (.Q (WindowDout_3__4__4), .QB (nx6206), .D (
        nx2851), .CLK (CLK)) ;
    nand03 ix6209 (.Y (nx6208), .A0 (nx8080), .A1 (WindowDout_4__4__4), .A2 (
           nx7944)) ;
    oai21 ix2862 (.Y (nx2861), .A0 (nx6212), .A1 (nx7944), .B0 (nx6214)) ;
    dff L0_3_L1_4_Wij_reg_Dout_5 (.Q (WindowDout_3__4__5), .QB (nx6212), .D (
        nx2861), .CLK (CLK)) ;
    nand03 ix6215 (.Y (nx6214), .A0 (nx8080), .A1 (WindowDout_4__4__5), .A2 (
           nx7944)) ;
    oai21 ix2872 (.Y (nx2871), .A0 (nx6218), .A1 (nx7944), .B0 (nx6220)) ;
    dff L0_3_L1_4_Wij_reg_Dout_6 (.Q (WindowDout_3__4__6), .QB (nx6218), .D (
        nx2871), .CLK (CLK)) ;
    nand03 ix6221 (.Y (nx6220), .A0 (nx8080), .A1 (WindowDout_4__4__6), .A2 (
           nx7944)) ;
    oai21 ix2882 (.Y (nx2881), .A0 (nx6224), .A1 (nx7946), .B0 (nx6226)) ;
    dff L0_3_L1_4_Wij_reg_Dout_7 (.Q (WindowDout_3__4__7), .QB (nx6224), .D (
        nx2881), .CLK (CLK)) ;
    nand03 ix6227 (.Y (nx6226), .A0 (nx8080), .A1 (WindowDout_4__4__7), .A2 (
           nx7946)) ;
    oai21 ix2972 (.Y (nx2971), .A0 (nx6230), .A1 (nx7946), .B0 (nx6232)) ;
    dff L0_3_L1_3_Wij_reg_Dout_0 (.Q (WindowDout_3__3__0), .QB (nx6230), .D (
        nx2971), .CLK (CLK)) ;
    nand03 ix6233 (.Y (nx6232), .A0 (nx8080), .A1 (WindowDout_4__3__0), .A2 (
           nx7946)) ;
    oai21 ix2982 (.Y (nx2981), .A0 (nx6236), .A1 (nx7946), .B0 (nx6238)) ;
    dff L0_3_L1_3_Wij_reg_Dout_1 (.Q (WindowDout_3__3__1), .QB (nx6236), .D (
        nx2981), .CLK (CLK)) ;
    nand03 ix6239 (.Y (nx6238), .A0 (nx8080), .A1 (WindowDout_4__3__1), .A2 (
           nx7946)) ;
    oai21 ix2992 (.Y (nx2991), .A0 (nx6242), .A1 (nx7946), .B0 (nx6244)) ;
    dff L0_3_L1_3_Wij_reg_Dout_2 (.Q (WindowDout_3__3__2), .QB (nx6242), .D (
        nx2991), .CLK (CLK)) ;
    nand03 ix6245 (.Y (nx6244), .A0 (nx8082), .A1 (WindowDout_4__3__2), .A2 (
           nx7948)) ;
    oai21 ix3002 (.Y (nx3001), .A0 (nx6248), .A1 (nx7948), .B0 (nx6250)) ;
    dff L0_3_L1_3_Wij_reg_Dout_3 (.Q (WindowDout_3__3__3), .QB (nx6248), .D (
        nx3001), .CLK (CLK)) ;
    nand03 ix6251 (.Y (nx6250), .A0 (nx8082), .A1 (WindowDout_4__3__3), .A2 (
           nx7948)) ;
    oai21 ix3012 (.Y (nx3011), .A0 (nx6254), .A1 (nx7948), .B0 (nx6256)) ;
    dff L0_3_L1_3_Wij_reg_Dout_4 (.Q (WindowDout_3__3__4), .QB (nx6254), .D (
        nx3011), .CLK (CLK)) ;
    nand03 ix6257 (.Y (nx6256), .A0 (nx8082), .A1 (WindowDout_4__3__4), .A2 (
           nx7948)) ;
    oai21 ix3022 (.Y (nx3021), .A0 (nx6260), .A1 (nx7948), .B0 (nx6262)) ;
    dff L0_3_L1_3_Wij_reg_Dout_5 (.Q (WindowDout_3__3__5), .QB (nx6260), .D (
        nx3021), .CLK (CLK)) ;
    nand03 ix6263 (.Y (nx6262), .A0 (nx8082), .A1 (WindowDout_4__3__5), .A2 (
           nx7948)) ;
    oai21 ix3032 (.Y (nx3031), .A0 (nx6266), .A1 (nx7950), .B0 (nx6268)) ;
    dff L0_3_L1_3_Wij_reg_Dout_6 (.Q (WindowDout_3__3__6), .QB (nx6266), .D (
        nx3031), .CLK (CLK)) ;
    nand03 ix6269 (.Y (nx6268), .A0 (nx8082), .A1 (WindowDout_4__3__6), .A2 (
           nx7950)) ;
    oai21 ix3042 (.Y (nx3041), .A0 (nx6272), .A1 (nx7950), .B0 (nx6274)) ;
    dff L0_3_L1_3_Wij_reg_Dout_7 (.Q (WindowDout_3__3__7), .QB (nx6272), .D (
        nx3041), .CLK (CLK)) ;
    nand03 ix6275 (.Y (nx6274), .A0 (nx8082), .A1 (WindowDout_4__3__7), .A2 (
           nx7950)) ;
    dff L0_3_L1_2_Wij_reg_Dout_0 (.Q (WindowDout_3__2__0), .QB (\$dummy [48]), .D (
        nx3131), .CLK (CLK)) ;
    ao32 ix3132 (.Y (nx3131), .A0 (nx8082), .A1 (WindowDout_4__2__0), .A2 (
         WindowWR), .B0 (WindowDout_3__2__0), .B1 (nx8200)) ;
    dff L0_3_L1_2_Wij_reg_Dout_1 (.Q (WindowDout_3__2__1), .QB (\$dummy [49]), .D (
        nx3141), .CLK (CLK)) ;
    ao32 ix3142 (.Y (nx3141), .A0 (nx8084), .A1 (WindowDout_4__2__1), .A2 (
         WindowWR), .B0 (WindowDout_3__2__1), .B1 (nx8200)) ;
    dff L0_3_L1_2_Wij_reg_Dout_2 (.Q (WindowDout_3__2__2), .QB (\$dummy [50]), .D (
        nx3151), .CLK (CLK)) ;
    ao32 ix3152 (.Y (nx3151), .A0 (nx8084), .A1 (WindowDout_4__2__2), .A2 (
         WindowWR), .B0 (WindowDout_3__2__2), .B1 (nx8200)) ;
    dff L0_3_L1_2_Wij_reg_Dout_3 (.Q (WindowDout_3__2__3), .QB (\$dummy [51]), .D (
        nx3161), .CLK (CLK)) ;
    ao32 ix3162 (.Y (nx3161), .A0 (nx8084), .A1 (WindowDout_4__2__3), .A2 (
         WindowWR), .B0 (WindowDout_3__2__3), .B1 (nx8200)) ;
    dff L0_3_L1_2_Wij_reg_Dout_4 (.Q (WindowDout_3__2__4), .QB (\$dummy [52]), .D (
        nx3171), .CLK (CLK)) ;
    ao32 ix3172 (.Y (nx3171), .A0 (nx8084), .A1 (WindowDout_4__2__4), .A2 (
         WindowWR), .B0 (WindowDout_3__2__4), .B1 (nx8202)) ;
    dff L0_3_L1_2_Wij_reg_Dout_5 (.Q (WindowDout_3__2__5), .QB (\$dummy [53]), .D (
        nx3181), .CLK (CLK)) ;
    ao32 ix3182 (.Y (nx3181), .A0 (nx8084), .A1 (WindowDout_4__2__5), .A2 (
         WindowWR), .B0 (WindowDout_3__2__5), .B1 (nx8202)) ;
    dff L0_3_L1_2_Wij_reg_Dout_6 (.Q (WindowDout_3__2__6), .QB (\$dummy [54]), .D (
        nx3191), .CLK (CLK)) ;
    ao32 ix3192 (.Y (nx3191), .A0 (nx8084), .A1 (WindowDout_4__2__6), .A2 (
         WindowWR), .B0 (WindowDout_3__2__6), .B1 (nx8202)) ;
    dff L0_3_L1_2_Wij_reg_Dout_7 (.Q (WindowDout_3__2__7), .QB (\$dummy [55]), .D (
        nx3201), .CLK (CLK)) ;
    ao32 ix3202 (.Y (nx3201), .A0 (nx8084), .A1 (WindowDout_4__2__7), .A2 (
         WindowWR), .B0 (WindowDout_3__2__7), .B1 (nx8202)) ;
    dff L0_3_L1_1_Wij_reg_Dout_0 (.Q (WindowDout_3__1__0), .QB (\$dummy [56]), .D (
        nx3291), .CLK (CLK)) ;
    ao32 ix3292 (.Y (nx3291), .A0 (nx8086), .A1 (WindowDout_4__1__0), .A2 (
         WindowWR), .B0 (WindowDout_3__1__0), .B1 (nx8202)) ;
    dff L0_3_L1_1_Wij_reg_Dout_1 (.Q (WindowDout_3__1__1), .QB (\$dummy [57]), .D (
        nx3301), .CLK (CLK)) ;
    ao32 ix3302 (.Y (nx3301), .A0 (nx8086), .A1 (WindowDout_4__1__1), .A2 (
         WindowWR), .B0 (WindowDout_3__1__1), .B1 (nx8202)) ;
    dff L0_3_L1_1_Wij_reg_Dout_2 (.Q (WindowDout_3__1__2), .QB (\$dummy [58]), .D (
        nx3311), .CLK (CLK)) ;
    ao32 ix3312 (.Y (nx3311), .A0 (nx8086), .A1 (WindowDout_4__1__2), .A2 (
         WindowWR), .B0 (WindowDout_3__1__2), .B1 (nx8202)) ;
    dff L0_3_L1_1_Wij_reg_Dout_3 (.Q (WindowDout_3__1__3), .QB (\$dummy [59]), .D (
        nx3321), .CLK (CLK)) ;
    ao32 ix3322 (.Y (nx3321), .A0 (nx8086), .A1 (WindowDout_4__1__3), .A2 (
         WindowWR), .B0 (WindowDout_3__1__3), .B1 (nx8204)) ;
    dff L0_3_L1_1_Wij_reg_Dout_4 (.Q (WindowDout_3__1__4), .QB (\$dummy [60]), .D (
        nx3331), .CLK (CLK)) ;
    ao32 ix3332 (.Y (nx3331), .A0 (nx8086), .A1 (WindowDout_4__1__4), .A2 (
         WindowWR), .B0 (WindowDout_3__1__4), .B1 (nx8204)) ;
    dff L0_3_L1_1_Wij_reg_Dout_5 (.Q (WindowDout_3__1__5), .QB (\$dummy [61]), .D (
        nx3341), .CLK (CLK)) ;
    ao32 ix3342 (.Y (nx3341), .A0 (nx8086), .A1 (WindowDout_4__1__5), .A2 (
         WindowWR), .B0 (WindowDout_3__1__5), .B1 (nx8204)) ;
    dff L0_3_L1_1_Wij_reg_Dout_6 (.Q (WindowDout_3__1__6), .QB (\$dummy [62]), .D (
        nx3351), .CLK (CLK)) ;
    ao32 ix3352 (.Y (nx3351), .A0 (nx8086), .A1 (WindowDout_4__1__6), .A2 (
         WindowWR), .B0 (WindowDout_3__1__6), .B1 (nx8204)) ;
    dff L0_3_L1_1_Wij_reg_Dout_7 (.Q (WindowDout_3__1__7), .QB (\$dummy [63]), .D (
        nx3361), .CLK (CLK)) ;
    ao32 ix3362 (.Y (nx3361), .A0 (nx8088), .A1 (WindowDout_4__1__7), .A2 (
         WindowWR), .B0 (WindowDout_3__1__7), .B1 (nx8204)) ;
    dff L0_3_L1_0_Wij_reg_Dout_0 (.Q (WindowDout_3__0__0), .QB (\$dummy [64]), .D (
        nx3451), .CLK (CLK)) ;
    ao32 ix3452 (.Y (nx3451), .A0 (nx8088), .A1 (WindowDout_4__0__0), .A2 (
         WindowWR), .B0 (WindowDout_3__0__0), .B1 (nx8204)) ;
    dff L0_3_L1_0_Wij_reg_Dout_1 (.Q (WindowDout_3__0__1), .QB (\$dummy [65]), .D (
        nx3461), .CLK (CLK)) ;
    ao32 ix3462 (.Y (nx3461), .A0 (nx8088), .A1 (WindowDout_4__0__1), .A2 (
         WindowWR), .B0 (WindowDout_3__0__1), .B1 (nx8204)) ;
    dff L0_3_L1_0_Wij_reg_Dout_2 (.Q (WindowDout_3__0__2), .QB (\$dummy [66]), .D (
        nx3471), .CLK (CLK)) ;
    ao32 ix3472 (.Y (nx3471), .A0 (nx8088), .A1 (WindowDout_4__0__2), .A2 (
         WindowWR), .B0 (WindowDout_3__0__2), .B1 (nx8206)) ;
    dff L0_3_L1_0_Wij_reg_Dout_3 (.Q (WindowDout_3__0__3), .QB (\$dummy [67]), .D (
        nx3481), .CLK (CLK)) ;
    ao32 ix3482 (.Y (nx3481), .A0 (nx8088), .A1 (WindowDout_4__0__3), .A2 (
         WindowWR), .B0 (WindowDout_3__0__3), .B1 (nx8206)) ;
    dff L0_3_L1_0_Wij_reg_Dout_4 (.Q (WindowDout_3__0__4), .QB (\$dummy [68]), .D (
        nx3491), .CLK (CLK)) ;
    ao32 ix3492 (.Y (nx3491), .A0 (nx8088), .A1 (WindowDout_4__0__4), .A2 (
         WindowWR), .B0 (WindowDout_3__0__4), .B1 (nx8206)) ;
    dff L0_3_L1_0_Wij_reg_Dout_5 (.Q (WindowDout_3__0__5), .QB (\$dummy [69]), .D (
        nx3501), .CLK (CLK)) ;
    ao32 ix3502 (.Y (nx3501), .A0 (nx8088), .A1 (WindowDout_4__0__5), .A2 (
         WindowWR), .B0 (WindowDout_3__0__5), .B1 (nx8206)) ;
    dff L0_3_L1_0_Wij_reg_Dout_6 (.Q (WindowDout_3__0__6), .QB (\$dummy [70]), .D (
        nx3511), .CLK (CLK)) ;
    ao32 ix3512 (.Y (nx3511), .A0 (nx8090), .A1 (WindowDout_4__0__6), .A2 (
         WindowWR), .B0 (WindowDout_3__0__6), .B1 (nx8206)) ;
    dff L0_3_L1_0_Wij_reg_Dout_7 (.Q (WindowDout_3__0__7), .QB (\$dummy [71]), .D (
        nx3521), .CLK (CLK)) ;
    ao32 ix3522 (.Y (nx3521), .A0 (nx8090), .A1 (WindowDout_4__0__7), .A2 (
         WindowWR), .B0 (WindowDout_3__0__7), .B1 (nx8206)) ;
    oai21 ix3612 (.Y (nx3611), .A0 (nx6350), .A1 (nx7950), .B0 (nx6352)) ;
    dff L0_2_L1_4_Wij_reg_Dout_0 (.Q (WindowDout_2__4__0), .QB (nx6350), .D (
        nx3611), .CLK (CLK)) ;
    oai21 ix3622 (.Y (nx3621), .A0 (nx6356), .A1 (nx7950), .B0 (nx6358)) ;
    dff L0_2_L1_4_Wij_reg_Dout_1 (.Q (WindowDout_2__4__1), .QB (nx6356), .D (
        nx3621), .CLK (CLK)) ;
    oai21 ix3632 (.Y (nx3631), .A0 (nx6362), .A1 (nx7952), .B0 (nx6364)) ;
    dff L0_2_L1_4_Wij_reg_Dout_2 (.Q (WindowDout_2__4__2), .QB (nx6362), .D (
        nx3631), .CLK (CLK)) ;
    oai21 ix3642 (.Y (nx3641), .A0 (nx6368), .A1 (nx7952), .B0 (nx6370)) ;
    dff L0_2_L1_4_Wij_reg_Dout_3 (.Q (WindowDout_2__4__3), .QB (nx6368), .D (
        nx3641), .CLK (CLK)) ;
    oai21 ix3652 (.Y (nx3651), .A0 (nx6374), .A1 (nx7952), .B0 (nx6376)) ;
    dff L0_2_L1_4_Wij_reg_Dout_4 (.Q (WindowDout_2__4__4), .QB (nx6374), .D (
        nx3651), .CLK (CLK)) ;
    oai21 ix3662 (.Y (nx3661), .A0 (nx6380), .A1 (nx7954), .B0 (nx6382)) ;
    dff L0_2_L1_4_Wij_reg_Dout_5 (.Q (WindowDout_2__4__5), .QB (nx6380), .D (
        nx3661), .CLK (CLK)) ;
    oai21 ix3672 (.Y (nx3671), .A0 (nx6386), .A1 (nx7954), .B0 (nx6388)) ;
    dff L0_2_L1_4_Wij_reg_Dout_6 (.Q (WindowDout_2__4__6), .QB (nx6386), .D (
        nx3671), .CLK (CLK)) ;
    oai21 ix3682 (.Y (nx3681), .A0 (nx6392), .A1 (nx7954), .B0 (nx6394)) ;
    dff L0_2_L1_4_Wij_reg_Dout_7 (.Q (WindowDout_2__4__7), .QB (nx6392), .D (
        nx3681), .CLK (CLK)) ;
    oai21 ix3772 (.Y (nx3771), .A0 (nx6398), .A1 (nx7954), .B0 (nx6400)) ;
    dff L0_2_L1_3_Wij_reg_Dout_0 (.Q (WindowDout_2__3__0), .QB (nx6398), .D (
        nx3771), .CLK (CLK)) ;
    oai21 ix3782 (.Y (nx3781), .A0 (nx6404), .A1 (nx7956), .B0 (nx6406)) ;
    dff L0_2_L1_3_Wij_reg_Dout_1 (.Q (WindowDout_2__3__1), .QB (nx6404), .D (
        nx3781), .CLK (CLK)) ;
    oai21 ix3792 (.Y (nx3791), .A0 (nx6410), .A1 (nx7956), .B0 (nx6412)) ;
    dff L0_2_L1_3_Wij_reg_Dout_2 (.Q (WindowDout_2__3__2), .QB (nx6410), .D (
        nx3791), .CLK (CLK)) ;
    oai21 ix3802 (.Y (nx3801), .A0 (nx6416), .A1 (nx7956), .B0 (nx6418)) ;
    dff L0_2_L1_3_Wij_reg_Dout_3 (.Q (WindowDout_2__3__3), .QB (nx6416), .D (
        nx3801), .CLK (CLK)) ;
    oai21 ix3812 (.Y (nx3811), .A0 (nx6422), .A1 (nx7958), .B0 (nx6424)) ;
    dff L0_2_L1_3_Wij_reg_Dout_4 (.Q (WindowDout_2__3__4), .QB (nx6422), .D (
        nx3811), .CLK (CLK)) ;
    oai21 ix3822 (.Y (nx3821), .A0 (nx6428), .A1 (nx7958), .B0 (nx6430)) ;
    dff L0_2_L1_3_Wij_reg_Dout_5 (.Q (WindowDout_2__3__5), .QB (nx6428), .D (
        nx3821), .CLK (CLK)) ;
    oai21 ix3832 (.Y (nx3831), .A0 (nx6434), .A1 (nx7958), .B0 (nx6436)) ;
    dff L0_2_L1_3_Wij_reg_Dout_6 (.Q (WindowDout_2__3__6), .QB (nx6434), .D (
        nx3831), .CLK (CLK)) ;
    oai21 ix3842 (.Y (nx3841), .A0 (nx6440), .A1 (nx7958), .B0 (nx6442)) ;
    dff L0_2_L1_3_Wij_reg_Dout_7 (.Q (WindowDout_2__3__7), .QB (nx6440), .D (
        nx3841), .CLK (CLK)) ;
    dff L0_2_L1_2_Wij_reg_Dout_0 (.Q (WindowDout_2__2__0), .QB (\$dummy [72]), .D (
        nx3931), .CLK (CLK)) ;
    ao32 ix3932 (.Y (nx3931), .A0 (nx8094), .A1 (WindowDout_3__2__0), .A2 (
         WindowWR), .B0 (WindowDout_2__2__0), .B1 (nx8206)) ;
    dff L0_2_L1_2_Wij_reg_Dout_1 (.Q (WindowDout_2__2__1), .QB (\$dummy [73]), .D (
        nx3941), .CLK (CLK)) ;
    ao32 ix3942 (.Y (nx3941), .A0 (nx8094), .A1 (WindowDout_3__2__1), .A2 (
         WindowWR), .B0 (WindowDout_2__2__1), .B1 (nx8208)) ;
    dff L0_2_L1_2_Wij_reg_Dout_2 (.Q (WindowDout_2__2__2), .QB (\$dummy [74]), .D (
        nx3951), .CLK (CLK)) ;
    ao32 ix3952 (.Y (nx3951), .A0 (nx8094), .A1 (WindowDout_3__2__2), .A2 (
         WindowWR), .B0 (WindowDout_2__2__2), .B1 (nx8208)) ;
    dff L0_2_L1_2_Wij_reg_Dout_3 (.Q (WindowDout_2__2__3), .QB (\$dummy [75]), .D (
        nx3961), .CLK (CLK)) ;
    ao32 ix3962 (.Y (nx3961), .A0 (nx8096), .A1 (WindowDout_3__2__3), .A2 (
         WindowWR), .B0 (WindowDout_2__2__3), .B1 (nx8208)) ;
    dff L0_2_L1_2_Wij_reg_Dout_4 (.Q (WindowDout_2__2__4), .QB (\$dummy [76]), .D (
        nx3971), .CLK (CLK)) ;
    ao32 ix3972 (.Y (nx3971), .A0 (nx8096), .A1 (WindowDout_3__2__4), .A2 (
         WindowWR), .B0 (WindowDout_2__2__4), .B1 (nx8208)) ;
    dff L0_2_L1_2_Wij_reg_Dout_5 (.Q (WindowDout_2__2__5), .QB (\$dummy [77]), .D (
        nx3981), .CLK (CLK)) ;
    ao32 ix3982 (.Y (nx3981), .A0 (nx8096), .A1 (WindowDout_3__2__5), .A2 (
         WindowWR), .B0 (WindowDout_2__2__5), .B1 (nx8208)) ;
    dff L0_2_L1_2_Wij_reg_Dout_6 (.Q (WindowDout_2__2__6), .QB (\$dummy [78]), .D (
        nx3991), .CLK (CLK)) ;
    ao32 ix3992 (.Y (nx3991), .A0 (nx8096), .A1 (WindowDout_3__2__6), .A2 (
         WindowWR), .B0 (WindowDout_2__2__6), .B1 (nx8208)) ;
    dff L0_2_L1_2_Wij_reg_Dout_7 (.Q (WindowDout_2__2__7), .QB (\$dummy [79]), .D (
        nx4001), .CLK (CLK)) ;
    ao32 ix4002 (.Y (nx4001), .A0 (nx8096), .A1 (WindowDout_3__2__7), .A2 (
         WindowWR), .B0 (WindowDout_2__2__7), .B1 (nx8208)) ;
    dff L0_2_L1_1_Wij_reg_Dout_0 (.Q (WindowDout_2__1__0), .QB (\$dummy [80]), .D (
        nx4091), .CLK (CLK)) ;
    ao32 ix4092 (.Y (nx4091), .A0 (nx8096), .A1 (WindowDout_3__1__0), .A2 (
         WindowWR), .B0 (WindowDout_2__1__0), .B1 (nx8210)) ;
    dff L0_2_L1_1_Wij_reg_Dout_1 (.Q (WindowDout_2__1__1), .QB (\$dummy [81]), .D (
        nx4101), .CLK (CLK)) ;
    ao32 ix4102 (.Y (nx4101), .A0 (nx8096), .A1 (WindowDout_3__1__1), .A2 (
         WindowWR), .B0 (WindowDout_2__1__1), .B1 (nx8210)) ;
    dff L0_2_L1_1_Wij_reg_Dout_2 (.Q (WindowDout_2__1__2), .QB (\$dummy [82]), .D (
        nx4111), .CLK (CLK)) ;
    ao32 ix4112 (.Y (nx4111), .A0 (nx8098), .A1 (WindowDout_3__1__2), .A2 (
         WindowWR), .B0 (WindowDout_2__1__2), .B1 (nx8210)) ;
    dff L0_2_L1_1_Wij_reg_Dout_3 (.Q (WindowDout_2__1__3), .QB (\$dummy [83]), .D (
        nx4121), .CLK (CLK)) ;
    ao32 ix4122 (.Y (nx4121), .A0 (nx8098), .A1 (WindowDout_3__1__3), .A2 (
         WindowWR), .B0 (WindowDout_2__1__3), .B1 (nx8210)) ;
    dff L0_2_L1_1_Wij_reg_Dout_4 (.Q (WindowDout_2__1__4), .QB (\$dummy [84]), .D (
        nx4131), .CLK (CLK)) ;
    ao32 ix4132 (.Y (nx4131), .A0 (nx8098), .A1 (WindowDout_3__1__4), .A2 (
         WindowWR), .B0 (WindowDout_2__1__4), .B1 (nx8210)) ;
    dff L0_2_L1_1_Wij_reg_Dout_5 (.Q (WindowDout_2__1__5), .QB (\$dummy [85]), .D (
        nx4141), .CLK (CLK)) ;
    ao32 ix4142 (.Y (nx4141), .A0 (nx8098), .A1 (WindowDout_3__1__5), .A2 (
         WindowWR), .B0 (WindowDout_2__1__5), .B1 (nx8210)) ;
    dff L0_2_L1_1_Wij_reg_Dout_6 (.Q (WindowDout_2__1__6), .QB (\$dummy [86]), .D (
        nx4151), .CLK (CLK)) ;
    ao32 ix4152 (.Y (nx4151), .A0 (nx8098), .A1 (WindowDout_3__1__6), .A2 (
         WindowWR), .B0 (WindowDout_2__1__6), .B1 (nx8210)) ;
    dff L0_2_L1_1_Wij_reg_Dout_7 (.Q (WindowDout_2__1__7), .QB (\$dummy [87]), .D (
        nx4161), .CLK (CLK)) ;
    ao32 ix4162 (.Y (nx4161), .A0 (nx8098), .A1 (WindowDout_3__1__7), .A2 (
         WindowWR), .B0 (WindowDout_2__1__7), .B1 (nx8212)) ;
    dff L0_2_L1_0_Wij_reg_Dout_0 (.Q (WindowDout_2__0__0), .QB (\$dummy [88]), .D (
        nx4251), .CLK (CLK)) ;
    ao32 ix4252 (.Y (nx4251), .A0 (nx8098), .A1 (WindowDout_3__0__0), .A2 (
         WindowWR), .B0 (WindowDout_2__0__0), .B1 (nx8212)) ;
    dff L0_2_L1_0_Wij_reg_Dout_1 (.Q (WindowDout_2__0__1), .QB (\$dummy [89]), .D (
        nx4261), .CLK (CLK)) ;
    ao32 ix4262 (.Y (nx4261), .A0 (nx8100), .A1 (WindowDout_3__0__1), .A2 (
         WindowWR), .B0 (WindowDout_2__0__1), .B1 (nx8212)) ;
    dff L0_2_L1_0_Wij_reg_Dout_2 (.Q (WindowDout_2__0__2), .QB (\$dummy [90]), .D (
        nx4271), .CLK (CLK)) ;
    ao32 ix4272 (.Y (nx4271), .A0 (nx8100), .A1 (WindowDout_3__0__2), .A2 (
         WindowWR), .B0 (WindowDout_2__0__2), .B1 (nx8212)) ;
    dff L0_2_L1_0_Wij_reg_Dout_3 (.Q (WindowDout_2__0__3), .QB (\$dummy [91]), .D (
        nx4281), .CLK (CLK)) ;
    ao32 ix4282 (.Y (nx4281), .A0 (nx8100), .A1 (WindowDout_3__0__3), .A2 (
         WindowWR), .B0 (WindowDout_2__0__3), .B1 (nx8212)) ;
    dff L0_2_L1_0_Wij_reg_Dout_4 (.Q (WindowDout_2__0__4), .QB (\$dummy [92]), .D (
        nx4291), .CLK (CLK)) ;
    ao32 ix4292 (.Y (nx4291), .A0 (nx8100), .A1 (WindowDout_3__0__4), .A2 (
         WindowWR), .B0 (WindowDout_2__0__4), .B1 (nx8212)) ;
    dff L0_2_L1_0_Wij_reg_Dout_5 (.Q (WindowDout_2__0__5), .QB (\$dummy [93]), .D (
        nx4301), .CLK (CLK)) ;
    ao32 ix4302 (.Y (nx4301), .A0 (nx8100), .A1 (WindowDout_3__0__5), .A2 (
         WindowWR), .B0 (WindowDout_2__0__5), .B1 (nx8212)) ;
    dff L0_2_L1_0_Wij_reg_Dout_6 (.Q (WindowDout_2__0__6), .QB (\$dummy [94]), .D (
        nx4311), .CLK (CLK)) ;
    ao32 ix4312 (.Y (nx4311), .A0 (nx8100), .A1 (WindowDout_3__0__6), .A2 (
         WindowWR), .B0 (WindowDout_2__0__6), .B1 (nx8214)) ;
    dff L0_2_L1_0_Wij_reg_Dout_7 (.Q (WindowDout_2__0__7), .QB (\$dummy [95]), .D (
        nx4321), .CLK (CLK)) ;
    ao32 ix4322 (.Y (nx4321), .A0 (nx8100), .A1 (WindowDout_3__0__7), .A2 (
         WindowWR), .B0 (WindowDout_2__0__7), .B1 (nx8214)) ;
    oai21 ix4412 (.Y (nx4411), .A0 (nx6518), .A1 (nx7960), .B0 (nx6520)) ;
    dff L0_1_L1_4_Wij_reg_Dout_0 (.Q (WindowDout_1__4__0), .QB (nx6518), .D (
        nx4411), .CLK (CLK)) ;
    oai21 ix4422 (.Y (nx4421), .A0 (nx6524), .A1 (nx7960), .B0 (nx6526)) ;
    dff L0_1_L1_4_Wij_reg_Dout_1 (.Q (WindowDout_1__4__1), .QB (nx6524), .D (
        nx4421), .CLK (CLK)) ;
    oai21 ix4432 (.Y (nx4431), .A0 (nx6530), .A1 (nx7960), .B0 (nx6532)) ;
    dff L0_1_L1_4_Wij_reg_Dout_2 (.Q (WindowDout_1__4__2), .QB (nx6530), .D (
        nx4431), .CLK (CLK)) ;
    oai21 ix4442 (.Y (nx4441), .A0 (nx6536), .A1 (nx7962), .B0 (nx6538)) ;
    dff L0_1_L1_4_Wij_reg_Dout_3 (.Q (WindowDout_1__4__3), .QB (nx6536), .D (
        nx4441), .CLK (CLK)) ;
    oai21 ix4452 (.Y (nx4451), .A0 (nx6542), .A1 (nx7962), .B0 (nx6544)) ;
    dff L0_1_L1_4_Wij_reg_Dout_4 (.Q (WindowDout_1__4__4), .QB (nx6542), .D (
        nx4451), .CLK (CLK)) ;
    oai21 ix4462 (.Y (nx4461), .A0 (nx6548), .A1 (nx7962), .B0 (nx6550)) ;
    dff L0_1_L1_4_Wij_reg_Dout_5 (.Q (WindowDout_1__4__5), .QB (nx6548), .D (
        nx4461), .CLK (CLK)) ;
    oai21 ix4472 (.Y (nx4471), .A0 (nx6554), .A1 (nx7962), .B0 (nx6556)) ;
    dff L0_1_L1_4_Wij_reg_Dout_6 (.Q (WindowDout_1__4__6), .QB (nx6554), .D (
        nx4471), .CLK (CLK)) ;
    oai21 ix4482 (.Y (nx4481), .A0 (nx6560), .A1 (nx7964), .B0 (nx6562)) ;
    dff L0_1_L1_4_Wij_reg_Dout_7 (.Q (WindowDout_1__4__7), .QB (nx6560), .D (
        nx4481), .CLK (CLK)) ;
    oai21 ix4732 (.Y (nx4731), .A0 (nx6566), .A1 (nx7964), .B0 (nx6568)) ;
    dff L0_1_L1_3_Wij_reg_Dout_0 (.Q (WindowDout_1__3__0), .QB (nx6566), .D (
        nx4731), .CLK (CLK)) ;
    oai21 ix4742 (.Y (nx4741), .A0 (nx6572), .A1 (nx7964), .B0 (nx6574)) ;
    dff L0_1_L1_3_Wij_reg_Dout_1 (.Q (WindowDout_1__3__1), .QB (nx6572), .D (
        nx4741), .CLK (CLK)) ;
    oai21 ix4752 (.Y (nx4751), .A0 (nx6578), .A1 (nx7966), .B0 (nx6580)) ;
    dff L0_1_L1_3_Wij_reg_Dout_2 (.Q (WindowDout_1__3__2), .QB (nx6578), .D (
        nx4751), .CLK (CLK)) ;
    oai21 ix4762 (.Y (nx4761), .A0 (nx6584), .A1 (nx7966), .B0 (nx6586)) ;
    dff L0_1_L1_3_Wij_reg_Dout_3 (.Q (WindowDout_1__3__3), .QB (nx6584), .D (
        nx4761), .CLK (CLK)) ;
    oai21 ix4772 (.Y (nx4771), .A0 (nx6590), .A1 (nx7966), .B0 (nx6592)) ;
    dff L0_1_L1_3_Wij_reg_Dout_4 (.Q (WindowDout_1__3__4), .QB (nx6590), .D (
        nx4771), .CLK (CLK)) ;
    oai21 ix4782 (.Y (nx4781), .A0 (nx6596), .A1 (nx7966), .B0 (nx6598)) ;
    dff L0_1_L1_3_Wij_reg_Dout_5 (.Q (WindowDout_1__3__5), .QB (nx6596), .D (
        nx4781), .CLK (CLK)) ;
    oai21 ix4792 (.Y (nx4791), .A0 (nx6602), .A1 (nx7968), .B0 (nx6604)) ;
    dff L0_1_L1_3_Wij_reg_Dout_6 (.Q (WindowDout_1__3__6), .QB (nx6602), .D (
        nx4791), .CLK (CLK)) ;
    oai21 ix4802 (.Y (nx4801), .A0 (nx6608), .A1 (nx7968), .B0 (nx6610)) ;
    dff L0_1_L1_3_Wij_reg_Dout_7 (.Q (WindowDout_1__3__7), .QB (nx6608), .D (
        nx4801), .CLK (CLK)) ;
    oai21 ix5052 (.Y (nx5051), .A0 (nx6614), .A1 (nx7968), .B0 (nx6616)) ;
    dff L0_1_L1_2_Wij_reg_Dout_0 (.Q (WindowDout_1__2__0), .QB (nx6614), .D (
        nx5051), .CLK (CLK)) ;
    nand03 ix6617 (.Y (nx6616), .A0 (nx8106), .A1 (WindowDout_2__2__0), .A2 (
           nx7968)) ;
    oai21 ix5062 (.Y (nx5061), .A0 (nx6620), .A1 (nx7970), .B0 (nx6622)) ;
    dff L0_1_L1_2_Wij_reg_Dout_1 (.Q (WindowDout_1__2__1), .QB (nx6620), .D (
        nx5061), .CLK (CLK)) ;
    nand03 ix6623 (.Y (nx6622), .A0 (nx8106), .A1 (WindowDout_2__2__1), .A2 (
           nx7970)) ;
    oai21 ix5072 (.Y (nx5071), .A0 (nx6626), .A1 (nx7970), .B0 (nx6628)) ;
    dff L0_1_L1_2_Wij_reg_Dout_2 (.Q (WindowDout_1__2__2), .QB (nx6626), .D (
        nx5071), .CLK (CLK)) ;
    nand03 ix6629 (.Y (nx6628), .A0 (nx8106), .A1 (WindowDout_2__2__2), .A2 (
           nx7970)) ;
    oai21 ix5082 (.Y (nx5081), .A0 (nx6632), .A1 (nx7970), .B0 (nx6634)) ;
    dff L0_1_L1_2_Wij_reg_Dout_3 (.Q (WindowDout_1__2__3), .QB (nx6632), .D (
        nx5081), .CLK (CLK)) ;
    nand03 ix6635 (.Y (nx6634), .A0 (nx8106), .A1 (WindowDout_2__2__3), .A2 (
           nx7970)) ;
    oai21 ix5092 (.Y (nx5091), .A0 (nx6638), .A1 (nx7970), .B0 (nx6640)) ;
    dff L0_1_L1_2_Wij_reg_Dout_4 (.Q (WindowDout_1__2__4), .QB (nx6638), .D (
        nx5091), .CLK (CLK)) ;
    nand03 ix6641 (.Y (nx6640), .A0 (nx8106), .A1 (WindowDout_2__2__4), .A2 (
           nx7972)) ;
    oai21 ix5102 (.Y (nx5101), .A0 (nx6644), .A1 (nx7972), .B0 (nx6646)) ;
    dff L0_1_L1_2_Wij_reg_Dout_5 (.Q (WindowDout_1__2__5), .QB (nx6644), .D (
        nx5101), .CLK (CLK)) ;
    nand03 ix6647 (.Y (nx6646), .A0 (nx8108), .A1 (WindowDout_2__2__5), .A2 (
           nx7972)) ;
    oai21 ix5112 (.Y (nx5111), .A0 (nx6650), .A1 (nx7972), .B0 (nx6652)) ;
    dff L0_1_L1_2_Wij_reg_Dout_6 (.Q (WindowDout_1__2__6), .QB (nx6650), .D (
        nx5111), .CLK (CLK)) ;
    nand03 ix6653 (.Y (nx6652), .A0 (nx8108), .A1 (WindowDout_2__2__6), .A2 (
           nx7972)) ;
    oai21 ix5122 (.Y (nx5121), .A0 (nx6656), .A1 (nx7972), .B0 (nx6658)) ;
    dff L0_1_L1_2_Wij_reg_Dout_7 (.Q (WindowDout_1__2__7), .QB (nx6656), .D (
        nx5121), .CLK (CLK)) ;
    nand03 ix6659 (.Y (nx6658), .A0 (nx8108), .A1 (WindowDout_2__2__7), .A2 (
           nx7972)) ;
    oai21 ix5372 (.Y (nx5371), .A0 (nx6662), .A1 (nx7974), .B0 (nx6664)) ;
    dff L0_1_L1_1_Wij_reg_Dout_0 (.Q (WindowDout_1__1__0), .QB (nx6662), .D (
        nx5371), .CLK (CLK)) ;
    nand03 ix6665 (.Y (nx6664), .A0 (nx8108), .A1 (WindowDout_2__1__0), .A2 (
           nx7974)) ;
    oai21 ix5382 (.Y (nx5381), .A0 (nx6668), .A1 (nx7974), .B0 (nx6670)) ;
    dff L0_1_L1_1_Wij_reg_Dout_1 (.Q (WindowDout_1__1__1), .QB (nx6668), .D (
        nx5381), .CLK (CLK)) ;
    nand03 ix6671 (.Y (nx6670), .A0 (nx8108), .A1 (WindowDout_2__1__1), .A2 (
           nx7974)) ;
    oai21 ix5392 (.Y (nx5391), .A0 (nx6674), .A1 (nx7974), .B0 (nx6676)) ;
    dff L0_1_L1_1_Wij_reg_Dout_2 (.Q (WindowDout_1__1__2), .QB (nx6674), .D (
        nx5391), .CLK (CLK)) ;
    nand03 ix6677 (.Y (nx6676), .A0 (nx8108), .A1 (WindowDout_2__1__2), .A2 (
           nx7974)) ;
    oai21 ix5402 (.Y (nx5401), .A0 (nx6680), .A1 (nx7974), .B0 (nx6682)) ;
    dff L0_1_L1_1_Wij_reg_Dout_3 (.Q (WindowDout_1__1__3), .QB (nx6680), .D (
        nx5401), .CLK (CLK)) ;
    nand03 ix6683 (.Y (nx6682), .A0 (nx8108), .A1 (WindowDout_2__1__3), .A2 (
           nx7976)) ;
    oai21 ix5412 (.Y (nx5411), .A0 (nx6686), .A1 (nx7976), .B0 (nx6688)) ;
    dff L0_1_L1_1_Wij_reg_Dout_4 (.Q (WindowDout_1__1__4), .QB (nx6686), .D (
        nx5411), .CLK (CLK)) ;
    nand03 ix6689 (.Y (nx6688), .A0 (nx8110), .A1 (WindowDout_2__1__4), .A2 (
           nx7976)) ;
    oai21 ix5422 (.Y (nx5421), .A0 (nx6692), .A1 (nx7976), .B0 (nx6694)) ;
    dff L0_1_L1_1_Wij_reg_Dout_5 (.Q (WindowDout_1__1__5), .QB (nx6692), .D (
        nx5421), .CLK (CLK)) ;
    nand03 ix6695 (.Y (nx6694), .A0 (nx8110), .A1 (WindowDout_2__1__5), .A2 (
           nx7976)) ;
    oai21 ix5432 (.Y (nx5431), .A0 (nx6698), .A1 (nx7976), .B0 (nx6700)) ;
    dff L0_1_L1_1_Wij_reg_Dout_6 (.Q (WindowDout_1__1__6), .QB (nx6698), .D (
        nx5431), .CLK (CLK)) ;
    nand03 ix6701 (.Y (nx6700), .A0 (nx8110), .A1 (WindowDout_2__1__6), .A2 (
           nx7976)) ;
    oai21 ix5442 (.Y (nx5441), .A0 (nx6704), .A1 (nx7978), .B0 (nx6706)) ;
    dff L0_1_L1_1_Wij_reg_Dout_7 (.Q (WindowDout_1__1__7), .QB (nx6704), .D (
        nx5441), .CLK (CLK)) ;
    nand03 ix6707 (.Y (nx6706), .A0 (nx8110), .A1 (WindowDout_2__1__7), .A2 (
           nx7978)) ;
    oai21 ix5692 (.Y (nx5691), .A0 (nx6710), .A1 (nx7978), .B0 (nx6712)) ;
    dff L0_1_L1_0_Wij_reg_Dout_0 (.Q (WindowDout_1__0__0), .QB (nx6710), .D (
        nx5691), .CLK (CLK)) ;
    nand03 ix6713 (.Y (nx6712), .A0 (nx8110), .A1 (WindowDout_2__0__0), .A2 (
           nx7978)) ;
    oai21 ix5702 (.Y (nx5701), .A0 (nx6716), .A1 (nx7978), .B0 (nx6718)) ;
    dff L0_1_L1_0_Wij_reg_Dout_1 (.Q (WindowDout_1__0__1), .QB (nx6716), .D (
        nx5701), .CLK (CLK)) ;
    nand03 ix6719 (.Y (nx6718), .A0 (nx8110), .A1 (WindowDout_2__0__1), .A2 (
           nx7978)) ;
    oai21 ix5712 (.Y (nx5711), .A0 (nx6722), .A1 (nx7978), .B0 (nx6724)) ;
    dff L0_1_L1_0_Wij_reg_Dout_2 (.Q (WindowDout_1__0__2), .QB (nx6722), .D (
        nx5711), .CLK (CLK)) ;
    nand03 ix6725 (.Y (nx6724), .A0 (nx8110), .A1 (WindowDout_2__0__2), .A2 (
           nx7980)) ;
    oai21 ix5722 (.Y (nx5721), .A0 (nx6728), .A1 (nx7980), .B0 (nx6730)) ;
    dff L0_1_L1_0_Wij_reg_Dout_3 (.Q (WindowDout_1__0__3), .QB (nx6728), .D (
        nx5721), .CLK (CLK)) ;
    nand03 ix6731 (.Y (nx6730), .A0 (nx8112), .A1 (WindowDout_2__0__3), .A2 (
           nx7980)) ;
    oai21 ix5732 (.Y (nx5731), .A0 (nx6734), .A1 (nx7980), .B0 (nx6736)) ;
    dff L0_1_L1_0_Wij_reg_Dout_4 (.Q (WindowDout_1__0__4), .QB (nx6734), .D (
        nx5731), .CLK (CLK)) ;
    nand03 ix6737 (.Y (nx6736), .A0 (nx8112), .A1 (WindowDout_2__0__4), .A2 (
           nx7980)) ;
    oai21 ix5742 (.Y (nx5741), .A0 (nx6740), .A1 (nx7980), .B0 (nx6742)) ;
    dff L0_1_L1_0_Wij_reg_Dout_5 (.Q (WindowDout_1__0__5), .QB (nx6740), .D (
        nx5741), .CLK (CLK)) ;
    nand03 ix6743 (.Y (nx6742), .A0 (nx8112), .A1 (WindowDout_2__0__5), .A2 (
           nx7980)) ;
    oai21 ix5752 (.Y (nx5751), .A0 (nx6746), .A1 (nx7982), .B0 (nx6748)) ;
    dff L0_1_L1_0_Wij_reg_Dout_6 (.Q (WindowDout_1__0__6), .QB (nx6746), .D (
        nx5751), .CLK (CLK)) ;
    nand03 ix6749 (.Y (nx6748), .A0 (nx8112), .A1 (WindowDout_2__0__6), .A2 (
           nx7982)) ;
    oai21 ix5762 (.Y (nx5761), .A0 (nx6752), .A1 (nx7982), .B0 (nx6754)) ;
    dff L0_1_L1_0_Wij_reg_Dout_7 (.Q (WindowDout_1__0__7), .QB (nx6752), .D (
        nx5761), .CLK (CLK)) ;
    nand03 ix6755 (.Y (nx6754), .A0 (nx8112), .A1 (WindowDout_2__0__7), .A2 (
           nx7982)) ;
    oai21 ix4492 (.Y (nx4491), .A0 (nx6758), .A1 (nx7982), .B0 (nx6760)) ;
    dff L0_0_L1_4_Wij_reg_Dout_0 (.Q (WindowDout_0__4__0), .QB (nx6758), .D (
        nx4491), .CLK (CLK)) ;
    oai21 ix4502 (.Y (nx4501), .A0 (nx6764), .A1 (nx7982), .B0 (nx6766)) ;
    dff L0_0_L1_4_Wij_reg_Dout_1 (.Q (WindowDout_0__4__1), .QB (nx6764), .D (
        nx4501), .CLK (CLK)) ;
    oai21 ix4512 (.Y (nx4511), .A0 (nx6770), .A1 (nx7984), .B0 (nx6772)) ;
    dff L0_0_L1_4_Wij_reg_Dout_2 (.Q (WindowDout_0__4__2), .QB (nx6770), .D (
        nx4511), .CLK (CLK)) ;
    oai21 ix4522 (.Y (nx4521), .A0 (nx6776), .A1 (nx7984), .B0 (nx6778)) ;
    dff L0_0_L1_4_Wij_reg_Dout_3 (.Q (WindowDout_0__4__3), .QB (nx6776), .D (
        nx4521), .CLK (CLK)) ;
    oai21 ix4532 (.Y (nx4531), .A0 (nx6782), .A1 (nx7984), .B0 (nx6784)) ;
    dff L0_0_L1_4_Wij_reg_Dout_4 (.Q (WindowDout_0__4__4), .QB (nx6782), .D (
        nx4531), .CLK (CLK)) ;
    oai21 ix4542 (.Y (nx4541), .A0 (nx6788), .A1 (nx7986), .B0 (nx6790)) ;
    dff L0_0_L1_4_Wij_reg_Dout_5 (.Q (WindowDout_0__4__5), .QB (nx6788), .D (
        nx4541), .CLK (CLK)) ;
    oai21 ix4552 (.Y (nx4551), .A0 (nx6794), .A1 (nx7986), .B0 (nx6796)) ;
    dff L0_0_L1_4_Wij_reg_Dout_6 (.Q (WindowDout_0__4__6), .QB (nx6794), .D (
        nx4551), .CLK (CLK)) ;
    oai21 ix4562 (.Y (nx4561), .A0 (nx6800), .A1 (nx7986), .B0 (nx6802)) ;
    dff L0_0_L1_4_Wij_reg_Dout_7 (.Q (WindowDout_0__4__7), .QB (nx6800), .D (
        nx4561), .CLK (CLK)) ;
    oai21 ix4812 (.Y (nx4811), .A0 (nx6806), .A1 (nx7986), .B0 (nx6808)) ;
    dff L0_0_L1_3_Wij_reg_Dout_0 (.Q (WindowDout_0__3__0), .QB (nx6806), .D (
        nx4811), .CLK (CLK)) ;
    oai21 ix4822 (.Y (nx4821), .A0 (nx6812), .A1 (nx7988), .B0 (nx6814)) ;
    dff L0_0_L1_3_Wij_reg_Dout_1 (.Q (WindowDout_0__3__1), .QB (nx6812), .D (
        nx4821), .CLK (CLK)) ;
    oai21 ix4832 (.Y (nx4831), .A0 (nx6818), .A1 (nx7988), .B0 (nx6820)) ;
    dff L0_0_L1_3_Wij_reg_Dout_2 (.Q (WindowDout_0__3__2), .QB (nx6818), .D (
        nx4831), .CLK (CLK)) ;
    oai21 ix4842 (.Y (nx4841), .A0 (nx6824), .A1 (nx7988), .B0 (nx6826)) ;
    dff L0_0_L1_3_Wij_reg_Dout_3 (.Q (WindowDout_0__3__3), .QB (nx6824), .D (
        nx4841), .CLK (CLK)) ;
    oai21 ix4852 (.Y (nx4851), .A0 (nx6830), .A1 (nx7990), .B0 (nx6832)) ;
    dff L0_0_L1_3_Wij_reg_Dout_4 (.Q (WindowDout_0__3__4), .QB (nx6830), .D (
        nx4851), .CLK (CLK)) ;
    oai21 ix4862 (.Y (nx4861), .A0 (nx6836), .A1 (nx7990), .B0 (nx6838)) ;
    dff L0_0_L1_3_Wij_reg_Dout_5 (.Q (WindowDout_0__3__5), .QB (nx6836), .D (
        nx4861), .CLK (CLK)) ;
    oai21 ix4872 (.Y (nx4871), .A0 (nx6842), .A1 (nx7990), .B0 (nx6844)) ;
    dff L0_0_L1_3_Wij_reg_Dout_6 (.Q (WindowDout_0__3__6), .QB (nx6842), .D (
        nx4871), .CLK (CLK)) ;
    oai21 ix4882 (.Y (nx4881), .A0 (nx6848), .A1 (nx7990), .B0 (nx6850)) ;
    dff L0_0_L1_3_Wij_reg_Dout_7 (.Q (WindowDout_0__3__7), .QB (nx6848), .D (
        nx4881), .CLK (CLK)) ;
    oai21 ix5132 (.Y (nx5131), .A0 (nx6854), .A1 (nx7992), .B0 (nx6856)) ;
    dff L0_0_L1_2_Wij_reg_Dout_0 (.Q (WindowDout_0__2__0), .QB (nx6854), .D (
        nx5131), .CLK (CLK)) ;
    oai21 ix5142 (.Y (nx5141), .A0 (nx6860), .A1 (nx7992), .B0 (nx6862)) ;
    dff L0_0_L1_2_Wij_reg_Dout_1 (.Q (WindowDout_0__2__1), .QB (nx6860), .D (
        nx5141), .CLK (CLK)) ;
    oai21 ix5152 (.Y (nx5151), .A0 (nx6866), .A1 (nx7992), .B0 (nx6868)) ;
    dff L0_0_L1_2_Wij_reg_Dout_2 (.Q (WindowDout_0__2__2), .QB (nx6866), .D (
        nx5151), .CLK (CLK)) ;
    oai21 ix5162 (.Y (nx5161), .A0 (nx6872), .A1 (nx7994), .B0 (nx6874)) ;
    dff L0_0_L1_2_Wij_reg_Dout_3 (.Q (WindowDout_0__2__3), .QB (nx6872), .D (
        nx5161), .CLK (CLK)) ;
    oai21 ix5172 (.Y (nx5171), .A0 (nx6878), .A1 (nx7994), .B0 (nx6880)) ;
    dff L0_0_L1_2_Wij_reg_Dout_4 (.Q (WindowDout_0__2__4), .QB (nx6878), .D (
        nx5171), .CLK (CLK)) ;
    oai21 ix5182 (.Y (nx5181), .A0 (nx6884), .A1 (nx7994), .B0 (nx6886)) ;
    dff L0_0_L1_2_Wij_reg_Dout_5 (.Q (WindowDout_0__2__5), .QB (nx6884), .D (
        nx5181), .CLK (CLK)) ;
    oai21 ix5192 (.Y (nx5191), .A0 (nx6890), .A1 (nx7994), .B0 (nx6892)) ;
    dff L0_0_L1_2_Wij_reg_Dout_6 (.Q (WindowDout_0__2__6), .QB (nx6890), .D (
        nx5191), .CLK (CLK)) ;
    oai21 ix5202 (.Y (nx5201), .A0 (nx6896), .A1 (nx7996), .B0 (nx6898)) ;
    dff L0_0_L1_2_Wij_reg_Dout_7 (.Q (WindowDout_0__2__7), .QB (nx6896), .D (
        nx5201), .CLK (CLK)) ;
    oai21 ix5452 (.Y (nx5451), .A0 (nx6902), .A1 (nx7996), .B0 (nx6904)) ;
    dff L0_0_L1_1_Wij_reg_Dout_0 (.Q (WindowDout_0__1__0), .QB (nx6902), .D (
        nx5451), .CLK (CLK)) ;
    oai21 ix5462 (.Y (nx5461), .A0 (nx6908), .A1 (nx7996), .B0 (nx6910)) ;
    dff L0_0_L1_1_Wij_reg_Dout_1 (.Q (WindowDout_0__1__1), .QB (nx6908), .D (
        nx5461), .CLK (CLK)) ;
    oai21 ix5472 (.Y (nx5471), .A0 (nx6914), .A1 (nx7998), .B0 (nx6916)) ;
    dff L0_0_L1_1_Wij_reg_Dout_2 (.Q (WindowDout_0__1__2), .QB (nx6914), .D (
        nx5471), .CLK (CLK)) ;
    oai21 ix5482 (.Y (nx5481), .A0 (nx6920), .A1 (nx7998), .B0 (nx6922)) ;
    dff L0_0_L1_1_Wij_reg_Dout_3 (.Q (WindowDout_0__1__3), .QB (nx6920), .D (
        nx5481), .CLK (CLK)) ;
    oai21 ix5492 (.Y (nx5491), .A0 (nx6926), .A1 (nx7998), .B0 (nx6928)) ;
    dff L0_0_L1_1_Wij_reg_Dout_4 (.Q (WindowDout_0__1__4), .QB (nx6926), .D (
        nx5491), .CLK (CLK)) ;
    oai21 ix5502 (.Y (nx5501), .A0 (nx6932), .A1 (nx7998), .B0 (nx6934)) ;
    dff L0_0_L1_1_Wij_reg_Dout_5 (.Q (WindowDout_0__1__5), .QB (nx6932), .D (
        nx5501), .CLK (CLK)) ;
    oai21 ix5512 (.Y (nx5511), .A0 (nx6938), .A1 (nx8000), .B0 (nx6940)) ;
    dff L0_0_L1_1_Wij_reg_Dout_6 (.Q (WindowDout_0__1__6), .QB (nx6938), .D (
        nx5511), .CLK (CLK)) ;
    oai21 ix5522 (.Y (nx5521), .A0 (nx6944), .A1 (nx8000), .B0 (nx6946)) ;
    dff L0_0_L1_1_Wij_reg_Dout_7 (.Q (WindowDout_0__1__7), .QB (nx6944), .D (
        nx5521), .CLK (CLK)) ;
    oai21 ix5772 (.Y (nx5771), .A0 (nx6950), .A1 (nx8000), .B0 (nx6952)) ;
    dff L0_0_L1_0_Wij_reg_Dout_0 (.Q (WindowDout_0__0__0), .QB (nx6950), .D (
        nx5771), .CLK (CLK)) ;
    oai21 ix5782 (.Y (nx5781), .A0 (nx6956), .A1 (nx8002), .B0 (nx6958)) ;
    dff L0_0_L1_0_Wij_reg_Dout_1 (.Q (WindowDout_0__0__1), .QB (nx6956), .D (
        nx5781), .CLK (CLK)) ;
    oai21 ix5792 (.Y (nx5791), .A0 (nx6962), .A1 (nx8002), .B0 (nx6964)) ;
    dff L0_0_L1_0_Wij_reg_Dout_2 (.Q (WindowDout_0__0__2), .QB (nx6962), .D (
        nx5791), .CLK (CLK)) ;
    oai21 ix5802 (.Y (nx5801), .A0 (nx6968), .A1 (nx8002), .B0 (nx6970)) ;
    dff L0_0_L1_0_Wij_reg_Dout_3 (.Q (WindowDout_0__0__3), .QB (nx6968), .D (
        nx5801), .CLK (CLK)) ;
    oai21 ix5812 (.Y (nx5811), .A0 (nx6974), .A1 (nx8002), .B0 (nx6976)) ;
    dff L0_0_L1_0_Wij_reg_Dout_4 (.Q (WindowDout_0__0__4), .QB (nx6974), .D (
        nx5811), .CLK (CLK)) ;
    oai21 ix5822 (.Y (nx5821), .A0 (nx6980), .A1 (nx8004), .B0 (nx6982)) ;
    dff L0_0_L1_0_Wij_reg_Dout_5 (.Q (WindowDout_0__0__5), .QB (nx6980), .D (
        nx5821), .CLK (CLK)) ;
    oai21 ix5832 (.Y (nx5831), .A0 (nx6986), .A1 (nx8004), .B0 (nx6988)) ;
    dff L0_0_L1_0_Wij_reg_Dout_6 (.Q (WindowDout_0__0__6), .QB (nx6986), .D (
        nx5831), .CLK (CLK)) ;
    oai21 ix5842 (.Y (nx5841), .A0 (nx6992), .A1 (nx8004), .B0 (nx6994)) ;
    dff L0_0_L1_0_Wij_reg_Dout_7 (.Q (WindowDout_0__0__7), .QB (nx6992), .D (
        nx5841), .CLK (CLK)) ;
    dff L0_4_L1_4_Fij_reg_Dout_0 (.Q (FilterDout_4__4__0), .QB (\$dummy [96]), .D (
        nx2091), .CLK (CLK)) ;
    aoi21 ix6999 (.Y (nx6998), .A0 (FilterSize), .A1 (FilterWR), .B0 (RST)) ;
    dff L0_4_L1_4_Fij_reg_Dout_1 (.Q (FilterDout_4__4__1), .QB (\$dummy [97]), .D (
        nx2101), .CLK (CLK)) ;
    dff L0_4_L1_4_Fij_reg_Dout_2 (.Q (FilterDout_4__4__2), .QB (\$dummy [98]), .D (
        nx2111), .CLK (CLK)) ;
    dff L0_4_L1_4_Fij_reg_Dout_3 (.Q (FilterDout_4__4__3), .QB (\$dummy [99]), .D (
        nx2121), .CLK (CLK)) ;
    dff L0_4_L1_4_Fij_reg_Dout_4 (.Q (FilterDout_4__4__4), .QB (\$dummy [100]), 
        .D (nx2131), .CLK (CLK)) ;
    dff L0_4_L1_4_Fij_reg_Dout_5 (.Q (FilterDout_4__4__5), .QB (\$dummy [101]), 
        .D (nx2141), .CLK (CLK)) ;
    dff L0_4_L1_4_Fij_reg_Dout_6 (.Q (FilterDout_4__4__6), .QB (\$dummy [102]), 
        .D (nx2151), .CLK (CLK)) ;
    dff L0_4_L1_4_Fij_reg_Dout_7 (.Q (FilterDout_4__4__7), .QB (\$dummy [103]), 
        .D (nx2161), .CLK (CLK)) ;
    dff L0_4_L1_3_Fij_reg_Dout_0 (.Q (FilterDout_4__3__0), .QB (\$dummy [104]), 
        .D (nx2251), .CLK (CLK)) ;
    dff L0_4_L1_3_Fij_reg_Dout_1 (.Q (FilterDout_4__3__1), .QB (\$dummy [105]), 
        .D (nx2261), .CLK (CLK)) ;
    dff L0_4_L1_3_Fij_reg_Dout_2 (.Q (FilterDout_4__3__2), .QB (\$dummy [106]), 
        .D (nx2271), .CLK (CLK)) ;
    dff L0_4_L1_3_Fij_reg_Dout_3 (.Q (FilterDout_4__3__3), .QB (\$dummy [107]), 
        .D (nx2281), .CLK (CLK)) ;
    dff L0_4_L1_3_Fij_reg_Dout_4 (.Q (FilterDout_4__3__4), .QB (\$dummy [108]), 
        .D (nx2291), .CLK (CLK)) ;
    dff L0_4_L1_3_Fij_reg_Dout_5 (.Q (FilterDout_4__3__5), .QB (\$dummy [109]), 
        .D (nx2301), .CLK (CLK)) ;
    dff L0_4_L1_3_Fij_reg_Dout_6 (.Q (FilterDout_4__3__6), .QB (\$dummy [110]), 
        .D (nx2311), .CLK (CLK)) ;
    dff L0_4_L1_3_Fij_reg_Dout_7 (.Q (FilterDout_4__3__7), .QB (\$dummy [111]), 
        .D (nx2321), .CLK (CLK)) ;
    dff L0_4_L1_2_Fij_reg_Dout_0 (.Q (FilterDout_4__2__0), .QB (\$dummy [112]), 
        .D (nx2411), .CLK (CLK)) ;
    ao32 ix2412 (.Y (nx2411), .A0 (Din[16]), .A1 (nx8124), .A2 (FilterWR), .B0 (
         FilterDout_4__2__0), .B1 (nx8232)) ;
    nor02_2x ix7049 (.Y (nx7048), .A0 (FilterWR), .A1 (RST)) ;
    dff L0_4_L1_2_Fij_reg_Dout_1 (.Q (FilterDout_4__2__1), .QB (\$dummy [113]), 
        .D (nx2421), .CLK (CLK)) ;
    ao32 ix2422 (.Y (nx2421), .A0 (Din[17]), .A1 (nx8124), .A2 (FilterWR), .B0 (
         FilterDout_4__2__1), .B1 (nx8232)) ;
    dff L0_4_L1_2_Fij_reg_Dout_2 (.Q (FilterDout_4__2__2), .QB (\$dummy [114]), 
        .D (nx2431), .CLK (CLK)) ;
    ao32 ix2432 (.Y (nx2431), .A0 (Din[18]), .A1 (nx8124), .A2 (FilterWR), .B0 (
         FilterDout_4__2__2), .B1 (nx8232)) ;
    dff L0_4_L1_2_Fij_reg_Dout_3 (.Q (FilterDout_4__2__3), .QB (\$dummy [115]), 
        .D (nx2441), .CLK (CLK)) ;
    ao32 ix2442 (.Y (nx2441), .A0 (Din[19]), .A1 (nx8124), .A2 (FilterWR), .B0 (
         FilterDout_4__2__3), .B1 (nx8232)) ;
    dff L0_4_L1_2_Fij_reg_Dout_4 (.Q (FilterDout_4__2__4), .QB (\$dummy [116]), 
        .D (nx2451), .CLK (CLK)) ;
    ao32 ix2452 (.Y (nx2451), .A0 (Din[20]), .A1 (nx8126), .A2 (FilterWR), .B0 (
         FilterDout_4__2__4), .B1 (nx8232)) ;
    dff L0_4_L1_2_Fij_reg_Dout_5 (.Q (FilterDout_4__2__5), .QB (\$dummy [117]), 
        .D (nx2461), .CLK (CLK)) ;
    ao32 ix2462 (.Y (nx2461), .A0 (Din[21]), .A1 (nx8126), .A2 (FilterWR), .B0 (
         FilterDout_4__2__5), .B1 (nx8232)) ;
    dff L0_4_L1_2_Fij_reg_Dout_6 (.Q (FilterDout_4__2__6), .QB (\$dummy [118]), 
        .D (nx2471), .CLK (CLK)) ;
    ao32 ix2472 (.Y (nx2471), .A0 (Din[22]), .A1 (nx8126), .A2 (FilterWR), .B0 (
         FilterDout_4__2__6), .B1 (nx8232)) ;
    dff L0_4_L1_2_Fij_reg_Dout_7 (.Q (FilterDout_4__2__7), .QB (\$dummy [119]), 
        .D (nx2481), .CLK (CLK)) ;
    ao32 ix2482 (.Y (nx2481), .A0 (Din[23]), .A1 (nx8126), .A2 (FilterWR), .B0 (
         FilterDout_4__2__7), .B1 (nx8234)) ;
    dff L0_4_L1_1_Fij_reg_Dout_0 (.Q (FilterDout_4__1__0), .QB (\$dummy [120]), 
        .D (nx2571), .CLK (CLK)) ;
    ao32 ix2572 (.Y (nx2571), .A0 (Din[8]), .A1 (nx8126), .A2 (FilterWR), .B0 (
         FilterDout_4__1__0), .B1 (nx8234)) ;
    dff L0_4_L1_1_Fij_reg_Dout_1 (.Q (FilterDout_4__1__1), .QB (\$dummy [121]), 
        .D (nx2581), .CLK (CLK)) ;
    ao32 ix2582 (.Y (nx2581), .A0 (Din[9]), .A1 (nx8126), .A2 (FilterWR), .B0 (
         FilterDout_4__1__1), .B1 (nx8234)) ;
    dff L0_4_L1_1_Fij_reg_Dout_2 (.Q (FilterDout_4__1__2), .QB (\$dummy [122]), 
        .D (nx2591), .CLK (CLK)) ;
    ao32 ix2592 (.Y (nx2591), .A0 (Din[10]), .A1 (nx8126), .A2 (FilterWR), .B0 (
         FilterDout_4__1__2), .B1 (nx8234)) ;
    dff L0_4_L1_1_Fij_reg_Dout_3 (.Q (FilterDout_4__1__3), .QB (\$dummy [123]), 
        .D (nx2601), .CLK (CLK)) ;
    ao32 ix2602 (.Y (nx2601), .A0 (Din[11]), .A1 (nx8128), .A2 (FilterWR), .B0 (
         FilterDout_4__1__3), .B1 (nx8234)) ;
    dff L0_4_L1_1_Fij_reg_Dout_4 (.Q (FilterDout_4__1__4), .QB (\$dummy [124]), 
        .D (nx2611), .CLK (CLK)) ;
    ao32 ix2612 (.Y (nx2611), .A0 (Din[12]), .A1 (nx8128), .A2 (FilterWR), .B0 (
         FilterDout_4__1__4), .B1 (nx8234)) ;
    dff L0_4_L1_1_Fij_reg_Dout_5 (.Q (FilterDout_4__1__5), .QB (\$dummy [125]), 
        .D (nx2621), .CLK (CLK)) ;
    ao32 ix2622 (.Y (nx2621), .A0 (Din[13]), .A1 (nx8128), .A2 (FilterWR), .B0 (
         FilterDout_4__1__5), .B1 (nx8234)) ;
    dff L0_4_L1_1_Fij_reg_Dout_6 (.Q (FilterDout_4__1__6), .QB (\$dummy [126]), 
        .D (nx2631), .CLK (CLK)) ;
    ao32 ix2632 (.Y (nx2631), .A0 (Din[14]), .A1 (nx8128), .A2 (FilterWR), .B0 (
         FilterDout_4__1__6), .B1 (nx8236)) ;
    dff L0_4_L1_1_Fij_reg_Dout_7 (.Q (FilterDout_4__1__7), .QB (\$dummy [127]), 
        .D (nx2641), .CLK (CLK)) ;
    ao32 ix2642 (.Y (nx2641), .A0 (Din[15]), .A1 (nx8128), .A2 (FilterWR), .B0 (
         FilterDout_4__1__7), .B1 (nx8236)) ;
    dff L0_4_L1_0_Fij_reg_Dout_0 (.Q (FilterDout_4__0__0), .QB (\$dummy [128]), 
        .D (nx2731), .CLK (CLK)) ;
    ao32 ix2732 (.Y (nx2731), .A0 (Din[0]), .A1 (nx8128), .A2 (FilterWR), .B0 (
         FilterDout_4__0__0), .B1 (nx8236)) ;
    dff L0_4_L1_0_Fij_reg_Dout_1 (.Q (FilterDout_4__0__1), .QB (\$dummy [129]), 
        .D (nx2741), .CLK (CLK)) ;
    ao32 ix2742 (.Y (nx2741), .A0 (Din[1]), .A1 (nx8128), .A2 (FilterWR), .B0 (
         FilterDout_4__0__1), .B1 (nx8236)) ;
    dff L0_4_L1_0_Fij_reg_Dout_2 (.Q (FilterDout_4__0__2), .QB (\$dummy [130]), 
        .D (nx2751), .CLK (CLK)) ;
    ao32 ix2752 (.Y (nx2751), .A0 (Din[2]), .A1 (nx8130), .A2 (FilterWR), .B0 (
         FilterDout_4__0__2), .B1 (nx8236)) ;
    dff L0_4_L1_0_Fij_reg_Dout_3 (.Q (FilterDout_4__0__3), .QB (\$dummy [131]), 
        .D (nx2761), .CLK (CLK)) ;
    ao32 ix2762 (.Y (nx2761), .A0 (Din[3]), .A1 (nx8130), .A2 (FilterWR), .B0 (
         FilterDout_4__0__3), .B1 (nx8236)) ;
    dff L0_4_L1_0_Fij_reg_Dout_4 (.Q (FilterDout_4__0__4), .QB (\$dummy [132]), 
        .D (nx2771), .CLK (CLK)) ;
    ao32 ix2772 (.Y (nx2771), .A0 (Din[4]), .A1 (nx8130), .A2 (FilterWR), .B0 (
         FilterDout_4__0__4), .B1 (nx8236)) ;
    dff L0_4_L1_0_Fij_reg_Dout_5 (.Q (FilterDout_4__0__5), .QB (\$dummy [133]), 
        .D (nx2781), .CLK (CLK)) ;
    ao32 ix2782 (.Y (nx2781), .A0 (Din[5]), .A1 (nx8130), .A2 (FilterWR), .B0 (
         FilterDout_4__0__5), .B1 (nx8238)) ;
    dff L0_4_L1_0_Fij_reg_Dout_6 (.Q (FilterDout_4__0__6), .QB (\$dummy [134]), 
        .D (nx2791), .CLK (CLK)) ;
    ao32 ix2792 (.Y (nx2791), .A0 (Din[6]), .A1 (nx8130), .A2 (FilterWR), .B0 (
         FilterDout_4__0__6), .B1 (nx8238)) ;
    dff L0_4_L1_0_Fij_reg_Dout_7 (.Q (FilterDout_4__0__7), .QB (\$dummy [135]), 
        .D (nx2801), .CLK (CLK)) ;
    ao32 ix2802 (.Y (nx2801), .A0 (Din[7]), .A1 (nx8130), .A2 (FilterWR), .B0 (
         FilterDout_4__0__7), .B1 (nx8238)) ;
    oai21 ix2892 (.Y (nx2891), .A0 (nx7122), .A1 (nx8006), .B0 (nx7125)) ;
    dff L0_3_L1_4_Fij_reg_Dout_0 (.Q (FilterDout_3__4__0), .QB (nx7122), .D (
        nx2891), .CLK (CLK)) ;
    nand03 ix7126 (.Y (nx7125), .A0 (nx8130), .A1 (FilterDout_4__4__0), .A2 (
           nx8006)) ;
    oai21 ix2902 (.Y (nx2901), .A0 (nx7129), .A1 (nx8006), .B0 (nx7131)) ;
    dff L0_3_L1_4_Fij_reg_Dout_1 (.Q (FilterDout_3__4__1), .QB (nx7129), .D (
        nx2901), .CLK (CLK)) ;
    nand03 ix7132 (.Y (nx7131), .A0 (nx8132), .A1 (FilterDout_4__4__1), .A2 (
           nx8006)) ;
    oai21 ix2912 (.Y (nx2911), .A0 (nx7135), .A1 (nx8006), .B0 (nx7137)) ;
    dff L0_3_L1_4_Fij_reg_Dout_2 (.Q (FilterDout_3__4__2), .QB (nx7135), .D (
        nx2911), .CLK (CLK)) ;
    nand03 ix7138 (.Y (nx7137), .A0 (nx8132), .A1 (FilterDout_4__4__2), .A2 (
           nx8006)) ;
    oai21 ix2922 (.Y (nx2921), .A0 (nx7141), .A1 (nx8006), .B0 (nx7143)) ;
    dff L0_3_L1_4_Fij_reg_Dout_3 (.Q (FilterDout_3__4__3), .QB (nx7141), .D (
        nx2921), .CLK (CLK)) ;
    nand03 ix7144 (.Y (nx7143), .A0 (nx8132), .A1 (FilterDout_4__4__3), .A2 (
           nx8008)) ;
    oai21 ix2932 (.Y (nx2931), .A0 (nx7147), .A1 (nx8008), .B0 (nx7149)) ;
    dff L0_3_L1_4_Fij_reg_Dout_4 (.Q (FilterDout_3__4__4), .QB (nx7147), .D (
        nx2931), .CLK (CLK)) ;
    nand03 ix7150 (.Y (nx7149), .A0 (nx8132), .A1 (FilterDout_4__4__4), .A2 (
           nx8008)) ;
    oai21 ix2942 (.Y (nx2941), .A0 (nx7153), .A1 (nx8008), .B0 (nx7155)) ;
    dff L0_3_L1_4_Fij_reg_Dout_5 (.Q (FilterDout_3__4__5), .QB (nx7153), .D (
        nx2941), .CLK (CLK)) ;
    nand03 ix7156 (.Y (nx7155), .A0 (nx8132), .A1 (FilterDout_4__4__5), .A2 (
           nx8008)) ;
    oai21 ix2952 (.Y (nx2951), .A0 (nx7159), .A1 (nx8008), .B0 (nx7161)) ;
    dff L0_3_L1_4_Fij_reg_Dout_6 (.Q (FilterDout_3__4__6), .QB (nx7159), .D (
        nx2951), .CLK (CLK)) ;
    nand03 ix7162 (.Y (nx7161), .A0 (nx8132), .A1 (FilterDout_4__4__6), .A2 (
           nx8008)) ;
    oai21 ix2962 (.Y (nx2961), .A0 (nx7165), .A1 (nx8010), .B0 (nx7167)) ;
    dff L0_3_L1_4_Fij_reg_Dout_7 (.Q (FilterDout_3__4__7), .QB (nx7165), .D (
        nx2961), .CLK (CLK)) ;
    nand03 ix7168 (.Y (nx7167), .A0 (nx8132), .A1 (FilterDout_4__4__7), .A2 (
           nx8010)) ;
    oai21 ix3052 (.Y (nx3051), .A0 (nx7171), .A1 (nx8010), .B0 (nx7173)) ;
    dff L0_3_L1_3_Fij_reg_Dout_0 (.Q (FilterDout_3__3__0), .QB (nx7171), .D (
        nx3051), .CLK (CLK)) ;
    nand03 ix7174 (.Y (nx7173), .A0 (nx8134), .A1 (FilterDout_4__3__0), .A2 (
           nx8010)) ;
    oai21 ix3062 (.Y (nx3061), .A0 (nx7177), .A1 (nx8010), .B0 (nx7179)) ;
    dff L0_3_L1_3_Fij_reg_Dout_1 (.Q (FilterDout_3__3__1), .QB (nx7177), .D (
        nx3061), .CLK (CLK)) ;
    nand03 ix7180 (.Y (nx7179), .A0 (nx8134), .A1 (FilterDout_4__3__1), .A2 (
           nx8010)) ;
    oai21 ix3072 (.Y (nx3071), .A0 (nx7183), .A1 (nx8010), .B0 (nx7185)) ;
    dff L0_3_L1_3_Fij_reg_Dout_2 (.Q (FilterDout_3__3__2), .QB (nx7183), .D (
        nx3071), .CLK (CLK)) ;
    nand03 ix7186 (.Y (nx7185), .A0 (nx8134), .A1 (FilterDout_4__3__2), .A2 (
           nx8012)) ;
    oai21 ix3082 (.Y (nx3081), .A0 (nx7189), .A1 (nx8012), .B0 (nx7191)) ;
    dff L0_3_L1_3_Fij_reg_Dout_3 (.Q (FilterDout_3__3__3), .QB (nx7189), .D (
        nx3081), .CLK (CLK)) ;
    nand03 ix7192 (.Y (nx7191), .A0 (nx8134), .A1 (FilterDout_4__3__3), .A2 (
           nx8012)) ;
    oai21 ix3092 (.Y (nx3091), .A0 (nx7195), .A1 (nx8012), .B0 (nx7197)) ;
    dff L0_3_L1_3_Fij_reg_Dout_4 (.Q (FilterDout_3__3__4), .QB (nx7195), .D (
        nx3091), .CLK (CLK)) ;
    nand03 ix7198 (.Y (nx7197), .A0 (nx8134), .A1 (FilterDout_4__3__4), .A2 (
           nx8012)) ;
    oai21 ix3102 (.Y (nx3101), .A0 (nx7201), .A1 (nx8012), .B0 (nx7203)) ;
    dff L0_3_L1_3_Fij_reg_Dout_5 (.Q (FilterDout_3__3__5), .QB (nx7201), .D (
        nx3101), .CLK (CLK)) ;
    nand03 ix7204 (.Y (nx7203), .A0 (nx8134), .A1 (FilterDout_4__3__5), .A2 (
           nx8012)) ;
    oai21 ix3112 (.Y (nx3111), .A0 (nx7207), .A1 (nx8014), .B0 (nx7209)) ;
    dff L0_3_L1_3_Fij_reg_Dout_6 (.Q (FilterDout_3__3__6), .QB (nx7207), .D (
        nx3111), .CLK (CLK)) ;
    nand03 ix7210 (.Y (nx7209), .A0 (nx8134), .A1 (FilterDout_4__3__6), .A2 (
           nx8014)) ;
    oai21 ix3122 (.Y (nx3121), .A0 (nx7213), .A1 (nx8014), .B0 (nx7215)) ;
    dff L0_3_L1_3_Fij_reg_Dout_7 (.Q (FilterDout_3__3__7), .QB (nx7213), .D (
        nx3121), .CLK (CLK)) ;
    nand03 ix7216 (.Y (nx7215), .A0 (nx8136), .A1 (FilterDout_4__3__7), .A2 (
           nx8014)) ;
    dff L0_3_L1_2_Fij_reg_Dout_0 (.Q (FilterDout_3__2__0), .QB (\$dummy [136]), 
        .D (nx3211), .CLK (CLK)) ;
    ao32 ix3212 (.Y (nx3211), .A0 (nx8136), .A1 (FilterDout_4__2__0), .A2 (
         FilterWR), .B0 (FilterDout_3__2__0), .B1 (nx8238)) ;
    dff L0_3_L1_2_Fij_reg_Dout_1 (.Q (FilterDout_3__2__1), .QB (\$dummy [137]), 
        .D (nx3221), .CLK (CLK)) ;
    ao32 ix3222 (.Y (nx3221), .A0 (nx8136), .A1 (FilterDout_4__2__1), .A2 (
         FilterWR), .B0 (FilterDout_3__2__1), .B1 (nx8238)) ;
    dff L0_3_L1_2_Fij_reg_Dout_2 (.Q (FilterDout_3__2__2), .QB (\$dummy [138]), 
        .D (nx3231), .CLK (CLK)) ;
    ao32 ix3232 (.Y (nx3231), .A0 (nx8136), .A1 (FilterDout_4__2__2), .A2 (
         FilterWR), .B0 (FilterDout_3__2__2), .B1 (nx8238)) ;
    dff L0_3_L1_2_Fij_reg_Dout_3 (.Q (FilterDout_3__2__3), .QB (\$dummy [139]), 
        .D (nx3241), .CLK (CLK)) ;
    ao32 ix3242 (.Y (nx3241), .A0 (nx8136), .A1 (FilterDout_4__2__3), .A2 (
         FilterWR), .B0 (FilterDout_3__2__3), .B1 (nx8238)) ;
    dff L0_3_L1_2_Fij_reg_Dout_4 (.Q (FilterDout_3__2__4), .QB (\$dummy [140]), 
        .D (nx3251), .CLK (CLK)) ;
    ao32 ix3252 (.Y (nx3251), .A0 (nx8136), .A1 (FilterDout_4__2__4), .A2 (
         FilterWR), .B0 (FilterDout_3__2__4), .B1 (nx8240)) ;
    dff L0_3_L1_2_Fij_reg_Dout_5 (.Q (FilterDout_3__2__5), .QB (\$dummy [141]), 
        .D (nx3261), .CLK (CLK)) ;
    ao32 ix3262 (.Y (nx3261), .A0 (nx8136), .A1 (FilterDout_4__2__5), .A2 (
         FilterWR), .B0 (FilterDout_3__2__5), .B1 (nx8240)) ;
    dff L0_3_L1_2_Fij_reg_Dout_6 (.Q (FilterDout_3__2__6), .QB (\$dummy [142]), 
        .D (nx3271), .CLK (CLK)) ;
    ao32 ix3272 (.Y (nx3271), .A0 (nx8138), .A1 (FilterDout_4__2__6), .A2 (
         FilterWR), .B0 (FilterDout_3__2__6), .B1 (nx8240)) ;
    dff L0_3_L1_2_Fij_reg_Dout_7 (.Q (FilterDout_3__2__7), .QB (\$dummy [143]), 
        .D (nx3281), .CLK (CLK)) ;
    ao32 ix3282 (.Y (nx3281), .A0 (nx8138), .A1 (FilterDout_4__2__7), .A2 (
         FilterWR), .B0 (FilterDout_3__2__7), .B1 (nx8240)) ;
    dff L0_3_L1_1_Fij_reg_Dout_0 (.Q (FilterDout_3__1__0), .QB (\$dummy [144]), 
        .D (nx3371), .CLK (CLK)) ;
    ao32 ix3372 (.Y (nx3371), .A0 (nx8138), .A1 (FilterDout_4__1__0), .A2 (
         FilterWR), .B0 (FilterDout_3__1__0), .B1 (nx8240)) ;
    dff L0_3_L1_1_Fij_reg_Dout_1 (.Q (FilterDout_3__1__1), .QB (\$dummy [145]), 
        .D (nx3381), .CLK (CLK)) ;
    ao32 ix3382 (.Y (nx3381), .A0 (nx8138), .A1 (FilterDout_4__1__1), .A2 (
         FilterWR), .B0 (FilterDout_3__1__1), .B1 (nx8240)) ;
    dff L0_3_L1_1_Fij_reg_Dout_2 (.Q (FilterDout_3__1__2), .QB (\$dummy [146]), 
        .D (nx3391), .CLK (CLK)) ;
    ao32 ix3392 (.Y (nx3391), .A0 (nx8138), .A1 (FilterDout_4__1__2), .A2 (
         FilterWR), .B0 (FilterDout_3__1__2), .B1 (nx8240)) ;
    dff L0_3_L1_1_Fij_reg_Dout_3 (.Q (FilterDout_3__1__3), .QB (\$dummy [147]), 
        .D (nx3401), .CLK (CLK)) ;
    ao32 ix3402 (.Y (nx3401), .A0 (nx8138), .A1 (FilterDout_4__1__3), .A2 (
         FilterWR), .B0 (FilterDout_3__1__3), .B1 (nx8242)) ;
    dff L0_3_L1_1_Fij_reg_Dout_4 (.Q (FilterDout_3__1__4), .QB (\$dummy [148]), 
        .D (nx3411), .CLK (CLK)) ;
    ao32 ix3412 (.Y (nx3411), .A0 (nx8138), .A1 (FilterDout_4__1__4), .A2 (
         FilterWR), .B0 (FilterDout_3__1__4), .B1 (nx8242)) ;
    dff L0_3_L1_1_Fij_reg_Dout_5 (.Q (FilterDout_3__1__5), .QB (\$dummy [149]), 
        .D (nx3421), .CLK (CLK)) ;
    ao32 ix3422 (.Y (nx3421), .A0 (nx8140), .A1 (FilterDout_4__1__5), .A2 (
         FilterWR), .B0 (FilterDout_3__1__5), .B1 (nx8242)) ;
    dff L0_3_L1_1_Fij_reg_Dout_6 (.Q (FilterDout_3__1__6), .QB (\$dummy [150]), 
        .D (nx3431), .CLK (CLK)) ;
    ao32 ix3432 (.Y (nx3431), .A0 (nx8140), .A1 (FilterDout_4__1__6), .A2 (
         FilterWR), .B0 (FilterDout_3__1__6), .B1 (nx8242)) ;
    dff L0_3_L1_1_Fij_reg_Dout_7 (.Q (FilterDout_3__1__7), .QB (\$dummy [151]), 
        .D (nx3441), .CLK (CLK)) ;
    ao32 ix3442 (.Y (nx3441), .A0 (nx8140), .A1 (FilterDout_4__1__7), .A2 (
         FilterWR), .B0 (FilterDout_3__1__7), .B1 (nx8242)) ;
    dff L0_3_L1_0_Fij_reg_Dout_0 (.Q (FilterDout_3__0__0), .QB (\$dummy [152]), 
        .D (nx3531), .CLK (CLK)) ;
    ao32 ix3532 (.Y (nx3531), .A0 (nx8140), .A1 (FilterDout_4__0__0), .A2 (
         FilterWR), .B0 (FilterDout_3__0__0), .B1 (nx8242)) ;
    dff L0_3_L1_0_Fij_reg_Dout_1 (.Q (FilterDout_3__0__1), .QB (\$dummy [153]), 
        .D (nx3541), .CLK (CLK)) ;
    ao32 ix3542 (.Y (nx3541), .A0 (nx8140), .A1 (FilterDout_4__0__1), .A2 (
         FilterWR), .B0 (FilterDout_3__0__1), .B1 (nx8242)) ;
    dff L0_3_L1_0_Fij_reg_Dout_2 (.Q (FilterDout_3__0__2), .QB (\$dummy [154]), 
        .D (nx3551), .CLK (CLK)) ;
    ao32 ix3552 (.Y (nx3551), .A0 (nx8140), .A1 (FilterDout_4__0__2), .A2 (
         FilterWR), .B0 (FilterDout_3__0__2), .B1 (nx8244)) ;
    dff L0_3_L1_0_Fij_reg_Dout_3 (.Q (FilterDout_3__0__3), .QB (\$dummy [155]), 
        .D (nx3561), .CLK (CLK)) ;
    ao32 ix3562 (.Y (nx3561), .A0 (nx8140), .A1 (FilterDout_4__0__3), .A2 (
         FilterWR), .B0 (FilterDout_3__0__3), .B1 (nx8244)) ;
    dff L0_3_L1_0_Fij_reg_Dout_4 (.Q (FilterDout_3__0__4), .QB (\$dummy [156]), 
        .D (nx3571), .CLK (CLK)) ;
    ao32 ix3572 (.Y (nx3571), .A0 (nx8142), .A1 (FilterDout_4__0__4), .A2 (
         FilterWR), .B0 (FilterDout_3__0__4), .B1 (nx8244)) ;
    dff L0_3_L1_0_Fij_reg_Dout_5 (.Q (FilterDout_3__0__5), .QB (\$dummy [157]), 
        .D (nx3581), .CLK (CLK)) ;
    ao32 ix3582 (.Y (nx3581), .A0 (nx8142), .A1 (FilterDout_4__0__5), .A2 (
         FilterWR), .B0 (FilterDout_3__0__5), .B1 (nx8244)) ;
    dff L0_3_L1_0_Fij_reg_Dout_6 (.Q (FilterDout_3__0__6), .QB (\$dummy [158]), 
        .D (nx3591), .CLK (CLK)) ;
    ao32 ix3592 (.Y (nx3591), .A0 (nx8142), .A1 (FilterDout_4__0__6), .A2 (
         FilterWR), .B0 (FilterDout_3__0__6), .B1 (nx8244)) ;
    dff L0_3_L1_0_Fij_reg_Dout_7 (.Q (FilterDout_3__0__7), .QB (\$dummy [159]), 
        .D (nx3601), .CLK (CLK)) ;
    ao32 ix3602 (.Y (nx3601), .A0 (nx8142), .A1 (FilterDout_4__0__7), .A2 (
         FilterWR), .B0 (FilterDout_3__0__7), .B1 (nx8244)) ;
    oai21 ix3692 (.Y (nx3691), .A0 (nx7291), .A1 (nx8014), .B0 (nx7293)) ;
    dff L0_2_L1_4_Fij_reg_Dout_0 (.Q (FilterDout_2__4__0), .QB (nx7291), .D (
        nx3691), .CLK (CLK)) ;
    oai21 ix3702 (.Y (nx3701), .A0 (nx7297), .A1 (nx8014), .B0 (nx7299)) ;
    dff L0_2_L1_4_Fij_reg_Dout_1 (.Q (FilterDout_2__4__1), .QB (nx7297), .D (
        nx3701), .CLK (CLK)) ;
    oai21 ix3712 (.Y (nx3711), .A0 (nx7303), .A1 (nx8016), .B0 (nx7305)) ;
    dff L0_2_L1_4_Fij_reg_Dout_2 (.Q (FilterDout_2__4__2), .QB (nx7303), .D (
        nx3711), .CLK (CLK)) ;
    oai21 ix3722 (.Y (nx3721), .A0 (nx7309), .A1 (nx8016), .B0 (nx7311)) ;
    dff L0_2_L1_4_Fij_reg_Dout_3 (.Q (FilterDout_2__4__3), .QB (nx7309), .D (
        nx3721), .CLK (CLK)) ;
    oai21 ix3732 (.Y (nx3731), .A0 (nx7315), .A1 (nx8016), .B0 (nx7317)) ;
    dff L0_2_L1_4_Fij_reg_Dout_4 (.Q (FilterDout_2__4__4), .QB (nx7315), .D (
        nx3731), .CLK (CLK)) ;
    oai21 ix3742 (.Y (nx3741), .A0 (nx7321), .A1 (nx8018), .B0 (nx7323)) ;
    dff L0_2_L1_4_Fij_reg_Dout_5 (.Q (FilterDout_2__4__5), .QB (nx7321), .D (
        nx3741), .CLK (CLK)) ;
    oai21 ix3752 (.Y (nx3751), .A0 (nx7327), .A1 (nx8018), .B0 (nx7329)) ;
    dff L0_2_L1_4_Fij_reg_Dout_6 (.Q (FilterDout_2__4__6), .QB (nx7327), .D (
        nx3751), .CLK (CLK)) ;
    oai21 ix3762 (.Y (nx3761), .A0 (nx7333), .A1 (nx8018), .B0 (nx7335)) ;
    dff L0_2_L1_4_Fij_reg_Dout_7 (.Q (FilterDout_2__4__7), .QB (nx7333), .D (
        nx3761), .CLK (CLK)) ;
    oai21 ix3852 (.Y (nx3851), .A0 (nx7339), .A1 (nx8018), .B0 (nx7341)) ;
    dff L0_2_L1_3_Fij_reg_Dout_0 (.Q (FilterDout_2__3__0), .QB (nx7339), .D (
        nx3851), .CLK (CLK)) ;
    oai21 ix3862 (.Y (nx3861), .A0 (nx7345), .A1 (nx8020), .B0 (nx7347)) ;
    dff L0_2_L1_3_Fij_reg_Dout_1 (.Q (FilterDout_2__3__1), .QB (nx7345), .D (
        nx3861), .CLK (CLK)) ;
    oai21 ix3872 (.Y (nx3871), .A0 (nx7351), .A1 (nx8020), .B0 (nx7353)) ;
    dff L0_2_L1_3_Fij_reg_Dout_2 (.Q (FilterDout_2__3__2), .QB (nx7351), .D (
        nx3871), .CLK (CLK)) ;
    oai21 ix3882 (.Y (nx3881), .A0 (nx7357), .A1 (nx8020), .B0 (nx7359)) ;
    dff L0_2_L1_3_Fij_reg_Dout_3 (.Q (FilterDout_2__3__3), .QB (nx7357), .D (
        nx3881), .CLK (CLK)) ;
    oai21 ix3892 (.Y (nx3891), .A0 (nx7363), .A1 (nx8022), .B0 (nx7365)) ;
    dff L0_2_L1_3_Fij_reg_Dout_4 (.Q (FilterDout_2__3__4), .QB (nx7363), .D (
        nx3891), .CLK (CLK)) ;
    oai21 ix3902 (.Y (nx3901), .A0 (nx7369), .A1 (nx8022), .B0 (nx7371)) ;
    dff L0_2_L1_3_Fij_reg_Dout_5 (.Q (FilterDout_2__3__5), .QB (nx7369), .D (
        nx3901), .CLK (CLK)) ;
    oai21 ix3912 (.Y (nx3911), .A0 (nx7375), .A1 (nx8022), .B0 (nx7377)) ;
    dff L0_2_L1_3_Fij_reg_Dout_6 (.Q (FilterDout_2__3__6), .QB (nx7375), .D (
        nx3911), .CLK (CLK)) ;
    oai21 ix3922 (.Y (nx3921), .A0 (nx7381), .A1 (nx8022), .B0 (nx7383)) ;
    dff L0_2_L1_3_Fij_reg_Dout_7 (.Q (FilterDout_2__3__7), .QB (nx7381), .D (
        nx3921), .CLK (CLK)) ;
    dff L0_2_L1_2_Fij_reg_Dout_0 (.Q (FilterDout_2__2__0), .QB (\$dummy [160]), 
        .D (nx4011), .CLK (CLK)) ;
    ao32 ix4012 (.Y (nx4011), .A0 (nx8146), .A1 (FilterDout_3__2__0), .A2 (
         FilterWR), .B0 (FilterDout_2__2__0), .B1 (nx8244)) ;
    dff L0_2_L1_2_Fij_reg_Dout_1 (.Q (FilterDout_2__2__1), .QB (\$dummy [161]), 
        .D (nx4021), .CLK (CLK)) ;
    ao32 ix4022 (.Y (nx4021), .A0 (nx8148), .A1 (FilterDout_3__2__1), .A2 (
         FilterWR), .B0 (FilterDout_2__2__1), .B1 (nx8246)) ;
    dff L0_2_L1_2_Fij_reg_Dout_2 (.Q (FilterDout_2__2__2), .QB (\$dummy [162]), 
        .D (nx4031), .CLK (CLK)) ;
    ao32 ix4032 (.Y (nx4031), .A0 (nx8148), .A1 (FilterDout_3__2__2), .A2 (
         FilterWR), .B0 (FilterDout_2__2__2), .B1 (nx8246)) ;
    dff L0_2_L1_2_Fij_reg_Dout_3 (.Q (FilterDout_2__2__3), .QB (\$dummy [163]), 
        .D (nx4041), .CLK (CLK)) ;
    ao32 ix4042 (.Y (nx4041), .A0 (nx8148), .A1 (FilterDout_3__2__3), .A2 (
         FilterWR), .B0 (FilterDout_2__2__3), .B1 (nx8246)) ;
    dff L0_2_L1_2_Fij_reg_Dout_4 (.Q (FilterDout_2__2__4), .QB (\$dummy [164]), 
        .D (nx4051), .CLK (CLK)) ;
    ao32 ix4052 (.Y (nx4051), .A0 (nx8148), .A1 (FilterDout_3__2__4), .A2 (
         FilterWR), .B0 (FilterDout_2__2__4), .B1 (nx8246)) ;
    dff L0_2_L1_2_Fij_reg_Dout_5 (.Q (FilterDout_2__2__5), .QB (\$dummy [165]), 
        .D (nx4061), .CLK (CLK)) ;
    ao32 ix4062 (.Y (nx4061), .A0 (nx8148), .A1 (FilterDout_3__2__5), .A2 (
         FilterWR), .B0 (FilterDout_2__2__5), .B1 (nx8246)) ;
    dff L0_2_L1_2_Fij_reg_Dout_6 (.Q (FilterDout_2__2__6), .QB (\$dummy [166]), 
        .D (nx4071), .CLK (CLK)) ;
    ao32 ix4072 (.Y (nx4071), .A0 (nx8148), .A1 (FilterDout_3__2__6), .A2 (
         FilterWR), .B0 (FilterDout_2__2__6), .B1 (nx8246)) ;
    dff L0_2_L1_2_Fij_reg_Dout_7 (.Q (FilterDout_2__2__7), .QB (\$dummy [167]), 
        .D (nx4081), .CLK (CLK)) ;
    ao32 ix4082 (.Y (nx4081), .A0 (nx8148), .A1 (FilterDout_3__2__7), .A2 (
         FilterWR), .B0 (FilterDout_2__2__7), .B1 (nx8246)) ;
    dff L0_2_L1_1_Fij_reg_Dout_0 (.Q (FilterDout_2__1__0), .QB (\$dummy [168]), 
        .D (nx4171), .CLK (CLK)) ;
    ao32 ix4172 (.Y (nx4171), .A0 (nx8150), .A1 (FilterDout_3__1__0), .A2 (
         FilterWR), .B0 (FilterDout_2__1__0), .B1 (nx8248)) ;
    dff L0_2_L1_1_Fij_reg_Dout_1 (.Q (FilterDout_2__1__1), .QB (\$dummy [169]), 
        .D (nx4181), .CLK (CLK)) ;
    ao32 ix4182 (.Y (nx4181), .A0 (nx8150), .A1 (FilterDout_3__1__1), .A2 (
         FilterWR), .B0 (FilterDout_2__1__1), .B1 (nx8248)) ;
    dff L0_2_L1_1_Fij_reg_Dout_2 (.Q (FilterDout_2__1__2), .QB (\$dummy [170]), 
        .D (nx4191), .CLK (CLK)) ;
    ao32 ix4192 (.Y (nx4191), .A0 (nx8150), .A1 (FilterDout_3__1__2), .A2 (
         FilterWR), .B0 (FilterDout_2__1__2), .B1 (nx8248)) ;
    dff L0_2_L1_1_Fij_reg_Dout_3 (.Q (FilterDout_2__1__3), .QB (\$dummy [171]), 
        .D (nx4201), .CLK (CLK)) ;
    ao32 ix4202 (.Y (nx4201), .A0 (nx8150), .A1 (FilterDout_3__1__3), .A2 (
         FilterWR), .B0 (FilterDout_2__1__3), .B1 (nx8248)) ;
    dff L0_2_L1_1_Fij_reg_Dout_4 (.Q (FilterDout_2__1__4), .QB (\$dummy [172]), 
        .D (nx4211), .CLK (CLK)) ;
    ao32 ix4212 (.Y (nx4211), .A0 (nx8150), .A1 (FilterDout_3__1__4), .A2 (
         FilterWR), .B0 (FilterDout_2__1__4), .B1 (nx8248)) ;
    dff L0_2_L1_1_Fij_reg_Dout_5 (.Q (FilterDout_2__1__5), .QB (\$dummy [173]), 
        .D (nx4221), .CLK (CLK)) ;
    ao32 ix4222 (.Y (nx4221), .A0 (nx8150), .A1 (FilterDout_3__1__5), .A2 (
         FilterWR), .B0 (FilterDout_2__1__5), .B1 (nx8248)) ;
    dff L0_2_L1_1_Fij_reg_Dout_6 (.Q (FilterDout_2__1__6), .QB (\$dummy [174]), 
        .D (nx4231), .CLK (CLK)) ;
    ao32 ix4232 (.Y (nx4231), .A0 (nx8150), .A1 (FilterDout_3__1__6), .A2 (
         FilterWR), .B0 (FilterDout_2__1__6), .B1 (nx8248)) ;
    dff L0_2_L1_1_Fij_reg_Dout_7 (.Q (FilterDout_2__1__7), .QB (\$dummy [175]), 
        .D (nx4241), .CLK (CLK)) ;
    ao32 ix4242 (.Y (nx4241), .A0 (nx8152), .A1 (FilterDout_3__1__7), .A2 (
         FilterWR), .B0 (FilterDout_2__1__7), .B1 (nx8250)) ;
    dff L0_2_L1_0_Fij_reg_Dout_0 (.Q (FilterDout_2__0__0), .QB (\$dummy [176]), 
        .D (nx4331), .CLK (CLK)) ;
    ao32 ix4332 (.Y (nx4331), .A0 (nx8152), .A1 (FilterDout_3__0__0), .A2 (
         FilterWR), .B0 (FilterDout_2__0__0), .B1 (nx8250)) ;
    dff L0_2_L1_0_Fij_reg_Dout_1 (.Q (FilterDout_2__0__1), .QB (\$dummy [177]), 
        .D (nx4341), .CLK (CLK)) ;
    ao32 ix4342 (.Y (nx4341), .A0 (nx8152), .A1 (FilterDout_3__0__1), .A2 (
         FilterWR), .B0 (FilterDout_2__0__1), .B1 (nx8250)) ;
    dff L0_2_L1_0_Fij_reg_Dout_2 (.Q (FilterDout_2__0__2), .QB (\$dummy [178]), 
        .D (nx4351), .CLK (CLK)) ;
    ao32 ix4352 (.Y (nx4351), .A0 (nx8152), .A1 (FilterDout_3__0__2), .A2 (
         FilterWR), .B0 (FilterDout_2__0__2), .B1 (nx8250)) ;
    dff L0_2_L1_0_Fij_reg_Dout_3 (.Q (FilterDout_2__0__3), .QB (\$dummy [179]), 
        .D (nx4361), .CLK (CLK)) ;
    ao32 ix4362 (.Y (nx4361), .A0 (nx8152), .A1 (FilterDout_3__0__3), .A2 (
         FilterWR), .B0 (FilterDout_2__0__3), .B1 (nx8250)) ;
    dff L0_2_L1_0_Fij_reg_Dout_4 (.Q (FilterDout_2__0__4), .QB (\$dummy [180]), 
        .D (nx4371), .CLK (CLK)) ;
    ao32 ix4372 (.Y (nx4371), .A0 (nx8152), .A1 (FilterDout_3__0__4), .A2 (
         FilterWR), .B0 (FilterDout_2__0__4), .B1 (nx8250)) ;
    dff L0_2_L1_0_Fij_reg_Dout_5 (.Q (FilterDout_2__0__5), .QB (\$dummy [181]), 
        .D (nx4381), .CLK (CLK)) ;
    ao32 ix4382 (.Y (nx4381), .A0 (nx8152), .A1 (FilterDout_3__0__5), .A2 (
         FilterWR), .B0 (FilterDout_2__0__5), .B1 (nx8250)) ;
    dff L0_2_L1_0_Fij_reg_Dout_6 (.Q (FilterDout_2__0__6), .QB (\$dummy [182]), 
        .D (nx4391), .CLK (CLK)) ;
    ao32 ix4392 (.Y (nx4391), .A0 (nx8154), .A1 (FilterDout_3__0__6), .A2 (
         FilterWR), .B0 (FilterDout_2__0__6), .B1 (nx8252)) ;
    dff L0_2_L1_0_Fij_reg_Dout_7 (.Q (FilterDout_2__0__7), .QB (\$dummy [183]), 
        .D (nx4401), .CLK (CLK)) ;
    ao32 ix4402 (.Y (nx4401), .A0 (nx8154), .A1 (FilterDout_3__0__7), .A2 (
         FilterWR), .B0 (FilterDout_2__0__7), .B1 (nx8252)) ;
    oai21 ix4572 (.Y (nx4571), .A0 (nx7459), .A1 (nx8024), .B0 (nx7461)) ;
    dff L0_1_L1_4_Fij_reg_Dout_0 (.Q (FilterDout_1__4__0), .QB (nx7459), .D (
        nx4571), .CLK (CLK)) ;
    oai21 ix4582 (.Y (nx4581), .A0 (nx7465), .A1 (nx8024), .B0 (nx7467)) ;
    dff L0_1_L1_4_Fij_reg_Dout_1 (.Q (FilterDout_1__4__1), .QB (nx7465), .D (
        nx4581), .CLK (CLK)) ;
    oai21 ix4592 (.Y (nx4591), .A0 (nx7471), .A1 (nx8024), .B0 (nx7473)) ;
    dff L0_1_L1_4_Fij_reg_Dout_2 (.Q (FilterDout_1__4__2), .QB (nx7471), .D (
        nx4591), .CLK (CLK)) ;
    oai21 ix4602 (.Y (nx4601), .A0 (nx7477), .A1 (nx8026), .B0 (nx7479)) ;
    dff L0_1_L1_4_Fij_reg_Dout_3 (.Q (FilterDout_1__4__3), .QB (nx7477), .D (
        nx4601), .CLK (CLK)) ;
    oai21 ix4612 (.Y (nx4611), .A0 (nx7483), .A1 (nx8026), .B0 (nx7485)) ;
    dff L0_1_L1_4_Fij_reg_Dout_4 (.Q (FilterDout_1__4__4), .QB (nx7483), .D (
        nx4611), .CLK (CLK)) ;
    oai21 ix4622 (.Y (nx4621), .A0 (nx7489), .A1 (nx8026), .B0 (nx7491)) ;
    dff L0_1_L1_4_Fij_reg_Dout_5 (.Q (FilterDout_1__4__5), .QB (nx7489), .D (
        nx4621), .CLK (CLK)) ;
    oai21 ix4632 (.Y (nx4631), .A0 (nx7495), .A1 (nx8026), .B0 (nx7497)) ;
    dff L0_1_L1_4_Fij_reg_Dout_6 (.Q (FilterDout_1__4__6), .QB (nx7495), .D (
        nx4631), .CLK (CLK)) ;
    oai21 ix4642 (.Y (nx4641), .A0 (nx7501), .A1 (nx8028), .B0 (nx7503)) ;
    dff L0_1_L1_4_Fij_reg_Dout_7 (.Q (FilterDout_1__4__7), .QB (nx7501), .D (
        nx4641), .CLK (CLK)) ;
    oai21 ix4892 (.Y (nx4891), .A0 (nx7507), .A1 (nx8028), .B0 (nx7509)) ;
    dff L0_1_L1_3_Fij_reg_Dout_0 (.Q (FilterDout_1__3__0), .QB (nx7507), .D (
        nx4891), .CLK (CLK)) ;
    oai21 ix4902 (.Y (nx4901), .A0 (nx7513), .A1 (nx8028), .B0 (nx7515)) ;
    dff L0_1_L1_3_Fij_reg_Dout_1 (.Q (FilterDout_1__3__1), .QB (nx7513), .D (
        nx4901), .CLK (CLK)) ;
    oai21 ix4912 (.Y (nx4911), .A0 (nx7519), .A1 (nx8030), .B0 (nx7521)) ;
    dff L0_1_L1_3_Fij_reg_Dout_2 (.Q (FilterDout_1__3__2), .QB (nx7519), .D (
        nx4911), .CLK (CLK)) ;
    oai21 ix4922 (.Y (nx4921), .A0 (nx7525), .A1 (nx8030), .B0 (nx7527)) ;
    dff L0_1_L1_3_Fij_reg_Dout_3 (.Q (FilterDout_1__3__3), .QB (nx7525), .D (
        nx4921), .CLK (CLK)) ;
    oai21 ix4932 (.Y (nx4931), .A0 (nx7531), .A1 (nx8030), .B0 (nx7533)) ;
    dff L0_1_L1_3_Fij_reg_Dout_4 (.Q (FilterDout_1__3__4), .QB (nx7531), .D (
        nx4931), .CLK (CLK)) ;
    oai21 ix4942 (.Y (nx4941), .A0 (nx7537), .A1 (nx8030), .B0 (nx7539)) ;
    dff L0_1_L1_3_Fij_reg_Dout_5 (.Q (FilterDout_1__3__5), .QB (nx7537), .D (
        nx4941), .CLK (CLK)) ;
    oai21 ix4952 (.Y (nx4951), .A0 (nx7543), .A1 (nx8032), .B0 (nx7545)) ;
    dff L0_1_L1_3_Fij_reg_Dout_6 (.Q (FilterDout_1__3__6), .QB (nx7543), .D (
        nx4951), .CLK (CLK)) ;
    oai21 ix4962 (.Y (nx4961), .A0 (nx7549), .A1 (nx8032), .B0 (nx7551)) ;
    dff L0_1_L1_3_Fij_reg_Dout_7 (.Q (FilterDout_1__3__7), .QB (nx7549), .D (
        nx4961), .CLK (CLK)) ;
    oai21 ix5212 (.Y (nx5211), .A0 (nx7555), .A1 (nx8032), .B0 (nx7557)) ;
    dff L0_1_L1_2_Fij_reg_Dout_0 (.Q (FilterDout_1__2__0), .QB (nx7555), .D (
        nx5211), .CLK (CLK)) ;
    nand03 ix7558 (.Y (nx7557), .A0 (nx8158), .A1 (FilterDout_2__2__0), .A2 (
           nx8032)) ;
    oai21 ix5222 (.Y (nx5221), .A0 (nx7561), .A1 (nx8034), .B0 (nx7563)) ;
    dff L0_1_L1_2_Fij_reg_Dout_1 (.Q (FilterDout_1__2__1), .QB (nx7561), .D (
        nx5221), .CLK (CLK)) ;
    nand03 ix7564 (.Y (nx7563), .A0 (nx8158), .A1 (FilterDout_2__2__1), .A2 (
           nx8034)) ;
    oai21 ix5232 (.Y (nx5231), .A0 (nx7567), .A1 (nx8034), .B0 (nx7569)) ;
    dff L0_1_L1_2_Fij_reg_Dout_2 (.Q (FilterDout_1__2__2), .QB (nx7567), .D (
        nx5231), .CLK (CLK)) ;
    nand03 ix7570 (.Y (nx7569), .A0 (nx8158), .A1 (FilterDout_2__2__2), .A2 (
           nx8034)) ;
    oai21 ix5242 (.Y (nx5241), .A0 (nx7573), .A1 (nx8034), .B0 (nx7575)) ;
    dff L0_1_L1_2_Fij_reg_Dout_3 (.Q (FilterDout_1__2__3), .QB (nx7573), .D (
        nx5241), .CLK (CLK)) ;
    nand03 ix7576 (.Y (nx7575), .A0 (nx8160), .A1 (FilterDout_2__2__3), .A2 (
           nx8034)) ;
    oai21 ix5252 (.Y (nx5251), .A0 (nx7579), .A1 (nx8034), .B0 (nx7581)) ;
    dff L0_1_L1_2_Fij_reg_Dout_4 (.Q (FilterDout_1__2__4), .QB (nx7579), .D (
        nx5251), .CLK (CLK)) ;
    nand03 ix7582 (.Y (nx7581), .A0 (nx8160), .A1 (FilterDout_2__2__4), .A2 (
           nx8036)) ;
    oai21 ix5262 (.Y (nx5261), .A0 (nx7585), .A1 (nx8036), .B0 (nx7587)) ;
    dff L0_1_L1_2_Fij_reg_Dout_5 (.Q (FilterDout_1__2__5), .QB (nx7585), .D (
        nx5261), .CLK (CLK)) ;
    nand03 ix7588 (.Y (nx7587), .A0 (nx8160), .A1 (FilterDout_2__2__5), .A2 (
           nx8036)) ;
    oai21 ix5272 (.Y (nx5271), .A0 (nx7591), .A1 (nx8036), .B0 (nx7593)) ;
    dff L0_1_L1_2_Fij_reg_Dout_6 (.Q (FilterDout_1__2__6), .QB (nx7591), .D (
        nx5271), .CLK (CLK)) ;
    nand03 ix7594 (.Y (nx7593), .A0 (nx8160), .A1 (FilterDout_2__2__6), .A2 (
           nx8036)) ;
    oai21 ix5282 (.Y (nx5281), .A0 (nx7597), .A1 (nx8036), .B0 (nx7599)) ;
    dff L0_1_L1_2_Fij_reg_Dout_7 (.Q (FilterDout_1__2__7), .QB (nx7597), .D (
        nx5281), .CLK (CLK)) ;
    nand03 ix7600 (.Y (nx7599), .A0 (nx8160), .A1 (FilterDout_2__2__7), .A2 (
           nx8036)) ;
    oai21 ix5532 (.Y (nx5531), .A0 (nx7603), .A1 (nx8038), .B0 (nx7605)) ;
    dff L0_1_L1_1_Fij_reg_Dout_0 (.Q (FilterDout_1__1__0), .QB (nx7603), .D (
        nx5531), .CLK (CLK)) ;
    nand03 ix7606 (.Y (nx7605), .A0 (nx8160), .A1 (FilterDout_2__1__0), .A2 (
           nx8038)) ;
    oai21 ix5542 (.Y (nx5541), .A0 (nx7609), .A1 (nx8038), .B0 (nx7611)) ;
    dff L0_1_L1_1_Fij_reg_Dout_1 (.Q (FilterDout_1__1__1), .QB (nx7609), .D (
        nx5541), .CLK (CLK)) ;
    nand03 ix7612 (.Y (nx7611), .A0 (nx8160), .A1 (FilterDout_2__1__1), .A2 (
           nx8038)) ;
    oai21 ix5552 (.Y (nx5551), .A0 (nx7615), .A1 (nx8038), .B0 (nx7617)) ;
    dff L0_1_L1_1_Fij_reg_Dout_2 (.Q (FilterDout_1__1__2), .QB (nx7615), .D (
        nx5551), .CLK (CLK)) ;
    nand03 ix7618 (.Y (nx7617), .A0 (nx8162), .A1 (FilterDout_2__1__2), .A2 (
           nx8038)) ;
    oai21 ix5562 (.Y (nx5561), .A0 (nx7621), .A1 (nx8038), .B0 (nx7623)) ;
    dff L0_1_L1_1_Fij_reg_Dout_3 (.Q (FilterDout_1__1__3), .QB (nx7621), .D (
        nx5561), .CLK (CLK)) ;
    nand03 ix7624 (.Y (nx7623), .A0 (nx8162), .A1 (FilterDout_2__1__3), .A2 (
           nx8040)) ;
    oai21 ix5572 (.Y (nx5571), .A0 (nx7627), .A1 (nx8040), .B0 (nx7629)) ;
    dff L0_1_L1_1_Fij_reg_Dout_4 (.Q (FilterDout_1__1__4), .QB (nx7627), .D (
        nx5571), .CLK (CLK)) ;
    nand03 ix7630 (.Y (nx7629), .A0 (nx8162), .A1 (FilterDout_2__1__4), .A2 (
           nx8040)) ;
    oai21 ix5582 (.Y (nx5581), .A0 (nx7633), .A1 (nx8040), .B0 (nx7635)) ;
    dff L0_1_L1_1_Fij_reg_Dout_5 (.Q (FilterDout_1__1__5), .QB (nx7633), .D (
        nx5581), .CLK (CLK)) ;
    nand03 ix7636 (.Y (nx7635), .A0 (nx8162), .A1 (FilterDout_2__1__5), .A2 (
           nx8040)) ;
    oai21 ix5592 (.Y (nx5591), .A0 (nx7639), .A1 (nx8040), .B0 (nx7641)) ;
    dff L0_1_L1_1_Fij_reg_Dout_6 (.Q (FilterDout_1__1__6), .QB (nx7639), .D (
        nx5591), .CLK (CLK)) ;
    nand03 ix7642 (.Y (nx7641), .A0 (nx8162), .A1 (FilterDout_2__1__6), .A2 (
           nx8040)) ;
    oai21 ix5602 (.Y (nx5601), .A0 (nx7645), .A1 (nx8042), .B0 (nx7647)) ;
    dff L0_1_L1_1_Fij_reg_Dout_7 (.Q (FilterDout_1__1__7), .QB (nx7645), .D (
        nx5601), .CLK (CLK)) ;
    nand03 ix7648 (.Y (nx7647), .A0 (nx8162), .A1 (FilterDout_2__1__7), .A2 (
           nx8042)) ;
    oai21 ix5852 (.Y (nx5851), .A0 (nx7651), .A1 (nx8042), .B0 (nx7653)) ;
    dff L0_1_L1_0_Fij_reg_Dout_0 (.Q (FilterDout_1__0__0), .QB (nx7651), .D (
        nx5851), .CLK (CLK)) ;
    nand03 ix7654 (.Y (nx7653), .A0 (nx8162), .A1 (FilterDout_2__0__0), .A2 (
           nx8042)) ;
    oai21 ix5862 (.Y (nx5861), .A0 (nx7657), .A1 (nx8042), .B0 (nx7659)) ;
    dff L0_1_L1_0_Fij_reg_Dout_1 (.Q (FilterDout_1__0__1), .QB (nx7657), .D (
        nx5861), .CLK (CLK)) ;
    nand03 ix7660 (.Y (nx7659), .A0 (nx8164), .A1 (FilterDout_2__0__1), .A2 (
           nx8042)) ;
    oai21 ix5872 (.Y (nx5871), .A0 (nx7663), .A1 (nx8042), .B0 (nx7665)) ;
    dff L0_1_L1_0_Fij_reg_Dout_2 (.Q (FilterDout_1__0__2), .QB (nx7663), .D (
        nx5871), .CLK (CLK)) ;
    nand03 ix7666 (.Y (nx7665), .A0 (nx8164), .A1 (FilterDout_2__0__2), .A2 (
           nx8044)) ;
    oai21 ix5882 (.Y (nx5881), .A0 (nx7669), .A1 (nx8044), .B0 (nx7671)) ;
    dff L0_1_L1_0_Fij_reg_Dout_3 (.Q (FilterDout_1__0__3), .QB (nx7669), .D (
        nx5881), .CLK (CLK)) ;
    nand03 ix7672 (.Y (nx7671), .A0 (nx8164), .A1 (FilterDout_2__0__3), .A2 (
           nx8044)) ;
    oai21 ix5892 (.Y (nx5891), .A0 (nx7675), .A1 (nx8044), .B0 (nx7677)) ;
    dff L0_1_L1_0_Fij_reg_Dout_4 (.Q (FilterDout_1__0__4), .QB (nx7675), .D (
        nx5891), .CLK (CLK)) ;
    nand03 ix7678 (.Y (nx7677), .A0 (nx8164), .A1 (FilterDout_2__0__4), .A2 (
           nx8044)) ;
    oai21 ix5902 (.Y (nx5901), .A0 (nx7681), .A1 (nx8044), .B0 (nx7683)) ;
    dff L0_1_L1_0_Fij_reg_Dout_5 (.Q (FilterDout_1__0__5), .QB (nx7681), .D (
        nx5901), .CLK (CLK)) ;
    nand03 ix7684 (.Y (nx7683), .A0 (nx8164), .A1 (FilterDout_2__0__5), .A2 (
           nx8044)) ;
    oai21 ix5912 (.Y (nx5911), .A0 (nx7687), .A1 (nx8046), .B0 (nx7689)) ;
    dff L0_1_L1_0_Fij_reg_Dout_6 (.Q (FilterDout_1__0__6), .QB (nx7687), .D (
        nx5911), .CLK (CLK)) ;
    nand03 ix7690 (.Y (nx7689), .A0 (nx8164), .A1 (FilterDout_2__0__6), .A2 (
           nx8046)) ;
    oai21 ix5922 (.Y (nx5921), .A0 (nx7693), .A1 (nx8046), .B0 (nx7695)) ;
    dff L0_1_L1_0_Fij_reg_Dout_7 (.Q (FilterDout_1__0__7), .QB (nx7693), .D (
        nx5921), .CLK (CLK)) ;
    nand03 ix7696 (.Y (nx7695), .A0 (nx8164), .A1 (FilterDout_2__0__7), .A2 (
           nx8046)) ;
    oai21 ix4652 (.Y (nx4651), .A0 (nx7699), .A1 (nx8046), .B0 (nx7701)) ;
    dff L0_0_L1_4_Fij_reg_Dout_0 (.Q (FilterDout_0__4__0), .QB (nx7699), .D (
        nx4651), .CLK (CLK)) ;
    oai21 ix4662 (.Y (nx4661), .A0 (nx7705), .A1 (nx8046), .B0 (nx7707)) ;
    dff L0_0_L1_4_Fij_reg_Dout_1 (.Q (FilterDout_0__4__1), .QB (nx7705), .D (
        nx4661), .CLK (CLK)) ;
    oai21 ix4672 (.Y (nx4671), .A0 (nx7711), .A1 (nx8048), .B0 (nx7713)) ;
    dff L0_0_L1_4_Fij_reg_Dout_2 (.Q (FilterDout_0__4__2), .QB (nx7711), .D (
        nx4671), .CLK (CLK)) ;
    oai21 ix4682 (.Y (nx4681), .A0 (nx7717), .A1 (nx8048), .B0 (nx7719)) ;
    dff L0_0_L1_4_Fij_reg_Dout_3 (.Q (FilterDout_0__4__3), .QB (nx7717), .D (
        nx4681), .CLK (CLK)) ;
    oai21 ix4692 (.Y (nx4691), .A0 (nx7723), .A1 (nx8048), .B0 (nx7725)) ;
    dff L0_0_L1_4_Fij_reg_Dout_4 (.Q (FilterDout_0__4__4), .QB (nx7723), .D (
        nx4691), .CLK (CLK)) ;
    oai21 ix4702 (.Y (nx4701), .A0 (nx7729), .A1 (nx8050), .B0 (nx7731)) ;
    dff L0_0_L1_4_Fij_reg_Dout_5 (.Q (FilterDout_0__4__5), .QB (nx7729), .D (
        nx4701), .CLK (CLK)) ;
    oai21 ix4712 (.Y (nx4711), .A0 (nx7735), .A1 (nx8050), .B0 (nx7737)) ;
    dff L0_0_L1_4_Fij_reg_Dout_6 (.Q (FilterDout_0__4__6), .QB (nx7735), .D (
        nx4711), .CLK (CLK)) ;
    oai21 ix4722 (.Y (nx4721), .A0 (nx7741), .A1 (nx8050), .B0 (nx7743)) ;
    dff L0_0_L1_4_Fij_reg_Dout_7 (.Q (FilterDout_0__4__7), .QB (nx7741), .D (
        nx4721), .CLK (CLK)) ;
    oai21 ix4972 (.Y (nx4971), .A0 (nx7747), .A1 (nx8050), .B0 (nx7749)) ;
    dff L0_0_L1_3_Fij_reg_Dout_0 (.Q (FilterDout_0__3__0), .QB (nx7747), .D (
        nx4971), .CLK (CLK)) ;
    oai21 ix4982 (.Y (nx4981), .A0 (nx7753), .A1 (nx8052), .B0 (nx7755)) ;
    dff L0_0_L1_3_Fij_reg_Dout_1 (.Q (FilterDout_0__3__1), .QB (nx7753), .D (
        nx4981), .CLK (CLK)) ;
    oai21 ix4992 (.Y (nx4991), .A0 (nx7759), .A1 (nx8052), .B0 (nx7761)) ;
    dff L0_0_L1_3_Fij_reg_Dout_2 (.Q (FilterDout_0__3__2), .QB (nx7759), .D (
        nx4991), .CLK (CLK)) ;
    oai21 ix5002 (.Y (nx5001), .A0 (nx7765), .A1 (nx8052), .B0 (nx7767)) ;
    dff L0_0_L1_3_Fij_reg_Dout_3 (.Q (FilterDout_0__3__3), .QB (nx7765), .D (
        nx5001), .CLK (CLK)) ;
    oai21 ix5012 (.Y (nx5011), .A0 (nx7771), .A1 (nx8054), .B0 (nx7773)) ;
    dff L0_0_L1_3_Fij_reg_Dout_4 (.Q (FilterDout_0__3__4), .QB (nx7771), .D (
        nx5011), .CLK (CLK)) ;
    oai21 ix5022 (.Y (nx5021), .A0 (nx7777), .A1 (nx8054), .B0 (nx7779)) ;
    dff L0_0_L1_3_Fij_reg_Dout_5 (.Q (FilterDout_0__3__5), .QB (nx7777), .D (
        nx5021), .CLK (CLK)) ;
    oai21 ix5032 (.Y (nx5031), .A0 (nx7783), .A1 (nx8054), .B0 (nx7785)) ;
    dff L0_0_L1_3_Fij_reg_Dout_6 (.Q (FilterDout_0__3__6), .QB (nx7783), .D (
        nx5031), .CLK (CLK)) ;
    oai21 ix5042 (.Y (nx5041), .A0 (nx7789), .A1 (nx8054), .B0 (nx7791)) ;
    dff L0_0_L1_3_Fij_reg_Dout_7 (.Q (FilterDout_0__3__7), .QB (nx7789), .D (
        nx5041), .CLK (CLK)) ;
    oai21 ix5292 (.Y (nx5291), .A0 (nx7795), .A1 (nx8056), .B0 (nx7797)) ;
    dff L0_0_L1_2_Fij_reg_Dout_0 (.Q (FilterDout_0__2__0), .QB (nx7795), .D (
        nx5291), .CLK (CLK)) ;
    oai21 ix5302 (.Y (nx5301), .A0 (nx7801), .A1 (nx8056), .B0 (nx7803)) ;
    dff L0_0_L1_2_Fij_reg_Dout_1 (.Q (FilterDout_0__2__1), .QB (nx7801), .D (
        nx5301), .CLK (CLK)) ;
    oai21 ix5312 (.Y (nx5311), .A0 (nx7807), .A1 (nx8056), .B0 (nx7809)) ;
    dff L0_0_L1_2_Fij_reg_Dout_2 (.Q (FilterDout_0__2__2), .QB (nx7807), .D (
        nx5311), .CLK (CLK)) ;
    oai21 ix5322 (.Y (nx5321), .A0 (nx7813), .A1 (nx8058), .B0 (nx7815)) ;
    dff L0_0_L1_2_Fij_reg_Dout_3 (.Q (FilterDout_0__2__3), .QB (nx7813), .D (
        nx5321), .CLK (CLK)) ;
    oai21 ix5332 (.Y (nx5331), .A0 (nx7819), .A1 (nx8058), .B0 (nx7821)) ;
    dff L0_0_L1_2_Fij_reg_Dout_4 (.Q (FilterDout_0__2__4), .QB (nx7819), .D (
        nx5331), .CLK (CLK)) ;
    oai21 ix5342 (.Y (nx5341), .A0 (nx7825), .A1 (nx8058), .B0 (nx7827)) ;
    dff L0_0_L1_2_Fij_reg_Dout_5 (.Q (FilterDout_0__2__5), .QB (nx7825), .D (
        nx5341), .CLK (CLK)) ;
    oai21 ix5352 (.Y (nx5351), .A0 (nx7831), .A1 (nx8058), .B0 (nx7833)) ;
    dff L0_0_L1_2_Fij_reg_Dout_6 (.Q (FilterDout_0__2__6), .QB (nx7831), .D (
        nx5351), .CLK (CLK)) ;
    oai21 ix5362 (.Y (nx5361), .A0 (nx7837), .A1 (nx8060), .B0 (nx7839)) ;
    dff L0_0_L1_2_Fij_reg_Dout_7 (.Q (FilterDout_0__2__7), .QB (nx7837), .D (
        nx5361), .CLK (CLK)) ;
    oai21 ix5612 (.Y (nx5611), .A0 (nx7843), .A1 (nx8060), .B0 (nx7845)) ;
    dff L0_0_L1_1_Fij_reg_Dout_0 (.Q (FilterDout_0__1__0), .QB (nx7843), .D (
        nx5611), .CLK (CLK)) ;
    oai21 ix5622 (.Y (nx5621), .A0 (nx7849), .A1 (nx8060), .B0 (nx7851)) ;
    dff L0_0_L1_1_Fij_reg_Dout_1 (.Q (FilterDout_0__1__1), .QB (nx7849), .D (
        nx5621), .CLK (CLK)) ;
    oai21 ix5632 (.Y (nx5631), .A0 (nx7855), .A1 (nx8062), .B0 (nx7857)) ;
    dff L0_0_L1_1_Fij_reg_Dout_2 (.Q (FilterDout_0__1__2), .QB (nx7855), .D (
        nx5631), .CLK (CLK)) ;
    oai21 ix5642 (.Y (nx5641), .A0 (nx7861), .A1 (nx8062), .B0 (nx7863)) ;
    dff L0_0_L1_1_Fij_reg_Dout_3 (.Q (FilterDout_0__1__3), .QB (nx7861), .D (
        nx5641), .CLK (CLK)) ;
    oai21 ix5652 (.Y (nx5651), .A0 (nx7867), .A1 (nx8062), .B0 (nx7869)) ;
    dff L0_0_L1_1_Fij_reg_Dout_4 (.Q (FilterDout_0__1__4), .QB (nx7867), .D (
        nx5651), .CLK (CLK)) ;
    oai21 ix5662 (.Y (nx5661), .A0 (nx7873), .A1 (nx8062), .B0 (nx7875)) ;
    dff L0_0_L1_1_Fij_reg_Dout_5 (.Q (FilterDout_0__1__5), .QB (nx7873), .D (
        nx5661), .CLK (CLK)) ;
    oai21 ix5672 (.Y (nx5671), .A0 (nx7879), .A1 (nx8064), .B0 (nx7881)) ;
    dff L0_0_L1_1_Fij_reg_Dout_6 (.Q (FilterDout_0__1__6), .QB (nx7879), .D (
        nx5671), .CLK (CLK)) ;
    oai21 ix5682 (.Y (nx5681), .A0 (nx7885), .A1 (nx8064), .B0 (nx7887)) ;
    dff L0_0_L1_1_Fij_reg_Dout_7 (.Q (FilterDout_0__1__7), .QB (nx7885), .D (
        nx5681), .CLK (CLK)) ;
    oai21 ix5932 (.Y (nx5931), .A0 (nx7891), .A1 (nx8064), .B0 (nx7893)) ;
    dff L0_0_L1_0_Fij_reg_Dout_0 (.Q (FilterDout_0__0__0), .QB (nx7891), .D (
        nx5931), .CLK (CLK)) ;
    oai21 ix5942 (.Y (nx5941), .A0 (nx7897), .A1 (nx8066), .B0 (nx7899)) ;
    dff L0_0_L1_0_Fij_reg_Dout_1 (.Q (FilterDout_0__0__1), .QB (nx7897), .D (
        nx5941), .CLK (CLK)) ;
    oai21 ix5952 (.Y (nx5951), .A0 (nx7903), .A1 (nx8066), .B0 (nx7905)) ;
    dff L0_0_L1_0_Fij_reg_Dout_2 (.Q (FilterDout_0__0__2), .QB (nx7903), .D (
        nx5951), .CLK (CLK)) ;
    oai21 ix5962 (.Y (nx5961), .A0 (nx7909), .A1 (nx8066), .B0 (nx7911)) ;
    dff L0_0_L1_0_Fij_reg_Dout_3 (.Q (FilterDout_0__0__3), .QB (nx7909), .D (
        nx5961), .CLK (CLK)) ;
    oai21 ix5972 (.Y (nx5971), .A0 (nx7915), .A1 (nx8066), .B0 (nx7917)) ;
    dff L0_0_L1_0_Fij_reg_Dout_4 (.Q (FilterDout_0__0__4), .QB (nx7915), .D (
        nx5971), .CLK (CLK)) ;
    oai21 ix5982 (.Y (nx5981), .A0 (nx7921), .A1 (nx8068), .B0 (nx7923)) ;
    dff L0_0_L1_0_Fij_reg_Dout_5 (.Q (FilterDout_0__0__5), .QB (nx7921), .D (
        nx5981), .CLK (CLK)) ;
    oai21 ix5992 (.Y (nx5991), .A0 (nx7927), .A1 (nx8068), .B0 (nx7929)) ;
    dff L0_0_L1_0_Fij_reg_Dout_6 (.Q (FilterDout_0__0__6), .QB (nx7927), .D (
        nx5991), .CLK (CLK)) ;
    oai21 ix6002 (.Y (nx6001), .A0 (nx7933), .A1 (nx8068), .B0 (nx7935)) ;
    dff L0_0_L1_0_Fij_reg_Dout_7 (.Q (FilterDout_0__0__7), .QB (nx7933), .D (
        nx6001), .CLK (CLK)) ;
    inv02 ix169 (.Y (nx168), .A (nx6998)) ;
    inv02 ix85 (.Y (nx84), .A (nx6042)) ;
    inv02 ix7941 (.Y (nx7942), .A (nx8182)) ;
    inv02 ix7943 (.Y (nx7944), .A (nx8182)) ;
    inv02 ix7945 (.Y (nx7946), .A (nx8182)) ;
    inv02 ix7947 (.Y (nx7948), .A (nx8182)) ;
    inv02 ix7949 (.Y (nx7950), .A (nx8182)) ;
    inv02 ix7951 (.Y (nx7952), .A (nx8278)) ;
    inv02 ix7953 (.Y (nx7954), .A (nx8278)) ;
    inv02 ix7955 (.Y (nx7956), .A (nx8278)) ;
    inv02 ix7957 (.Y (nx7958), .A (nx8278)) ;
    inv02 ix7959 (.Y (nx7960), .A (nx8278)) ;
    inv02 ix7961 (.Y (nx7962), .A (nx8278)) ;
    inv02 ix7963 (.Y (nx7964), .A (nx8278)) ;
    inv02 ix7965 (.Y (nx7966), .A (nx8286)) ;
    inv02 ix7967 (.Y (nx7968), .A (nx8286)) ;
    inv02 ix7969 (.Y (nx7970), .A (nx8286)) ;
    inv02 ix7971 (.Y (nx7972), .A (nx8286)) ;
    inv02 ix7973 (.Y (nx7974), .A (nx8286)) ;
    inv02 ix7975 (.Y (nx7976), .A (nx8286)) ;
    inv02 ix7977 (.Y (nx7978), .A (nx8286)) ;
    inv02 ix7979 (.Y (nx7980), .A (nx8288)) ;
    inv02 ix7981 (.Y (nx7982), .A (nx8288)) ;
    inv02 ix7983 (.Y (nx7984), .A (nx8288)) ;
    inv02 ix7985 (.Y (nx7986), .A (nx8288)) ;
    inv02 ix7987 (.Y (nx7988), .A (nx8288)) ;
    inv02 ix7989 (.Y (nx7990), .A (nx8288)) ;
    inv02 ix7991 (.Y (nx7992), .A (nx8288)) ;
    inv02 ix7993 (.Y (nx7994), .A (nx8294)) ;
    inv02 ix7995 (.Y (nx7996), .A (nx8294)) ;
    inv02 ix7997 (.Y (nx7998), .A (nx8294)) ;
    inv02 ix7999 (.Y (nx8000), .A (nx8294)) ;
    inv02 ix8001 (.Y (nx8002), .A (nx8294)) ;
    inv02 ix8003 (.Y (nx8004), .A (nx8294)) ;
    inv02 ix8005 (.Y (nx8006), .A (nx8220)) ;
    inv02 ix8007 (.Y (nx8008), .A (nx8220)) ;
    inv02 ix8009 (.Y (nx8010), .A (nx8220)) ;
    inv02 ix8011 (.Y (nx8012), .A (nx8220)) ;
    inv02 ix8013 (.Y (nx8014), .A (nx8220)) ;
    inv02 ix8015 (.Y (nx8016), .A (nx8300)) ;
    inv02 ix8017 (.Y (nx8018), .A (nx8300)) ;
    inv02 ix8019 (.Y (nx8020), .A (nx8300)) ;
    inv02 ix8021 (.Y (nx8022), .A (nx8300)) ;
    inv02 ix8023 (.Y (nx8024), .A (nx8300)) ;
    inv02 ix8025 (.Y (nx8026), .A (nx8300)) ;
    inv02 ix8027 (.Y (nx8028), .A (nx8300)) ;
    inv02 ix8029 (.Y (nx8030), .A (nx8308)) ;
    inv02 ix8031 (.Y (nx8032), .A (nx8308)) ;
    inv02 ix8033 (.Y (nx8034), .A (nx8308)) ;
    inv02 ix8035 (.Y (nx8036), .A (nx8308)) ;
    inv02 ix8037 (.Y (nx8038), .A (nx8308)) ;
    inv02 ix8039 (.Y (nx8040), .A (nx8308)) ;
    inv02 ix8041 (.Y (nx8042), .A (nx8308)) ;
    inv02 ix8043 (.Y (nx8044), .A (nx8310)) ;
    inv02 ix8045 (.Y (nx8046), .A (nx8310)) ;
    inv02 ix8047 (.Y (nx8048), .A (nx8310)) ;
    inv02 ix8049 (.Y (nx8050), .A (nx8310)) ;
    inv02 ix8051 (.Y (nx8052), .A (nx8310)) ;
    inv02 ix8053 (.Y (nx8054), .A (nx8310)) ;
    inv02 ix8055 (.Y (nx8056), .A (nx8310)) ;
    inv02 ix8057 (.Y (nx8058), .A (nx8316)) ;
    inv02 ix8059 (.Y (nx8060), .A (nx8316)) ;
    inv02 ix8061 (.Y (nx8062), .A (nx8316)) ;
    inv02 ix8063 (.Y (nx8064), .A (nx8316)) ;
    inv02 ix8065 (.Y (nx8066), .A (nx8316)) ;
    inv02 ix8067 (.Y (nx8068), .A (nx8316)) ;
    inv02 ix8069 (.Y (nx8070), .A (RST)) ;
    inv02 ix8071 (.Y (nx8072), .A (RST)) ;
    inv02 ix8073 (.Y (nx8074), .A (RST)) ;
    inv02 ix8075 (.Y (nx8076), .A (RST)) ;
    inv02 ix8077 (.Y (nx8078), .A (RST)) ;
    inv02 ix8079 (.Y (nx8080), .A (RST)) ;
    inv02 ix8081 (.Y (nx8082), .A (RST)) ;
    inv02 ix8083 (.Y (nx8084), .A (RST)) ;
    inv02 ix8085 (.Y (nx8086), .A (RST)) ;
    inv02 ix8087 (.Y (nx8088), .A (RST)) ;
    inv02 ix8089 (.Y (nx8090), .A (RST)) ;
    inv02 ix8093 (.Y (nx8094), .A (RST)) ;
    inv02 ix8095 (.Y (nx8096), .A (RST)) ;
    inv02 ix8097 (.Y (nx8098), .A (RST)) ;
    inv02 ix8099 (.Y (nx8100), .A (RST)) ;
    inv02 ix8105 (.Y (nx8106), .A (RST)) ;
    inv02 ix8107 (.Y (nx8108), .A (RST)) ;
    inv02 ix8109 (.Y (nx8110), .A (RST)) ;
    inv02 ix8111 (.Y (nx8112), .A (RST)) ;
    inv02 ix8123 (.Y (nx8124), .A (RST)) ;
    inv02 ix8125 (.Y (nx8126), .A (RST)) ;
    inv02 ix8127 (.Y (nx8128), .A (RST)) ;
    inv02 ix8129 (.Y (nx8130), .A (RST)) ;
    inv02 ix8131 (.Y (nx8132), .A (RST)) ;
    inv02 ix8133 (.Y (nx8134), .A (RST)) ;
    inv02 ix8135 (.Y (nx8136), .A (RST)) ;
    inv02 ix8137 (.Y (nx8138), .A (RST)) ;
    inv02 ix8139 (.Y (nx8140), .A (RST)) ;
    inv02 ix8141 (.Y (nx8142), .A (RST)) ;
    inv02 ix8145 (.Y (nx8146), .A (RST)) ;
    inv02 ix8147 (.Y (nx8148), .A (RST)) ;
    inv02 ix8149 (.Y (nx8150), .A (RST)) ;
    inv02 ix8151 (.Y (nx8152), .A (RST)) ;
    inv02 ix8153 (.Y (nx8154), .A (RST)) ;
    inv02 ix8157 (.Y (nx8158), .A (RST)) ;
    inv02 ix8159 (.Y (nx8160), .A (RST)) ;
    inv02 ix8161 (.Y (nx8162), .A (RST)) ;
    inv02 ix8163 (.Y (nx8164), .A (RST)) ;
    inv02 ix8181 (.Y (nx8182), .A (nx8322)) ;
    inv02 ix8183 (.Y (nx8184), .A (nx8322)) ;
    inv02 ix8185 (.Y (nx8186), .A (nx8322)) ;
    inv02 ix8187 (.Y (nx8188), .A (nx8322)) ;
    inv02 ix8189 (.Y (nx8190), .A (nx8322)) ;
    inv02 ix8193 (.Y (nx8194), .A (nx8254)) ;
    inv02 ix8195 (.Y (nx8196), .A (nx8254)) ;
    inv02 ix8197 (.Y (nx8198), .A (nx8254)) ;
    inv02 ix8199 (.Y (nx8200), .A (nx8254)) ;
    inv02 ix8201 (.Y (nx8202), .A (nx8254)) ;
    inv02 ix8203 (.Y (nx8204), .A (nx8254)) ;
    inv02 ix8205 (.Y (nx8206), .A (nx8254)) ;
    inv02 ix8207 (.Y (nx8208), .A (nx8256)) ;
    inv02 ix8209 (.Y (nx8210), .A (nx8256)) ;
    inv02 ix8211 (.Y (nx8212), .A (nx8256)) ;
    inv02 ix8213 (.Y (nx8214), .A (nx8256)) ;
    inv02 ix8219 (.Y (nx8220), .A (nx8326)) ;
    inv02 ix8221 (.Y (nx8222), .A (nx8326)) ;
    inv02 ix8223 (.Y (nx8224), .A (nx8326)) ;
    inv02 ix8225 (.Y (nx8226), .A (nx8326)) ;
    inv02 ix8227 (.Y (nx8228), .A (nx8326)) ;
    inv02 ix8231 (.Y (nx8232), .A (nx8258)) ;
    inv02 ix8233 (.Y (nx8234), .A (nx8258)) ;
    inv02 ix8235 (.Y (nx8236), .A (nx8258)) ;
    inv02 ix8237 (.Y (nx8238), .A (nx8258)) ;
    inv02 ix8239 (.Y (nx8240), .A (nx8258)) ;
    inv02 ix8241 (.Y (nx8242), .A (nx8258)) ;
    inv02 ix8243 (.Y (nx8244), .A (nx8258)) ;
    inv02 ix8245 (.Y (nx8246), .A (nx8260)) ;
    inv02 ix8247 (.Y (nx8248), .A (nx8260)) ;
    inv02 ix8249 (.Y (nx8250), .A (nx8260)) ;
    inv02 ix8251 (.Y (nx8252), .A (nx8260)) ;
    inv02 ix8253 (.Y (nx8254), .A (nx6107)) ;
    inv02 ix8255 (.Y (nx8256), .A (nx6107)) ;
    inv02 ix8257 (.Y (nx8258), .A (nx7048)) ;
    inv02 ix8259 (.Y (nx8260), .A (nx7048)) ;
    mux21_ni ix2012 (.Y (nx2011), .A0 (WindowDout_4__4__0), .A1 (nx88), .S0 (
             nx8322)) ;
    mux21_ni ix2022 (.Y (nx2021), .A0 (WindowDout_4__4__1), .A1 (nx98), .S0 (
             nx8322)) ;
    mux21_ni ix2032 (.Y (nx2031), .A0 (WindowDout_4__4__2), .A1 (nx108), .S0 (
             nx8272)) ;
    mux21_ni ix2042 (.Y (nx2041), .A0 (WindowDout_4__4__3), .A1 (nx118), .S0 (
             nx8272)) ;
    mux21_ni ix2052 (.Y (nx2051), .A0 (WindowDout_4__4__4), .A1 (nx128), .S0 (
             nx8272)) ;
    mux21_ni ix2062 (.Y (nx2061), .A0 (WindowDout_4__4__5), .A1 (nx138), .S0 (
             nx8272)) ;
    mux21_ni ix2072 (.Y (nx2071), .A0 (WindowDout_4__4__6), .A1 (nx148), .S0 (
             nx8272)) ;
    mux21_ni ix2082 (.Y (nx2081), .A0 (WindowDout_4__4__7), .A1 (nx158), .S0 (
             nx8272)) ;
    mux21_ni ix2172 (.Y (nx2171), .A0 (WindowDout_4__3__0), .A1 (nx220), .S0 (
             nx8272)) ;
    mux21_ni ix2182 (.Y (nx2181), .A0 (WindowDout_4__3__1), .A1 (nx230), .S0 (
             nx84)) ;
    mux21_ni ix2192 (.Y (nx2191), .A0 (WindowDout_4__3__2), .A1 (nx240), .S0 (
             nx84)) ;
    mux21_ni ix2202 (.Y (nx2201), .A0 (WindowDout_4__3__3), .A1 (nx250), .S0 (
             nx84)) ;
    mux21_ni ix2212 (.Y (nx2211), .A0 (WindowDout_4__3__4), .A1 (nx260), .S0 (
             nx84)) ;
    mux21_ni ix2222 (.Y (nx2221), .A0 (WindowDout_4__3__5), .A1 (nx270), .S0 (
             nx84)) ;
    mux21_ni ix2232 (.Y (nx2231), .A0 (WindowDout_4__3__6), .A1 (nx280), .S0 (
             nx84)) ;
    mux21_ni ix2242 (.Y (nx2241), .A0 (WindowDout_4__3__7), .A1 (nx290), .S0 (
             nx84)) ;
    or03 ix6353 (.Y (nx6352), .A0 (RST), .A1 (nx6181), .A2 (nx8182)) ;
    or03 ix6359 (.Y (nx6358), .A0 (RST), .A1 (nx6188), .A2 (nx8280)) ;
    or03 ix6365 (.Y (nx6364), .A0 (RST), .A1 (nx6194), .A2 (nx8280)) ;
    or03 ix6371 (.Y (nx6370), .A0 (RST), .A1 (nx6200), .A2 (nx8280)) ;
    or03 ix6377 (.Y (nx6376), .A0 (RST), .A1 (nx6206), .A2 (nx8280)) ;
    or03 ix6383 (.Y (nx6382), .A0 (RST), .A1 (nx6212), .A2 (nx8280)) ;
    or03 ix6389 (.Y (nx6388), .A0 (RST), .A1 (nx6218), .A2 (nx8280)) ;
    or03 ix6395 (.Y (nx6394), .A0 (RST), .A1 (nx6224), .A2 (nx8280)) ;
    or03 ix6401 (.Y (nx6400), .A0 (RST), .A1 (nx6230), .A2 (nx8282)) ;
    or03 ix6407 (.Y (nx6406), .A0 (RST), .A1 (nx6236), .A2 (nx8282)) ;
    or03 ix6413 (.Y (nx6412), .A0 (RST), .A1 (nx6242), .A2 (nx8282)) ;
    or03 ix6419 (.Y (nx6418), .A0 (RST), .A1 (nx6248), .A2 (nx8282)) ;
    or03 ix6425 (.Y (nx6424), .A0 (RST), .A1 (nx6254), .A2 (nx8282)) ;
    or03 ix6431 (.Y (nx6430), .A0 (RST), .A1 (nx6260), .A2 (nx8282)) ;
    or03 ix6437 (.Y (nx6436), .A0 (RST), .A1 (nx6266), .A2 (nx8282)) ;
    or03 ix6443 (.Y (nx6442), .A0 (RST), .A1 (nx6272), .A2 (nx8284)) ;
    or03 ix6521 (.Y (nx6520), .A0 (RST), .A1 (nx6350), .A2 (nx8284)) ;
    or03 ix6527 (.Y (nx6526), .A0 (RST), .A1 (nx6356), .A2 (nx8284)) ;
    or03 ix6533 (.Y (nx6532), .A0 (RST), .A1 (nx6362), .A2 (nx8284)) ;
    or03 ix6539 (.Y (nx6538), .A0 (RST), .A1 (nx6368), .A2 (nx8284)) ;
    or03 ix6545 (.Y (nx6544), .A0 (RST), .A1 (nx6374), .A2 (nx8284)) ;
    or03 ix6551 (.Y (nx6550), .A0 (RST), .A1 (nx6380), .A2 (nx8284)) ;
    or03 ix6557 (.Y (nx6556), .A0 (RST), .A1 (nx6386), .A2 (nx8184)) ;
    or03 ix6563 (.Y (nx6562), .A0 (RST), .A1 (nx6392), .A2 (nx8184)) ;
    or03 ix6569 (.Y (nx6568), .A0 (RST), .A1 (nx6398), .A2 (nx8184)) ;
    or03 ix6575 (.Y (nx6574), .A0 (RST), .A1 (nx6404), .A2 (nx8184)) ;
    or03 ix6581 (.Y (nx6580), .A0 (RST), .A1 (nx6410), .A2 (nx8186)) ;
    or03 ix6587 (.Y (nx6586), .A0 (RST), .A1 (nx6416), .A2 (nx8186)) ;
    or03 ix6593 (.Y (nx6592), .A0 (RST), .A1 (nx6422), .A2 (nx8186)) ;
    or03 ix6599 (.Y (nx6598), .A0 (RST), .A1 (nx6428), .A2 (nx8186)) ;
    or03 ix6605 (.Y (nx6604), .A0 (RST), .A1 (nx6434), .A2 (nx8186)) ;
    or03 ix6611 (.Y (nx6610), .A0 (RST), .A1 (nx6440), .A2 (nx8186)) ;
    or03 ix6761 (.Y (nx6760), .A0 (RST), .A1 (nx6518), .A2 (nx8290)) ;
    or03 ix6767 (.Y (nx6766), .A0 (RST), .A1 (nx6524), .A2 (nx8290)) ;
    or03 ix6773 (.Y (nx6772), .A0 (RST), .A1 (nx6530), .A2 (nx8290)) ;
    or03 ix6779 (.Y (nx6778), .A0 (RST), .A1 (nx6536), .A2 (nx8290)) ;
    or03 ix6785 (.Y (nx6784), .A0 (RST), .A1 (nx6542), .A2 (nx8290)) ;
    or03 ix6791 (.Y (nx6790), .A0 (RST), .A1 (nx6548), .A2 (nx8290)) ;
    or03 ix6797 (.Y (nx6796), .A0 (RST), .A1 (nx6554), .A2 (nx8290)) ;
    or03 ix6803 (.Y (nx6802), .A0 (RST), .A1 (nx6560), .A2 (nx8292)) ;
    or03 ix6809 (.Y (nx6808), .A0 (RST), .A1 (nx6566), .A2 (nx8292)) ;
    or03 ix6815 (.Y (nx6814), .A0 (RST), .A1 (nx6572), .A2 (nx8292)) ;
    or03 ix6821 (.Y (nx6820), .A0 (RST), .A1 (nx6578), .A2 (nx8292)) ;
    or03 ix6827 (.Y (nx6826), .A0 (RST), .A1 (nx6584), .A2 (nx8292)) ;
    or03 ix6833 (.Y (nx6832), .A0 (RST), .A1 (nx6590), .A2 (nx8292)) ;
    or03 ix6839 (.Y (nx6838), .A0 (RST), .A1 (nx6596), .A2 (nx8292)) ;
    or03 ix6845 (.Y (nx6844), .A0 (RST), .A1 (nx6602), .A2 (nx8188)) ;
    or03 ix6851 (.Y (nx6850), .A0 (RST), .A1 (nx6608), .A2 (nx8188)) ;
    or03 ix6857 (.Y (nx6856), .A0 (RST), .A1 (nx6614), .A2 (nx8188)) ;
    or03 ix6863 (.Y (nx6862), .A0 (RST), .A1 (nx6620), .A2 (nx8188)) ;
    or03 ix6869 (.Y (nx6868), .A0 (RST), .A1 (nx6626), .A2 (nx8188)) ;
    or03 ix6875 (.Y (nx6874), .A0 (RST), .A1 (nx6632), .A2 (nx8294)) ;
    or03 ix6881 (.Y (nx6880), .A0 (RST), .A1 (nx6638), .A2 (nx8296)) ;
    or03 ix6887 (.Y (nx6886), .A0 (RST), .A1 (nx6644), .A2 (nx8296)) ;
    or03 ix6893 (.Y (nx6892), .A0 (RST), .A1 (nx6650), .A2 (nx8296)) ;
    or03 ix6899 (.Y (nx6898), .A0 (RST), .A1 (nx6656), .A2 (nx8296)) ;
    or03 ix6905 (.Y (nx6904), .A0 (RST), .A1 (nx6662), .A2 (nx8296)) ;
    or03 ix6911 (.Y (nx6910), .A0 (RST), .A1 (nx6668), .A2 (nx8296)) ;
    or03 ix6917 (.Y (nx6916), .A0 (RST), .A1 (nx6674), .A2 (nx8296)) ;
    or03 ix6923 (.Y (nx6922), .A0 (RST), .A1 (nx6680), .A2 (nx8298)) ;
    or03 ix6929 (.Y (nx6928), .A0 (RST), .A1 (nx6686), .A2 (nx8298)) ;
    or03 ix6935 (.Y (nx6934), .A0 (RST), .A1 (nx6692), .A2 (nx8298)) ;
    or03 ix6941 (.Y (nx6940), .A0 (RST), .A1 (nx6698), .A2 (nx8298)) ;
    or03 ix6947 (.Y (nx6946), .A0 (RST), .A1 (nx6704), .A2 (nx8298)) ;
    or03 ix6953 (.Y (nx6952), .A0 (RST), .A1 (nx6710), .A2 (nx8298)) ;
    or03 ix6959 (.Y (nx6958), .A0 (RST), .A1 (nx6716), .A2 (nx8298)) ;
    or03 ix6965 (.Y (nx6964), .A0 (RST), .A1 (nx6722), .A2 (nx8190)) ;
    or03 ix6971 (.Y (nx6970), .A0 (RST), .A1 (nx6728), .A2 (nx8190)) ;
    or03 ix6977 (.Y (nx6976), .A0 (RST), .A1 (nx6734), .A2 (nx8190)) ;
    or03 ix6983 (.Y (nx6982), .A0 (RST), .A1 (nx6740), .A2 (nx8190)) ;
    or03 ix6989 (.Y (nx6988), .A0 (RST), .A1 (nx6746), .A2 (nx8190)) ;
    or03 ix6995 (.Y (nx6994), .A0 (RST), .A1 (nx6752), .A2 (nx8190)) ;
    mux21_ni ix2092 (.Y (nx2091), .A0 (FilterDout_4__4__0), .A1 (nx88), .S0 (
             nx8326)) ;
    mux21_ni ix2102 (.Y (nx2101), .A0 (FilterDout_4__4__1), .A1 (nx98), .S0 (
             nx8326)) ;
    mux21_ni ix2112 (.Y (nx2111), .A0 (FilterDout_4__4__2), .A1 (nx108), .S0 (
             nx8276)) ;
    mux21_ni ix2122 (.Y (nx2121), .A0 (FilterDout_4__4__3), .A1 (nx118), .S0 (
             nx8276)) ;
    mux21_ni ix2132 (.Y (nx2131), .A0 (FilterDout_4__4__4), .A1 (nx128), .S0 (
             nx8276)) ;
    mux21_ni ix2142 (.Y (nx2141), .A0 (FilterDout_4__4__5), .A1 (nx138), .S0 (
             nx8276)) ;
    mux21_ni ix2152 (.Y (nx2151), .A0 (FilterDout_4__4__6), .A1 (nx148), .S0 (
             nx8276)) ;
    mux21_ni ix2162 (.Y (nx2161), .A0 (FilterDout_4__4__7), .A1 (nx158), .S0 (
             nx8276)) ;
    mux21_ni ix2252 (.Y (nx2251), .A0 (FilterDout_4__3__0), .A1 (nx220), .S0 (
             nx8276)) ;
    mux21_ni ix2262 (.Y (nx2261), .A0 (FilterDout_4__3__1), .A1 (nx230), .S0 (
             nx168)) ;
    mux21_ni ix2272 (.Y (nx2271), .A0 (FilterDout_4__3__2), .A1 (nx240), .S0 (
             nx168)) ;
    mux21_ni ix2282 (.Y (nx2281), .A0 (FilterDout_4__3__3), .A1 (nx250), .S0 (
             nx168)) ;
    mux21_ni ix2292 (.Y (nx2291), .A0 (FilterDout_4__3__4), .A1 (nx260), .S0 (
             nx168)) ;
    mux21_ni ix2302 (.Y (nx2301), .A0 (FilterDout_4__3__5), .A1 (nx270), .S0 (
             nx168)) ;
    mux21_ni ix2312 (.Y (nx2311), .A0 (FilterDout_4__3__6), .A1 (nx280), .S0 (
             nx168)) ;
    mux21_ni ix2322 (.Y (nx2321), .A0 (FilterDout_4__3__7), .A1 (nx290), .S0 (
             nx168)) ;
    or03 ix7294 (.Y (nx7293), .A0 (RST), .A1 (nx7122), .A2 (nx8220)) ;
    or03 ix7300 (.Y (nx7299), .A0 (RST), .A1 (nx7129), .A2 (nx8302)) ;
    or03 ix7306 (.Y (nx7305), .A0 (RST), .A1 (nx7135), .A2 (nx8302)) ;
    or03 ix7312 (.Y (nx7311), .A0 (RST), .A1 (nx7141), .A2 (nx8302)) ;
    or03 ix7318 (.Y (nx7317), .A0 (RST), .A1 (nx7147), .A2 (nx8302)) ;
    or03 ix7324 (.Y (nx7323), .A0 (RST), .A1 (nx7153), .A2 (nx8302)) ;
    or03 ix7330 (.Y (nx7329), .A0 (RST), .A1 (nx7159), .A2 (nx8302)) ;
    or03 ix7336 (.Y (nx7335), .A0 (RST), .A1 (nx7165), .A2 (nx8302)) ;
    or03 ix7342 (.Y (nx7341), .A0 (RST), .A1 (nx7171), .A2 (nx8304)) ;
    or03 ix7348 (.Y (nx7347), .A0 (RST), .A1 (nx7177), .A2 (nx8304)) ;
    or03 ix7354 (.Y (nx7353), .A0 (RST), .A1 (nx7183), .A2 (nx8304)) ;
    or03 ix7360 (.Y (nx7359), .A0 (RST), .A1 (nx7189), .A2 (nx8304)) ;
    or03 ix7366 (.Y (nx7365), .A0 (RST), .A1 (nx7195), .A2 (nx8304)) ;
    or03 ix7372 (.Y (nx7371), .A0 (RST), .A1 (nx7201), .A2 (nx8304)) ;
    or03 ix7378 (.Y (nx7377), .A0 (RST), .A1 (nx7207), .A2 (nx8304)) ;
    or03 ix7384 (.Y (nx7383), .A0 (RST), .A1 (nx7213), .A2 (nx8306)) ;
    or03 ix7462 (.Y (nx7461), .A0 (RST), .A1 (nx7291), .A2 (nx8306)) ;
    or03 ix7468 (.Y (nx7467), .A0 (RST), .A1 (nx7297), .A2 (nx8306)) ;
    or03 ix7474 (.Y (nx7473), .A0 (RST), .A1 (nx7303), .A2 (nx8306)) ;
    or03 ix7480 (.Y (nx7479), .A0 (RST), .A1 (nx7309), .A2 (nx8306)) ;
    or03 ix7486 (.Y (nx7485), .A0 (RST), .A1 (nx7315), .A2 (nx8306)) ;
    or03 ix7492 (.Y (nx7491), .A0 (RST), .A1 (nx7321), .A2 (nx8306)) ;
    or03 ix7498 (.Y (nx7497), .A0 (RST), .A1 (nx7327), .A2 (nx8222)) ;
    or03 ix7504 (.Y (nx7503), .A0 (RST), .A1 (nx7333), .A2 (nx8222)) ;
    or03 ix7510 (.Y (nx7509), .A0 (RST), .A1 (nx7339), .A2 (nx8222)) ;
    or03 ix7516 (.Y (nx7515), .A0 (RST), .A1 (nx7345), .A2 (nx8222)) ;
    or03 ix7522 (.Y (nx7521), .A0 (RST), .A1 (nx7351), .A2 (nx8224)) ;
    or03 ix7528 (.Y (nx7527), .A0 (RST), .A1 (nx7357), .A2 (nx8224)) ;
    or03 ix7534 (.Y (nx7533), .A0 (RST), .A1 (nx7363), .A2 (nx8224)) ;
    or03 ix7540 (.Y (nx7539), .A0 (RST), .A1 (nx7369), .A2 (nx8224)) ;
    or03 ix7546 (.Y (nx7545), .A0 (RST), .A1 (nx7375), .A2 (nx8224)) ;
    or03 ix7552 (.Y (nx7551), .A0 (RST), .A1 (nx7381), .A2 (nx8224)) ;
    or03 ix7702 (.Y (nx7701), .A0 (RST), .A1 (nx7459), .A2 (nx8312)) ;
    or03 ix7708 (.Y (nx7707), .A0 (RST), .A1 (nx7465), .A2 (nx8312)) ;
    or03 ix7714 (.Y (nx7713), .A0 (RST), .A1 (nx7471), .A2 (nx8312)) ;
    or03 ix7720 (.Y (nx7719), .A0 (RST), .A1 (nx7477), .A2 (nx8312)) ;
    or03 ix7726 (.Y (nx7725), .A0 (RST), .A1 (nx7483), .A2 (nx8312)) ;
    or03 ix7732 (.Y (nx7731), .A0 (RST), .A1 (nx7489), .A2 (nx8312)) ;
    or03 ix7738 (.Y (nx7737), .A0 (RST), .A1 (nx7495), .A2 (nx8312)) ;
    or03 ix7744 (.Y (nx7743), .A0 (RST), .A1 (nx7501), .A2 (nx8314)) ;
    or03 ix7750 (.Y (nx7749), .A0 (RST), .A1 (nx7507), .A2 (nx8314)) ;
    or03 ix7756 (.Y (nx7755), .A0 (RST), .A1 (nx7513), .A2 (nx8314)) ;
    or03 ix7762 (.Y (nx7761), .A0 (RST), .A1 (nx7519), .A2 (nx8314)) ;
    or03 ix7768 (.Y (nx7767), .A0 (RST), .A1 (nx7525), .A2 (nx8314)) ;
    or03 ix7774 (.Y (nx7773), .A0 (RST), .A1 (nx7531), .A2 (nx8314)) ;
    or03 ix7780 (.Y (nx7779), .A0 (RST), .A1 (nx7537), .A2 (nx8314)) ;
    or03 ix7786 (.Y (nx7785), .A0 (RST), .A1 (nx7543), .A2 (nx8226)) ;
    or03 ix7792 (.Y (nx7791), .A0 (RST), .A1 (nx7549), .A2 (nx8226)) ;
    or03 ix7798 (.Y (nx7797), .A0 (RST), .A1 (nx7555), .A2 (nx8226)) ;
    or03 ix7804 (.Y (nx7803), .A0 (RST), .A1 (nx7561), .A2 (nx8226)) ;
    or03 ix7810 (.Y (nx7809), .A0 (RST), .A1 (nx7567), .A2 (nx8226)) ;
    or03 ix7816 (.Y (nx7815), .A0 (RST), .A1 (nx7573), .A2 (nx8316)) ;
    or03 ix7822 (.Y (nx7821), .A0 (RST), .A1 (nx7579), .A2 (nx8318)) ;
    or03 ix7828 (.Y (nx7827), .A0 (RST), .A1 (nx7585), .A2 (nx8318)) ;
    or03 ix7834 (.Y (nx7833), .A0 (RST), .A1 (nx7591), .A2 (nx8318)) ;
    or03 ix7840 (.Y (nx7839), .A0 (RST), .A1 (nx7597), .A2 (nx8318)) ;
    or03 ix7846 (.Y (nx7845), .A0 (RST), .A1 (nx7603), .A2 (nx8318)) ;
    or03 ix7852 (.Y (nx7851), .A0 (RST), .A1 (nx7609), .A2 (nx8318)) ;
    or03 ix7858 (.Y (nx7857), .A0 (RST), .A1 (nx7615), .A2 (nx8318)) ;
    or03 ix7864 (.Y (nx7863), .A0 (RST), .A1 (nx7621), .A2 (nx8320)) ;
    or03 ix7870 (.Y (nx7869), .A0 (RST), .A1 (nx7627), .A2 (nx8320)) ;
    or03 ix7876 (.Y (nx7875), .A0 (RST), .A1 (nx7633), .A2 (nx8320)) ;
    or03 ix7882 (.Y (nx7881), .A0 (RST), .A1 (nx7639), .A2 (nx8320)) ;
    or03 ix7888 (.Y (nx7887), .A0 (RST), .A1 (nx7645), .A2 (nx8320)) ;
    or03 ix7894 (.Y (nx7893), .A0 (RST), .A1 (nx7651), .A2 (nx8320)) ;
    or03 ix7900 (.Y (nx7899), .A0 (RST), .A1 (nx7657), .A2 (nx8320)) ;
    or03 ix7906 (.Y (nx7905), .A0 (RST), .A1 (nx7663), .A2 (nx8228)) ;
    or03 ix7912 (.Y (nx7911), .A0 (RST), .A1 (nx7669), .A2 (nx8228)) ;
    or03 ix7918 (.Y (nx7917), .A0 (RST), .A1 (nx7675), .A2 (nx8228)) ;
    or03 ix7924 (.Y (nx7923), .A0 (RST), .A1 (nx7681), .A2 (nx8228)) ;
    or03 ix7930 (.Y (nx7929), .A0 (RST), .A1 (nx7687), .A2 (nx8228)) ;
    or03 ix7936 (.Y (nx7935), .A0 (RST), .A1 (nx7693), .A2 (nx8228)) ;
    inv02 ix8269 (.Y (nx8270), .A (nx8334)) ;
    inv02 ix8271 (.Y (nx8272), .A (nx8334)) ;
    inv02 ix8273 (.Y (nx8274), .A (nx8336)) ;
    inv02 ix8275 (.Y (nx8276), .A (nx8336)) ;
    inv02 ix8277 (.Y (nx8278), .A (nx8324)) ;
    inv02 ix8279 (.Y (nx8280), .A (nx8324)) ;
    inv02 ix8281 (.Y (nx8282), .A (nx8324)) ;
    inv02 ix8283 (.Y (nx8284), .A (nx8324)) ;
    inv02 ix8285 (.Y (nx8286), .A (nx8324)) ;
    inv02 ix8287 (.Y (nx8288), .A (nx8324)) ;
    inv02 ix8289 (.Y (nx8290), .A (nx8324)) ;
    inv02 ix8291 (.Y (nx8292), .A (nx8270)) ;
    inv02 ix8293 (.Y (nx8294), .A (nx8270)) ;
    inv02 ix8295 (.Y (nx8296), .A (nx8270)) ;
    inv02 ix8297 (.Y (nx8298), .A (nx8270)) ;
    inv02 ix8299 (.Y (nx8300), .A (nx8328)) ;
    inv02 ix8301 (.Y (nx8302), .A (nx8328)) ;
    inv02 ix8303 (.Y (nx8304), .A (nx8328)) ;
    inv02 ix8305 (.Y (nx8306), .A (nx8328)) ;
    inv02 ix8307 (.Y (nx8308), .A (nx8328)) ;
    inv02 ix8309 (.Y (nx8310), .A (nx8328)) ;
    inv02 ix8311 (.Y (nx8312), .A (nx8328)) ;
    inv02 ix8313 (.Y (nx8314), .A (nx8274)) ;
    inv02 ix8315 (.Y (nx8316), .A (nx8274)) ;
    inv02 ix8317 (.Y (nx8318), .A (nx8274)) ;
    inv02 ix8319 (.Y (nx8320), .A (nx8274)) ;
    inv02 ix8321 (.Y (nx8322), .A (nx8334)) ;
    inv02 ix8323 (.Y (nx8324), .A (nx8334)) ;
    inv02 ix8325 (.Y (nx8326), .A (nx8336)) ;
    inv02 ix8327 (.Y (nx8328), .A (nx8336)) ;
    inv01 ix8333 (.Y (nx8334), .A (nx84)) ;
    inv01 ix8335 (.Y (nx8336), .A (nx168)) ;
endmodule


module RAM_8_18 ( CLK, WR, Address, Din, Dout ) ;

    input CLK ;
    input WR ;
    input [17:0]Address ;
    input [7:0]Din ;
    output [39:0]Dout ;




endmodule


module accelerator ( CLK, RST, Start, FilterSize, Instr, FilterDin_0__0__7, 
                     FilterDin_0__0__6, FilterDin_0__0__5, FilterDin_0__0__4, 
                     FilterDin_0__0__3, FilterDin_0__0__2, FilterDin_0__0__1, 
                     FilterDin_0__0__0, FilterDin_0__1__7, FilterDin_0__1__6, 
                     FilterDin_0__1__5, FilterDin_0__1__4, FilterDin_0__1__3, 
                     FilterDin_0__1__2, FilterDin_0__1__1, FilterDin_0__1__0, 
                     FilterDin_0__2__7, FilterDin_0__2__6, FilterDin_0__2__5, 
                     FilterDin_0__2__4, FilterDin_0__2__3, FilterDin_0__2__2, 
                     FilterDin_0__2__1, FilterDin_0__2__0, FilterDin_0__3__7, 
                     FilterDin_0__3__6, FilterDin_0__3__5, FilterDin_0__3__4, 
                     FilterDin_0__3__3, FilterDin_0__3__2, FilterDin_0__3__1, 
                     FilterDin_0__3__0, FilterDin_0__4__7, FilterDin_0__4__6, 
                     FilterDin_0__4__5, FilterDin_0__4__4, FilterDin_0__4__3, 
                     FilterDin_0__4__2, FilterDin_0__4__1, FilterDin_0__4__0, 
                     FilterDin_1__0__7, FilterDin_1__0__6, FilterDin_1__0__5, 
                     FilterDin_1__0__4, FilterDin_1__0__3, FilterDin_1__0__2, 
                     FilterDin_1__0__1, FilterDin_1__0__0, FilterDin_1__1__7, 
                     FilterDin_1__1__6, FilterDin_1__1__5, FilterDin_1__1__4, 
                     FilterDin_1__1__3, FilterDin_1__1__2, FilterDin_1__1__1, 
                     FilterDin_1__1__0, FilterDin_1__2__7, FilterDin_1__2__6, 
                     FilterDin_1__2__5, FilterDin_1__2__4, FilterDin_1__2__3, 
                     FilterDin_1__2__2, FilterDin_1__2__1, FilterDin_1__2__0, 
                     FilterDin_1__3__7, FilterDin_1__3__6, FilterDin_1__3__5, 
                     FilterDin_1__3__4, FilterDin_1__3__3, FilterDin_1__3__2, 
                     FilterDin_1__3__1, FilterDin_1__3__0, FilterDin_1__4__7, 
                     FilterDin_1__4__6, FilterDin_1__4__5, FilterDin_1__4__4, 
                     FilterDin_1__4__3, FilterDin_1__4__2, FilterDin_1__4__1, 
                     FilterDin_1__4__0, FilterDin_2__0__7, FilterDin_2__0__6, 
                     FilterDin_2__0__5, FilterDin_2__0__4, FilterDin_2__0__3, 
                     FilterDin_2__0__2, FilterDin_2__0__1, FilterDin_2__0__0, 
                     FilterDin_2__1__7, FilterDin_2__1__6, FilterDin_2__1__5, 
                     FilterDin_2__1__4, FilterDin_2__1__3, FilterDin_2__1__2, 
                     FilterDin_2__1__1, FilterDin_2__1__0, FilterDin_2__2__7, 
                     FilterDin_2__2__6, FilterDin_2__2__5, FilterDin_2__2__4, 
                     FilterDin_2__2__3, FilterDin_2__2__2, FilterDin_2__2__1, 
                     FilterDin_2__2__0, FilterDin_2__3__7, FilterDin_2__3__6, 
                     FilterDin_2__3__5, FilterDin_2__3__4, FilterDin_2__3__3, 
                     FilterDin_2__3__2, FilterDin_2__3__1, FilterDin_2__3__0, 
                     FilterDin_2__4__7, FilterDin_2__4__6, FilterDin_2__4__5, 
                     FilterDin_2__4__4, FilterDin_2__4__3, FilterDin_2__4__2, 
                     FilterDin_2__4__1, FilterDin_2__4__0, FilterDin_3__0__7, 
                     FilterDin_3__0__6, FilterDin_3__0__5, FilterDin_3__0__4, 
                     FilterDin_3__0__3, FilterDin_3__0__2, FilterDin_3__0__1, 
                     FilterDin_3__0__0, FilterDin_3__1__7, FilterDin_3__1__6, 
                     FilterDin_3__1__5, FilterDin_3__1__4, FilterDin_3__1__3, 
                     FilterDin_3__1__2, FilterDin_3__1__1, FilterDin_3__1__0, 
                     FilterDin_3__2__7, FilterDin_3__2__6, FilterDin_3__2__5, 
                     FilterDin_3__2__4, FilterDin_3__2__3, FilterDin_3__2__2, 
                     FilterDin_3__2__1, FilterDin_3__2__0, FilterDin_3__3__7, 
                     FilterDin_3__3__6, FilterDin_3__3__5, FilterDin_3__3__4, 
                     FilterDin_3__3__3, FilterDin_3__3__2, FilterDin_3__3__1, 
                     FilterDin_3__3__0, FilterDin_3__4__7, FilterDin_3__4__6, 
                     FilterDin_3__4__5, FilterDin_3__4__4, FilterDin_3__4__3, 
                     FilterDin_3__4__2, FilterDin_3__4__1, FilterDin_3__4__0, 
                     FilterDin_4__0__7, FilterDin_4__0__6, FilterDin_4__0__5, 
                     FilterDin_4__0__4, FilterDin_4__0__3, FilterDin_4__0__2, 
                     FilterDin_4__0__1, FilterDin_4__0__0, FilterDin_4__1__7, 
                     FilterDin_4__1__6, FilterDin_4__1__5, FilterDin_4__1__4, 
                     FilterDin_4__1__3, FilterDin_4__1__2, FilterDin_4__1__1, 
                     FilterDin_4__1__0, FilterDin_4__2__7, FilterDin_4__2__6, 
                     FilterDin_4__2__5, FilterDin_4__2__4, FilterDin_4__2__3, 
                     FilterDin_4__2__2, FilterDin_4__2__1, FilterDin_4__2__0, 
                     FilterDin_4__3__7, FilterDin_4__3__6, FilterDin_4__3__5, 
                     FilterDin_4__3__4, FilterDin_4__3__3, FilterDin_4__3__2, 
                     FilterDin_4__3__1, FilterDin_4__3__0, FilterDin_4__4__7, 
                     FilterDin_4__4__6, FilterDin_4__4__5, FilterDin_4__4__4, 
                     FilterDin_4__4__3, FilterDin_4__4__2, FilterDin_4__4__1, 
                     FilterDin_4__4__0, WindowDin_0__0__7, WindowDin_0__0__6, 
                     WindowDin_0__0__5, WindowDin_0__0__4, WindowDin_0__0__3, 
                     WindowDin_0__0__2, WindowDin_0__0__1, WindowDin_0__0__0, 
                     WindowDin_0__1__7, WindowDin_0__1__6, WindowDin_0__1__5, 
                     WindowDin_0__1__4, WindowDin_0__1__3, WindowDin_0__1__2, 
                     WindowDin_0__1__1, WindowDin_0__1__0, WindowDin_0__2__7, 
                     WindowDin_0__2__6, WindowDin_0__2__5, WindowDin_0__2__4, 
                     WindowDin_0__2__3, WindowDin_0__2__2, WindowDin_0__2__1, 
                     WindowDin_0__2__0, WindowDin_0__3__7, WindowDin_0__3__6, 
                     WindowDin_0__3__5, WindowDin_0__3__4, WindowDin_0__3__3, 
                     WindowDin_0__3__2, WindowDin_0__3__1, WindowDin_0__3__0, 
                     WindowDin_0__4__7, WindowDin_0__4__6, WindowDin_0__4__5, 
                     WindowDin_0__4__4, WindowDin_0__4__3, WindowDin_0__4__2, 
                     WindowDin_0__4__1, WindowDin_0__4__0, WindowDin_1__0__7, 
                     WindowDin_1__0__6, WindowDin_1__0__5, WindowDin_1__0__4, 
                     WindowDin_1__0__3, WindowDin_1__0__2, WindowDin_1__0__1, 
                     WindowDin_1__0__0, WindowDin_1__1__7, WindowDin_1__1__6, 
                     WindowDin_1__1__5, WindowDin_1__1__4, WindowDin_1__1__3, 
                     WindowDin_1__1__2, WindowDin_1__1__1, WindowDin_1__1__0, 
                     WindowDin_1__2__7, WindowDin_1__2__6, WindowDin_1__2__5, 
                     WindowDin_1__2__4, WindowDin_1__2__3, WindowDin_1__2__2, 
                     WindowDin_1__2__1, WindowDin_1__2__0, WindowDin_1__3__7, 
                     WindowDin_1__3__6, WindowDin_1__3__5, WindowDin_1__3__4, 
                     WindowDin_1__3__3, WindowDin_1__3__2, WindowDin_1__3__1, 
                     WindowDin_1__3__0, WindowDin_1__4__7, WindowDin_1__4__6, 
                     WindowDin_1__4__5, WindowDin_1__4__4, WindowDin_1__4__3, 
                     WindowDin_1__4__2, WindowDin_1__4__1, WindowDin_1__4__0, 
                     WindowDin_2__0__7, WindowDin_2__0__6, WindowDin_2__0__5, 
                     WindowDin_2__0__4, WindowDin_2__0__3, WindowDin_2__0__2, 
                     WindowDin_2__0__1, WindowDin_2__0__0, WindowDin_2__1__7, 
                     WindowDin_2__1__6, WindowDin_2__1__5, WindowDin_2__1__4, 
                     WindowDin_2__1__3, WindowDin_2__1__2, WindowDin_2__1__1, 
                     WindowDin_2__1__0, WindowDin_2__2__7, WindowDin_2__2__6, 
                     WindowDin_2__2__5, WindowDin_2__2__4, WindowDin_2__2__3, 
                     WindowDin_2__2__2, WindowDin_2__2__1, WindowDin_2__2__0, 
                     WindowDin_2__3__7, WindowDin_2__3__6, WindowDin_2__3__5, 
                     WindowDin_2__3__4, WindowDin_2__3__3, WindowDin_2__3__2, 
                     WindowDin_2__3__1, WindowDin_2__3__0, WindowDin_2__4__7, 
                     WindowDin_2__4__6, WindowDin_2__4__5, WindowDin_2__4__4, 
                     WindowDin_2__4__3, WindowDin_2__4__2, WindowDin_2__4__1, 
                     WindowDin_2__4__0, WindowDin_3__0__7, WindowDin_3__0__6, 
                     WindowDin_3__0__5, WindowDin_3__0__4, WindowDin_3__0__3, 
                     WindowDin_3__0__2, WindowDin_3__0__1, WindowDin_3__0__0, 
                     WindowDin_3__1__7, WindowDin_3__1__6, WindowDin_3__1__5, 
                     WindowDin_3__1__4, WindowDin_3__1__3, WindowDin_3__1__2, 
                     WindowDin_3__1__1, WindowDin_3__1__0, WindowDin_3__2__7, 
                     WindowDin_3__2__6, WindowDin_3__2__5, WindowDin_3__2__4, 
                     WindowDin_3__2__3, WindowDin_3__2__2, WindowDin_3__2__1, 
                     WindowDin_3__2__0, WindowDin_3__3__7, WindowDin_3__3__6, 
                     WindowDin_3__3__5, WindowDin_3__3__4, WindowDin_3__3__3, 
                     WindowDin_3__3__2, WindowDin_3__3__1, WindowDin_3__3__0, 
                     WindowDin_3__4__7, WindowDin_3__4__6, WindowDin_3__4__5, 
                     WindowDin_3__4__4, WindowDin_3__4__3, WindowDin_3__4__2, 
                     WindowDin_3__4__1, WindowDin_3__4__0, WindowDin_4__0__7, 
                     WindowDin_4__0__6, WindowDin_4__0__5, WindowDin_4__0__4, 
                     WindowDin_4__0__3, WindowDin_4__0__2, WindowDin_4__0__1, 
                     WindowDin_4__0__0, WindowDin_4__1__7, WindowDin_4__1__6, 
                     WindowDin_4__1__5, WindowDin_4__1__4, WindowDin_4__1__3, 
                     WindowDin_4__1__2, WindowDin_4__1__1, WindowDin_4__1__0, 
                     WindowDin_4__2__7, WindowDin_4__2__6, WindowDin_4__2__5, 
                     WindowDin_4__2__4, WindowDin_4__2__3, WindowDin_4__2__2, 
                     WindowDin_4__2__1, WindowDin_4__2__0, WindowDin_4__3__7, 
                     WindowDin_4__3__6, WindowDin_4__3__5, WindowDin_4__3__4, 
                     WindowDin_4__3__3, WindowDin_4__3__2, WindowDin_4__3__1, 
                     WindowDin_4__3__0, WindowDin_4__4__7, WindowDin_4__4__6, 
                     WindowDin_4__4__5, WindowDin_4__4__4, WindowDin_4__4__3, 
                     WindowDin_4__4__2, WindowDin_4__4__1, WindowDin_4__4__0, 
                     Done, Result ) ;

    input CLK ;
    input RST ;
    input Start ;
    input FilterSize ;
    input Instr ;
    input FilterDin_0__0__7 ;
    input FilterDin_0__0__6 ;
    input FilterDin_0__0__5 ;
    input FilterDin_0__0__4 ;
    input FilterDin_0__0__3 ;
    input FilterDin_0__0__2 ;
    input FilterDin_0__0__1 ;
    input FilterDin_0__0__0 ;
    input FilterDin_0__1__7 ;
    input FilterDin_0__1__6 ;
    input FilterDin_0__1__5 ;
    input FilterDin_0__1__4 ;
    input FilterDin_0__1__3 ;
    input FilterDin_0__1__2 ;
    input FilterDin_0__1__1 ;
    input FilterDin_0__1__0 ;
    input FilterDin_0__2__7 ;
    input FilterDin_0__2__6 ;
    input FilterDin_0__2__5 ;
    input FilterDin_0__2__4 ;
    input FilterDin_0__2__3 ;
    input FilterDin_0__2__2 ;
    input FilterDin_0__2__1 ;
    input FilterDin_0__2__0 ;
    input FilterDin_0__3__7 ;
    input FilterDin_0__3__6 ;
    input FilterDin_0__3__5 ;
    input FilterDin_0__3__4 ;
    input FilterDin_0__3__3 ;
    input FilterDin_0__3__2 ;
    input FilterDin_0__3__1 ;
    input FilterDin_0__3__0 ;
    input FilterDin_0__4__7 ;
    input FilterDin_0__4__6 ;
    input FilterDin_0__4__5 ;
    input FilterDin_0__4__4 ;
    input FilterDin_0__4__3 ;
    input FilterDin_0__4__2 ;
    input FilterDin_0__4__1 ;
    input FilterDin_0__4__0 ;
    input FilterDin_1__0__7 ;
    input FilterDin_1__0__6 ;
    input FilterDin_1__0__5 ;
    input FilterDin_1__0__4 ;
    input FilterDin_1__0__3 ;
    input FilterDin_1__0__2 ;
    input FilterDin_1__0__1 ;
    input FilterDin_1__0__0 ;
    input FilterDin_1__1__7 ;
    input FilterDin_1__1__6 ;
    input FilterDin_1__1__5 ;
    input FilterDin_1__1__4 ;
    input FilterDin_1__1__3 ;
    input FilterDin_1__1__2 ;
    input FilterDin_1__1__1 ;
    input FilterDin_1__1__0 ;
    input FilterDin_1__2__7 ;
    input FilterDin_1__2__6 ;
    input FilterDin_1__2__5 ;
    input FilterDin_1__2__4 ;
    input FilterDin_1__2__3 ;
    input FilterDin_1__2__2 ;
    input FilterDin_1__2__1 ;
    input FilterDin_1__2__0 ;
    input FilterDin_1__3__7 ;
    input FilterDin_1__3__6 ;
    input FilterDin_1__3__5 ;
    input FilterDin_1__3__4 ;
    input FilterDin_1__3__3 ;
    input FilterDin_1__3__2 ;
    input FilterDin_1__3__1 ;
    input FilterDin_1__3__0 ;
    input FilterDin_1__4__7 ;
    input FilterDin_1__4__6 ;
    input FilterDin_1__4__5 ;
    input FilterDin_1__4__4 ;
    input FilterDin_1__4__3 ;
    input FilterDin_1__4__2 ;
    input FilterDin_1__4__1 ;
    input FilterDin_1__4__0 ;
    input FilterDin_2__0__7 ;
    input FilterDin_2__0__6 ;
    input FilterDin_2__0__5 ;
    input FilterDin_2__0__4 ;
    input FilterDin_2__0__3 ;
    input FilterDin_2__0__2 ;
    input FilterDin_2__0__1 ;
    input FilterDin_2__0__0 ;
    input FilterDin_2__1__7 ;
    input FilterDin_2__1__6 ;
    input FilterDin_2__1__5 ;
    input FilterDin_2__1__4 ;
    input FilterDin_2__1__3 ;
    input FilterDin_2__1__2 ;
    input FilterDin_2__1__1 ;
    input FilterDin_2__1__0 ;
    input FilterDin_2__2__7 ;
    input FilterDin_2__2__6 ;
    input FilterDin_2__2__5 ;
    input FilterDin_2__2__4 ;
    input FilterDin_2__2__3 ;
    input FilterDin_2__2__2 ;
    input FilterDin_2__2__1 ;
    input FilterDin_2__2__0 ;
    input FilterDin_2__3__7 ;
    input FilterDin_2__3__6 ;
    input FilterDin_2__3__5 ;
    input FilterDin_2__3__4 ;
    input FilterDin_2__3__3 ;
    input FilterDin_2__3__2 ;
    input FilterDin_2__3__1 ;
    input FilterDin_2__3__0 ;
    input FilterDin_2__4__7 ;
    input FilterDin_2__4__6 ;
    input FilterDin_2__4__5 ;
    input FilterDin_2__4__4 ;
    input FilterDin_2__4__3 ;
    input FilterDin_2__4__2 ;
    input FilterDin_2__4__1 ;
    input FilterDin_2__4__0 ;
    input FilterDin_3__0__7 ;
    input FilterDin_3__0__6 ;
    input FilterDin_3__0__5 ;
    input FilterDin_3__0__4 ;
    input FilterDin_3__0__3 ;
    input FilterDin_3__0__2 ;
    input FilterDin_3__0__1 ;
    input FilterDin_3__0__0 ;
    input FilterDin_3__1__7 ;
    input FilterDin_3__1__6 ;
    input FilterDin_3__1__5 ;
    input FilterDin_3__1__4 ;
    input FilterDin_3__1__3 ;
    input FilterDin_3__1__2 ;
    input FilterDin_3__1__1 ;
    input FilterDin_3__1__0 ;
    input FilterDin_3__2__7 ;
    input FilterDin_3__2__6 ;
    input FilterDin_3__2__5 ;
    input FilterDin_3__2__4 ;
    input FilterDin_3__2__3 ;
    input FilterDin_3__2__2 ;
    input FilterDin_3__2__1 ;
    input FilterDin_3__2__0 ;
    input FilterDin_3__3__7 ;
    input FilterDin_3__3__6 ;
    input FilterDin_3__3__5 ;
    input FilterDin_3__3__4 ;
    input FilterDin_3__3__3 ;
    input FilterDin_3__3__2 ;
    input FilterDin_3__3__1 ;
    input FilterDin_3__3__0 ;
    input FilterDin_3__4__7 ;
    input FilterDin_3__4__6 ;
    input FilterDin_3__4__5 ;
    input FilterDin_3__4__4 ;
    input FilterDin_3__4__3 ;
    input FilterDin_3__4__2 ;
    input FilterDin_3__4__1 ;
    input FilterDin_3__4__0 ;
    input FilterDin_4__0__7 ;
    input FilterDin_4__0__6 ;
    input FilterDin_4__0__5 ;
    input FilterDin_4__0__4 ;
    input FilterDin_4__0__3 ;
    input FilterDin_4__0__2 ;
    input FilterDin_4__0__1 ;
    input FilterDin_4__0__0 ;
    input FilterDin_4__1__7 ;
    input FilterDin_4__1__6 ;
    input FilterDin_4__1__5 ;
    input FilterDin_4__1__4 ;
    input FilterDin_4__1__3 ;
    input FilterDin_4__1__2 ;
    input FilterDin_4__1__1 ;
    input FilterDin_4__1__0 ;
    input FilterDin_4__2__7 ;
    input FilterDin_4__2__6 ;
    input FilterDin_4__2__5 ;
    input FilterDin_4__2__4 ;
    input FilterDin_4__2__3 ;
    input FilterDin_4__2__2 ;
    input FilterDin_4__2__1 ;
    input FilterDin_4__2__0 ;
    input FilterDin_4__3__7 ;
    input FilterDin_4__3__6 ;
    input FilterDin_4__3__5 ;
    input FilterDin_4__3__4 ;
    input FilterDin_4__3__3 ;
    input FilterDin_4__3__2 ;
    input FilterDin_4__3__1 ;
    input FilterDin_4__3__0 ;
    input FilterDin_4__4__7 ;
    input FilterDin_4__4__6 ;
    input FilterDin_4__4__5 ;
    input FilterDin_4__4__4 ;
    input FilterDin_4__4__3 ;
    input FilterDin_4__4__2 ;
    input FilterDin_4__4__1 ;
    input FilterDin_4__4__0 ;
    input WindowDin_0__0__7 ;
    input WindowDin_0__0__6 ;
    input WindowDin_0__0__5 ;
    input WindowDin_0__0__4 ;
    input WindowDin_0__0__3 ;
    input WindowDin_0__0__2 ;
    input WindowDin_0__0__1 ;
    input WindowDin_0__0__0 ;
    input WindowDin_0__1__7 ;
    input WindowDin_0__1__6 ;
    input WindowDin_0__1__5 ;
    input WindowDin_0__1__4 ;
    input WindowDin_0__1__3 ;
    input WindowDin_0__1__2 ;
    input WindowDin_0__1__1 ;
    input WindowDin_0__1__0 ;
    input WindowDin_0__2__7 ;
    input WindowDin_0__2__6 ;
    input WindowDin_0__2__5 ;
    input WindowDin_0__2__4 ;
    input WindowDin_0__2__3 ;
    input WindowDin_0__2__2 ;
    input WindowDin_0__2__1 ;
    input WindowDin_0__2__0 ;
    input WindowDin_0__3__7 ;
    input WindowDin_0__3__6 ;
    input WindowDin_0__3__5 ;
    input WindowDin_0__3__4 ;
    input WindowDin_0__3__3 ;
    input WindowDin_0__3__2 ;
    input WindowDin_0__3__1 ;
    input WindowDin_0__3__0 ;
    input WindowDin_0__4__7 ;
    input WindowDin_0__4__6 ;
    input WindowDin_0__4__5 ;
    input WindowDin_0__4__4 ;
    input WindowDin_0__4__3 ;
    input WindowDin_0__4__2 ;
    input WindowDin_0__4__1 ;
    input WindowDin_0__4__0 ;
    input WindowDin_1__0__7 ;
    input WindowDin_1__0__6 ;
    input WindowDin_1__0__5 ;
    input WindowDin_1__0__4 ;
    input WindowDin_1__0__3 ;
    input WindowDin_1__0__2 ;
    input WindowDin_1__0__1 ;
    input WindowDin_1__0__0 ;
    input WindowDin_1__1__7 ;
    input WindowDin_1__1__6 ;
    input WindowDin_1__1__5 ;
    input WindowDin_1__1__4 ;
    input WindowDin_1__1__3 ;
    input WindowDin_1__1__2 ;
    input WindowDin_1__1__1 ;
    input WindowDin_1__1__0 ;
    input WindowDin_1__2__7 ;
    input WindowDin_1__2__6 ;
    input WindowDin_1__2__5 ;
    input WindowDin_1__2__4 ;
    input WindowDin_1__2__3 ;
    input WindowDin_1__2__2 ;
    input WindowDin_1__2__1 ;
    input WindowDin_1__2__0 ;
    input WindowDin_1__3__7 ;
    input WindowDin_1__3__6 ;
    input WindowDin_1__3__5 ;
    input WindowDin_1__3__4 ;
    input WindowDin_1__3__3 ;
    input WindowDin_1__3__2 ;
    input WindowDin_1__3__1 ;
    input WindowDin_1__3__0 ;
    input WindowDin_1__4__7 ;
    input WindowDin_1__4__6 ;
    input WindowDin_1__4__5 ;
    input WindowDin_1__4__4 ;
    input WindowDin_1__4__3 ;
    input WindowDin_1__4__2 ;
    input WindowDin_1__4__1 ;
    input WindowDin_1__4__0 ;
    input WindowDin_2__0__7 ;
    input WindowDin_2__0__6 ;
    input WindowDin_2__0__5 ;
    input WindowDin_2__0__4 ;
    input WindowDin_2__0__3 ;
    input WindowDin_2__0__2 ;
    input WindowDin_2__0__1 ;
    input WindowDin_2__0__0 ;
    input WindowDin_2__1__7 ;
    input WindowDin_2__1__6 ;
    input WindowDin_2__1__5 ;
    input WindowDin_2__1__4 ;
    input WindowDin_2__1__3 ;
    input WindowDin_2__1__2 ;
    input WindowDin_2__1__1 ;
    input WindowDin_2__1__0 ;
    input WindowDin_2__2__7 ;
    input WindowDin_2__2__6 ;
    input WindowDin_2__2__5 ;
    input WindowDin_2__2__4 ;
    input WindowDin_2__2__3 ;
    input WindowDin_2__2__2 ;
    input WindowDin_2__2__1 ;
    input WindowDin_2__2__0 ;
    input WindowDin_2__3__7 ;
    input WindowDin_2__3__6 ;
    input WindowDin_2__3__5 ;
    input WindowDin_2__3__4 ;
    input WindowDin_2__3__3 ;
    input WindowDin_2__3__2 ;
    input WindowDin_2__3__1 ;
    input WindowDin_2__3__0 ;
    input WindowDin_2__4__7 ;
    input WindowDin_2__4__6 ;
    input WindowDin_2__4__5 ;
    input WindowDin_2__4__4 ;
    input WindowDin_2__4__3 ;
    input WindowDin_2__4__2 ;
    input WindowDin_2__4__1 ;
    input WindowDin_2__4__0 ;
    input WindowDin_3__0__7 ;
    input WindowDin_3__0__6 ;
    input WindowDin_3__0__5 ;
    input WindowDin_3__0__4 ;
    input WindowDin_3__0__3 ;
    input WindowDin_3__0__2 ;
    input WindowDin_3__0__1 ;
    input WindowDin_3__0__0 ;
    input WindowDin_3__1__7 ;
    input WindowDin_3__1__6 ;
    input WindowDin_3__1__5 ;
    input WindowDin_3__1__4 ;
    input WindowDin_3__1__3 ;
    input WindowDin_3__1__2 ;
    input WindowDin_3__1__1 ;
    input WindowDin_3__1__0 ;
    input WindowDin_3__2__7 ;
    input WindowDin_3__2__6 ;
    input WindowDin_3__2__5 ;
    input WindowDin_3__2__4 ;
    input WindowDin_3__2__3 ;
    input WindowDin_3__2__2 ;
    input WindowDin_3__2__1 ;
    input WindowDin_3__2__0 ;
    input WindowDin_3__3__7 ;
    input WindowDin_3__3__6 ;
    input WindowDin_3__3__5 ;
    input WindowDin_3__3__4 ;
    input WindowDin_3__3__3 ;
    input WindowDin_3__3__2 ;
    input WindowDin_3__3__1 ;
    input WindowDin_3__3__0 ;
    input WindowDin_3__4__7 ;
    input WindowDin_3__4__6 ;
    input WindowDin_3__4__5 ;
    input WindowDin_3__4__4 ;
    input WindowDin_3__4__3 ;
    input WindowDin_3__4__2 ;
    input WindowDin_3__4__1 ;
    input WindowDin_3__4__0 ;
    input WindowDin_4__0__7 ;
    input WindowDin_4__0__6 ;
    input WindowDin_4__0__5 ;
    input WindowDin_4__0__4 ;
    input WindowDin_4__0__3 ;
    input WindowDin_4__0__2 ;
    input WindowDin_4__0__1 ;
    input WindowDin_4__0__0 ;
    input WindowDin_4__1__7 ;
    input WindowDin_4__1__6 ;
    input WindowDin_4__1__5 ;
    input WindowDin_4__1__4 ;
    input WindowDin_4__1__3 ;
    input WindowDin_4__1__2 ;
    input WindowDin_4__1__1 ;
    input WindowDin_4__1__0 ;
    input WindowDin_4__2__7 ;
    input WindowDin_4__2__6 ;
    input WindowDin_4__2__5 ;
    input WindowDin_4__2__4 ;
    input WindowDin_4__2__3 ;
    input WindowDin_4__2__2 ;
    input WindowDin_4__2__1 ;
    input WindowDin_4__2__0 ;
    input WindowDin_4__3__7 ;
    input WindowDin_4__3__6 ;
    input WindowDin_4__3__5 ;
    input WindowDin_4__3__4 ;
    input WindowDin_4__3__3 ;
    input WindowDin_4__3__2 ;
    input WindowDin_4__3__1 ;
    input WindowDin_4__3__0 ;
    input WindowDin_4__4__7 ;
    input WindowDin_4__4__6 ;
    input WindowDin_4__4__5 ;
    input WindowDin_4__4__4 ;
    input WindowDin_4__4__3 ;
    input WindowDin_4__4__2 ;
    input WindowDin_4__4__1 ;
    input WindowDin_4__4__0 ;
    output Done ;
    output [7:0]Result ;

    wire LoopingAndResultNotReady, L1FirstOperands_0__15, L1FirstOperands_0__14, 
         L1FirstOperands_0__13, L1FirstOperands_0__12, L1FirstOperands_0__11, 
         L1FirstOperands_0__10, L1FirstOperands_0__9, L1FirstOperands_0__8, 
         L1FirstOperands_0__7, L1FirstOperands_0__6, L1FirstOperands_0__5, 
         L1FirstOperands_0__4, L1FirstOperands_0__3, L1FirstOperands_0__2, 
         L1FirstOperands_0__1, L1FirstOperands_0__0, L1FirstOperands_2__15, 
         L1FirstOperands_2__14, L1FirstOperands_2__13, L1FirstOperands_2__12, 
         L1FirstOperands_2__11, L1FirstOperands_2__10, L1FirstOperands_2__9, 
         L1FirstOperands_2__8, L1FirstOperands_2__7, L1FirstOperands_2__6, 
         L1FirstOperands_2__5, L1FirstOperands_2__4, L1FirstOperands_2__3, 
         L1FirstOperands_2__2, L1FirstOperands_2__1, L1FirstOperands_2__0, 
         L1FirstOperands_3__15, L1FirstOperands_3__14, L1FirstOperands_3__13, 
         L1FirstOperands_3__12, L1FirstOperands_3__11, L1FirstOperands_3__10, 
         L1FirstOperands_3__9, L1FirstOperands_3__8, L1FirstOperands_3__7, 
         L1FirstOperands_3__6, L1FirstOperands_3__5, L1FirstOperands_3__4, 
         L1FirstOperands_3__3, L1FirstOperands_3__2, L1FirstOperands_3__1, 
         L1FirstOperands_3__0, L1FirstOperands_4__15, L1FirstOperands_4__14, 
         L1FirstOperands_4__13, L1FirstOperands_4__12, L1FirstOperands_4__11, 
         L1FirstOperands_4__10, L1FirstOperands_4__9, L1FirstOperands_4__8, 
         L1FirstOperands_4__7, L1FirstOperands_4__6, L1FirstOperands_4__5, 
         L1FirstOperands_4__4, L1FirstOperands_4__3, L1FirstOperands_4__2, 
         L1FirstOperands_4__1, L1FirstOperands_4__0, L1FirstOperands_6__15, 
         L1FirstOperands_6__14, L1FirstOperands_6__13, L1FirstOperands_6__12, 
         L1FirstOperands_6__11, L1FirstOperands_6__10, L1FirstOperands_6__9, 
         L1FirstOperands_6__8, L1FirstOperands_6__7, L1FirstOperands_6__6, 
         L1FirstOperands_6__5, L1FirstOperands_6__4, L1FirstOperands_6__3, 
         L1FirstOperands_6__2, L1FirstOperands_6__1, L1FirstOperands_6__0, 
         L1FirstOperands_7__15, L1FirstOperands_7__14, L1FirstOperands_7__13, 
         L1FirstOperands_7__12, L1FirstOperands_7__11, L1FirstOperands_7__10, 
         L1FirstOperands_7__9, L1FirstOperands_7__8, L1FirstOperands_7__7, 
         L1FirstOperands_7__6, L1FirstOperands_7__5, L1FirstOperands_7__4, 
         L1FirstOperands_7__3, L1FirstOperands_7__2, L1FirstOperands_7__1, 
         L1FirstOperands_7__0, L1FirstOperands_8__15, L1FirstOperands_8__14, 
         L1FirstOperands_8__13, L1FirstOperands_8__12, L1FirstOperands_8__11, 
         L1FirstOperands_8__10, L1FirstOperands_8__9, L1FirstOperands_8__8, 
         L1FirstOperands_8__7, L1FirstOperands_8__6, L1FirstOperands_8__5, 
         L1FirstOperands_8__4, L1FirstOperands_8__3, L1FirstOperands_8__2, 
         L1FirstOperands_8__1, L1FirstOperands_8__0, L1FirstOperands_10__15, 
         L1FirstOperands_10__14, L1FirstOperands_10__13, L1FirstOperands_10__12, 
         L1FirstOperands_10__11, L1FirstOperands_10__10, L1FirstOperands_10__9, 
         L1FirstOperands_10__8, L1FirstOperands_10__7, L1FirstOperands_10__6, 
         L1FirstOperands_10__5, L1FirstOperands_10__4, L1FirstOperands_10__3, 
         L1FirstOperands_10__2, L1FirstOperands_10__1, L1FirstOperands_10__0, 
         L1FirstOperands_11__15, L1FirstOperands_11__14, L1FirstOperands_11__13, 
         L1FirstOperands_11__12, L1FirstOperands_11__11, L1FirstOperands_11__10, 
         L1FirstOperands_11__9, L1FirstOperands_11__8, L1FirstOperands_11__7, 
         L1FirstOperands_11__6, L1FirstOperands_11__5, L1FirstOperands_11__4, 
         L1FirstOperands_11__3, L1FirstOperands_11__2, L1FirstOperands_11__1, 
         L1FirstOperands_11__0, L1ResultsLarge_0__16, L1ResultsLarge_0__15, 
         L1ResultsLarge_0__14, L1ResultsLarge_0__13, L1ResultsLarge_0__12, 
         L1ResultsLarge_0__11, L1ResultsLarge_0__10, L1ResultsLarge_0__9, 
         L1ResultsLarge_0__8, L1ResultsLarge_0__7, L1ResultsLarge_0__6, 
         L1ResultsLarge_0__5, L1ResultsLarge_0__4, L1ResultsLarge_0__3, 
         L1ResultsLarge_0__2, L1ResultsLarge_0__1, L1ResultsLarge_0__0, 
         L1ResultsLarge_1__16, L1ResultsLarge_1__15, L1ResultsLarge_1__14, 
         L1ResultsLarge_1__13, L1ResultsLarge_1__12, L1ResultsLarge_1__11, 
         L1ResultsLarge_1__10, L1ResultsLarge_1__9, L1ResultsLarge_1__8, 
         L1ResultsLarge_1__7, L1ResultsLarge_1__6, L1ResultsLarge_1__5, 
         L1ResultsLarge_1__4, L1ResultsLarge_1__3, L1ResultsLarge_1__2, 
         L1ResultsLarge_1__1, L1ResultsLarge_1__0, L1ResultsLarge_2__16, 
         L1ResultsLarge_2__15, L1ResultsLarge_2__14, L1ResultsLarge_2__13, 
         L1ResultsLarge_2__12, L1ResultsLarge_2__11, L1ResultsLarge_2__10, 
         L1ResultsLarge_2__9, L1ResultsLarge_2__8, L1ResultsLarge_2__7, 
         L1ResultsLarge_2__6, L1ResultsLarge_2__5, L1ResultsLarge_2__4, 
         L1ResultsLarge_2__3, L1ResultsLarge_2__2, L1ResultsLarge_2__1, 
         L1ResultsLarge_2__0, L1ResultsLarge_3__16, L1ResultsLarge_3__15, 
         L1ResultsLarge_3__14, L1ResultsLarge_3__13, L1ResultsLarge_3__12, 
         L1ResultsLarge_3__11, L1ResultsLarge_3__10, L1ResultsLarge_3__9, 
         L1ResultsLarge_3__8, L1ResultsLarge_3__7, L1ResultsLarge_3__6, 
         L1ResultsLarge_3__5, L1ResultsLarge_3__4, L1ResultsLarge_3__3, 
         L1ResultsLarge_3__2, L1ResultsLarge_3__1, L1ResultsLarge_3__0, 
         L1ResultsLarge_4__16, L1ResultsLarge_4__15, L1ResultsLarge_4__14, 
         L1ResultsLarge_4__13, L1ResultsLarge_4__12, L1ResultsLarge_4__11, 
         L1ResultsLarge_4__10, L1ResultsLarge_4__9, L1ResultsLarge_4__8, 
         L1ResultsLarge_4__7, L1ResultsLarge_4__6, L1ResultsLarge_4__5, 
         L1ResultsLarge_4__4, L1ResultsLarge_4__3, L1ResultsLarge_4__2, 
         L1ResultsLarge_4__1, L1ResultsLarge_4__0, L1ResultsLarge_5__16, 
         L1ResultsLarge_5__15, L1ResultsLarge_5__14, L1ResultsLarge_5__13, 
         L1ResultsLarge_5__12, L1ResultsLarge_5__11, L1ResultsLarge_5__10, 
         L1ResultsLarge_5__9, L1ResultsLarge_5__8, L1ResultsLarge_5__7, 
         L1ResultsLarge_5__6, L1ResultsLarge_5__5, L1ResultsLarge_5__4, 
         L1ResultsLarge_5__3, L1ResultsLarge_5__2, L1ResultsLarge_5__1, 
         L1ResultsLarge_5__0, L1ResultsLarge_6__16, L1ResultsLarge_6__15, 
         L1ResultsLarge_6__14, L1ResultsLarge_6__13, L1ResultsLarge_6__12, 
         L1ResultsLarge_6__11, L1ResultsLarge_6__10, L1ResultsLarge_6__9, 
         L1ResultsLarge_6__8, L1ResultsLarge_6__7, L1ResultsLarge_6__6, 
         L1ResultsLarge_6__5, L1ResultsLarge_6__4, L1ResultsLarge_6__3, 
         L1ResultsLarge_6__2, L1ResultsLarge_6__1, L1ResultsLarge_6__0, 
         L1ResultsLarge_7__16, L1ResultsLarge_7__15, L1ResultsLarge_7__14, 
         L1ResultsLarge_7__13, L1ResultsLarge_7__12, L1ResultsLarge_7__11, 
         L1ResultsLarge_7__10, L1ResultsLarge_7__9, L1ResultsLarge_7__8, 
         L1ResultsLarge_7__7, L1ResultsLarge_7__6, L1ResultsLarge_7__5, 
         L1ResultsLarge_7__4, L1ResultsLarge_7__3, L1ResultsLarge_7__2, 
         L1ResultsLarge_7__1, L1ResultsLarge_7__0, L1ResultsLarge_8__16, 
         L1ResultsLarge_8__15, L1ResultsLarge_8__14, L1ResultsLarge_8__13, 
         L1ResultsLarge_8__12, L1ResultsLarge_8__11, L1ResultsLarge_8__10, 
         L1ResultsLarge_8__9, L1ResultsLarge_8__8, L1ResultsLarge_8__7, 
         L1ResultsLarge_8__6, L1ResultsLarge_8__5, L1ResultsLarge_8__4, 
         L1ResultsLarge_8__3, L1ResultsLarge_8__2, L1ResultsLarge_8__1, 
         L1ResultsLarge_8__0, L1ResultsLarge_9__16, L1ResultsLarge_9__15, 
         L1ResultsLarge_9__14, L1ResultsLarge_9__13, L1ResultsLarge_9__12, 
         L1ResultsLarge_9__11, L1ResultsLarge_9__10, L1ResultsLarge_9__9, 
         L1ResultsLarge_9__8, L1ResultsLarge_9__7, L1ResultsLarge_9__6, 
         L1ResultsLarge_9__5, L1ResultsLarge_9__4, L1ResultsLarge_9__3, 
         L1ResultsLarge_9__2, L1ResultsLarge_9__1, L1ResultsLarge_9__0, 
         L1ResultsLarge_10__16, L1ResultsLarge_10__15, L1ResultsLarge_10__14, 
         L1ResultsLarge_10__13, L1ResultsLarge_10__12, L1ResultsLarge_10__11, 
         L1ResultsLarge_10__10, L1ResultsLarge_10__9, L1ResultsLarge_10__8, 
         L1ResultsLarge_10__7, L1ResultsLarge_10__6, L1ResultsLarge_10__5, 
         L1ResultsLarge_10__4, L1ResultsLarge_10__3, L1ResultsLarge_10__2, 
         L1ResultsLarge_10__1, L1ResultsLarge_10__0, L1ResultsLarge_11__16, 
         L1ResultsLarge_11__15, L1ResultsLarge_11__14, L1ResultsLarge_11__13, 
         L1ResultsLarge_11__12, L1ResultsLarge_11__11, L1ResultsLarge_11__10, 
         L1ResultsLarge_11__9, L1ResultsLarge_11__8, L1ResultsLarge_11__7, 
         L1ResultsLarge_11__6, L1ResultsLarge_11__5, L1ResultsLarge_11__4, 
         L1ResultsLarge_11__3, L1ResultsLarge_11__2, L1ResultsLarge_11__1, 
         L1ResultsLarge_11__0, L2ResultsLarge_0__16, L2ResultsLarge_0__15, 
         L2ResultsLarge_0__14, L2ResultsLarge_0__13, L2ResultsLarge_0__12, 
         L2ResultsLarge_0__11, L2ResultsLarge_0__10, L2ResultsLarge_0__9, 
         L2ResultsLarge_0__8, L2ResultsLarge_0__7, L2ResultsLarge_0__6, 
         L2ResultsLarge_0__5, L2ResultsLarge_0__4, L2ResultsLarge_0__3, 
         L2ResultsLarge_0__2, L2ResultsLarge_0__1, L2ResultsLarge_0__0, 
         L2ResultsLarge_1__16, L2ResultsLarge_1__15, L2ResultsLarge_1__14, 
         L2ResultsLarge_1__13, L2ResultsLarge_1__12, L2ResultsLarge_1__11, 
         L2ResultsLarge_1__10, L2ResultsLarge_1__9, L2ResultsLarge_1__8, 
         L2ResultsLarge_1__7, L2ResultsLarge_1__6, L2ResultsLarge_1__5, 
         L2ResultsLarge_1__4, L2ResultsLarge_1__3, L2ResultsLarge_1__2, 
         L2ResultsLarge_1__1, L2ResultsLarge_1__0, L2ResultsLarge_2__16, 
         L2ResultsLarge_2__15, L2ResultsLarge_2__14, L2ResultsLarge_2__13, 
         L2ResultsLarge_2__12, L2ResultsLarge_2__11, L2ResultsLarge_2__10, 
         L2ResultsLarge_2__9, L2ResultsLarge_2__8, L2ResultsLarge_2__7, 
         L2ResultsLarge_2__6, L2ResultsLarge_2__5, L2ResultsLarge_2__4, 
         L2ResultsLarge_2__3, L2ResultsLarge_2__2, L2ResultsLarge_2__1, 
         L2ResultsLarge_2__0, L2ResultsLarge_3__16, L2ResultsLarge_3__15, 
         L2ResultsLarge_3__14, L2ResultsLarge_3__13, L2ResultsLarge_3__12, 
         L2ResultsLarge_3__11, L2ResultsLarge_3__10, L2ResultsLarge_3__9, 
         L2ResultsLarge_3__8, L2ResultsLarge_3__7, L2ResultsLarge_3__6, 
         L2ResultsLarge_3__5, L2ResultsLarge_3__4, L2ResultsLarge_3__3, 
         L2ResultsLarge_3__2, L2ResultsLarge_3__1, L2ResultsLarge_3__0, 
         L2ResultsLarge_4__16, L2ResultsLarge_4__15, L2ResultsLarge_4__14, 
         L2ResultsLarge_4__13, L2ResultsLarge_4__12, L2ResultsLarge_4__11, 
         L2ResultsLarge_4__10, L2ResultsLarge_4__9, L2ResultsLarge_4__8, 
         L2ResultsLarge_4__7, L2ResultsLarge_4__6, L2ResultsLarge_4__5, 
         L2ResultsLarge_4__4, L2ResultsLarge_4__3, L2ResultsLarge_4__2, 
         L2ResultsLarge_4__1, L2ResultsLarge_4__0, L2ResultsLarge_5__16, 
         L2ResultsLarge_5__15, L2ResultsLarge_5__14, L2ResultsLarge_5__13, 
         L2ResultsLarge_5__12, L2ResultsLarge_5__11, L2ResultsLarge_5__10, 
         L2ResultsLarge_5__9, L2ResultsLarge_5__8, L2ResultsLarge_5__7, 
         L2ResultsLarge_5__6, L2ResultsLarge_5__5, L2ResultsLarge_5__4, 
         L2ResultsLarge_5__3, L2ResultsLarge_5__2, L2ResultsLarge_5__1, 
         L2ResultsLarge_5__0, L3ResultsLarge_0__16, L3ResultsLarge_0__15, 
         L3ResultsLarge_0__14, L3ResultsLarge_0__13, L3ResultsLarge_0__12, 
         L3ResultsLarge_0__11, L3ResultsLarge_0__10, L3ResultsLarge_0__9, 
         L3ResultsLarge_0__8, L3ResultsLarge_0__7, L3ResultsLarge_0__6, 
         L3ResultsLarge_0__5, L3ResultsLarge_0__4, L3ResultsLarge_0__3, 
         L3ResultsLarge_0__2, L3ResultsLarge_0__1, L3ResultsLarge_0__0, 
         L3ResultsLarge_1__16, L3ResultsLarge_1__15, L3ResultsLarge_1__14, 
         L3ResultsLarge_1__13, L3ResultsLarge_1__12, L3ResultsLarge_1__11, 
         L3ResultsLarge_1__10, L3ResultsLarge_1__9, L3ResultsLarge_1__8, 
         L3ResultsLarge_1__7, L3ResultsLarge_1__6, L3ResultsLarge_1__5, 
         L3ResultsLarge_1__4, L3ResultsLarge_1__3, L3ResultsLarge_1__2, 
         L3ResultsLarge_1__1, L3ResultsLarge_1__0, L3ResultsLarge_2__16, 
         L3ResultsLarge_2__15, L3ResultsLarge_2__14, L3ResultsLarge_2__13, 
         L3ResultsLarge_2__12, L3ResultsLarge_2__11, L3ResultsLarge_2__10, 
         L3ResultsLarge_2__9, L3ResultsLarge_2__8, L3ResultsLarge_2__7, 
         L3ResultsLarge_2__6, L3ResultsLarge_2__5, L3ResultsLarge_2__4, 
         L3ResultsLarge_2__3, L3ResultsLarge_2__2, L3ResultsLarge_2__1, 
         L3ResultsLarge_2__0, L4ResultsLarge_0__16, L4ResultsLarge_0__15, 
         L4ResultsLarge_0__14, L4ResultsLarge_0__13, L4ResultsLarge_0__12, 
         L4ResultsLarge_0__11, L4ResultsLarge_0__10, L4ResultsLarge_0__9, 
         L4ResultsLarge_0__8, L4ResultsLarge_0__7, L4ResultsLarge_0__6, 
         L4ResultsLarge_0__5, L4ResultsLarge_0__4, L4ResultsLarge_0__3, 
         L4ResultsLarge_0__2, L4ResultsLarge_0__1, L4ResultsLarge_0__0, 
         L5FirstOperands_1__16, L5FirstOperands_1__15, L5FirstOperands_1__14, 
         L5FirstOperands_1__13, L5FirstOperands_1__12, L5FirstOperands_1__11, 
         L5FirstOperands_1__10, L5FirstOperands_1__9, L5FirstOperands_1__8, 
         L5FirstOperands_1__7, L5FirstOperands_1__6, L5FirstOperands_1__5, 
         L5FirstOperands_1__4, L5FirstOperands_1__3, L5FirstOperands_1__2, 
         L5FirstOperands_1__1, L5FirstOperands_1__0, 
         L1_0_L2_0_G1_MINI_ALU_OperationResult_15, 
         L1_0_L2_0_G1_MINI_ALU_OperationResult_14, 
         L1_0_L2_0_G1_MINI_ALU_OperationResult_13, 
         L1_0_L2_0_G1_MINI_ALU_OperationResult_12, 
         L1_0_L2_0_G1_MINI_ALU_OperationResult_11, 
         L1_0_L2_0_G1_MINI_ALU_OperationResult_10, 
         L1_0_L2_0_G1_MINI_ALU_OperationResult_9, 
         L1_0_L2_0_G1_MINI_ALU_OperationResult_8, 
         L1_0_L2_0_G1_MINI_ALU_OperationResult_7, 
         L1_0_L2_0_G1_MINI_ALU_OperationResult_6, 
         L1_0_L2_0_G1_MINI_ALU_OperationResult_5, 
         L1_0_L2_0_G1_MINI_ALU_OperationResult_4, 
         L1_0_L2_0_G1_MINI_ALU_OperationResult_3, 
         L1_0_L2_0_G1_MINI_ALU_OperationResult_2, 
         L1_0_L2_0_G1_MINI_ALU_OperationResult_1, 
         L1_0_L2_0_G1_MINI_ALU_OperationResult_0, 
         L1_0_L2_0_G1_MINI_ALU_BoothXORCheck, 
         L1_0_L2_0_G1_MINI_ALU_BoothOperand_16, 
         L1_0_L2_0_G1_MINI_ALU_BoothOperand_15, 
         L1_0_L2_0_G1_MINI_ALU_BoothOperand_14, 
         L1_0_L2_0_G1_MINI_ALU_BoothOperand_13, 
         L1_0_L2_0_G1_MINI_ALU_BoothOperand_12, 
         L1_0_L2_0_G1_MINI_ALU_BoothOperand_11, 
         L1_0_L2_0_G1_MINI_ALU_BoothOperand_10, 
         L1_0_L2_0_G1_MINI_ALU_BoothOperand_9, L1_0_L2_0_G1_MINI_ALU_BoothP_16, 
         L1_0_L2_0_G1_MINI_ALU_BoothP_15, L1_0_L2_0_G1_MINI_ALU_BoothP_14, 
         L1_0_L2_0_G1_MINI_ALU_BoothP_13, L1_0_L2_0_G1_MINI_ALU_BoothP_12, 
         L1_0_L2_0_G1_MINI_ALU_BoothP_11, L1_0_L2_0_G1_MINI_ALU_BoothP_10, 
         L1_0_L2_0_G1_MINI_ALU_BoothP_9, L1_0_L2_0_G1_MINI_ALU_BoothP_8, 
         L1_0_L2_0_G1_MINI_ALU_BoothP_7, L1_0_L2_0_G1_MINI_ALU_BoothP_6, 
         L1_0_L2_0_G1_MINI_ALU_BoothP_5, L1_0_L2_0_G1_MINI_ALU_BoothP_4, 
         L1_0_L2_0_G1_MINI_ALU_BoothP_3, L1_0_L2_0_G1_MINI_ALU_BoothP_2, 
         L1_0_L2_0_G1_MINI_ALU_BoothP_1, L1_0_L2_0_G1_MINI_ALU_BoothP_0, 
         L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_15, 
         L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_14, 
         L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_13, 
         L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_12, 
         L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_11, 
         L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_10, 
         L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_9, 
         L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_8, 
         L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_7, 
         L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_6, 
         L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_5, 
         L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_4, 
         L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_3, 
         L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_2, 
         L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_1, 
         L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_0, 
         L1_0_L2_1_G1_MINI_ALU_OperationResult_15, 
         L1_0_L2_1_G1_MINI_ALU_OperationResult_14, 
         L1_0_L2_1_G1_MINI_ALU_OperationResult_13, 
         L1_0_L2_1_G1_MINI_ALU_OperationResult_12, 
         L1_0_L2_1_G1_MINI_ALU_OperationResult_11, 
         L1_0_L2_1_G1_MINI_ALU_OperationResult_10, 
         L1_0_L2_1_G1_MINI_ALU_OperationResult_9, 
         L1_0_L2_1_G1_MINI_ALU_OperationResult_8, 
         L1_0_L2_1_G1_MINI_ALU_OperationResult_7, 
         L1_0_L2_1_G1_MINI_ALU_OperationResult_6, 
         L1_0_L2_1_G1_MINI_ALU_OperationResult_5, 
         L1_0_L2_1_G1_MINI_ALU_OperationResult_4, 
         L1_0_L2_1_G1_MINI_ALU_OperationResult_3, 
         L1_0_L2_1_G1_MINI_ALU_OperationResult_2, 
         L1_0_L2_1_G1_MINI_ALU_OperationResult_1, 
         L1_0_L2_1_G1_MINI_ALU_OperationResult_0, 
         L1_0_L2_1_G1_MINI_ALU_BoothXORCheck, 
         L1_0_L2_1_G1_MINI_ALU_BoothOperand_16, 
         L1_0_L2_1_G1_MINI_ALU_BoothOperand_15, 
         L1_0_L2_1_G1_MINI_ALU_BoothOperand_14, 
         L1_0_L2_1_G1_MINI_ALU_BoothOperand_13, 
         L1_0_L2_1_G1_MINI_ALU_BoothOperand_12, 
         L1_0_L2_1_G1_MINI_ALU_BoothOperand_11, 
         L1_0_L2_1_G1_MINI_ALU_BoothOperand_10, 
         L1_0_L2_1_G1_MINI_ALU_BoothOperand_9, L1_0_L2_1_G1_MINI_ALU_BoothP_16, 
         L1_0_L2_1_G1_MINI_ALU_BoothP_15, L1_0_L2_1_G1_MINI_ALU_BoothP_14, 
         L1_0_L2_1_G1_MINI_ALU_BoothP_13, L1_0_L2_1_G1_MINI_ALU_BoothP_12, 
         L1_0_L2_1_G1_MINI_ALU_BoothP_11, L1_0_L2_1_G1_MINI_ALU_BoothP_10, 
         L1_0_L2_1_G1_MINI_ALU_BoothP_9, L1_0_L2_1_G1_MINI_ALU_BoothP_8, 
         L1_0_L2_1_G1_MINI_ALU_BoothP_7, L1_0_L2_1_G1_MINI_ALU_BoothP_6, 
         L1_0_L2_1_G1_MINI_ALU_BoothP_5, L1_0_L2_1_G1_MINI_ALU_BoothP_4, 
         L1_0_L2_1_G1_MINI_ALU_BoothP_3, L1_0_L2_1_G1_MINI_ALU_BoothP_2, 
         L1_0_L2_1_G1_MINI_ALU_BoothP_1, L1_0_L2_1_G1_MINI_ALU_BoothP_0, 
         L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_15, 
         L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_14, 
         L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_13, 
         L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_12, 
         L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_11, 
         L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_10, 
         L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_9, 
         L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_8, 
         L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_7, 
         L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_6, 
         L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_5, 
         L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_4, 
         L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_3, 
         L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_2, 
         L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_1, 
         L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_0, 
         L1_0_L2_2_G1_MINI_ALU_OperationResult_15, 
         L1_0_L2_2_G1_MINI_ALU_OperationResult_14, 
         L1_0_L2_2_G1_MINI_ALU_OperationResult_13, 
         L1_0_L2_2_G1_MINI_ALU_OperationResult_12, 
         L1_0_L2_2_G1_MINI_ALU_OperationResult_11, 
         L1_0_L2_2_G1_MINI_ALU_OperationResult_10, 
         L1_0_L2_2_G1_MINI_ALU_OperationResult_9, 
         L1_0_L2_2_G1_MINI_ALU_OperationResult_8, 
         L1_0_L2_2_G1_MINI_ALU_OperationResult_7, 
         L1_0_L2_2_G1_MINI_ALU_OperationResult_6, 
         L1_0_L2_2_G1_MINI_ALU_OperationResult_5, 
         L1_0_L2_2_G1_MINI_ALU_OperationResult_4, 
         L1_0_L2_2_G1_MINI_ALU_OperationResult_3, 
         L1_0_L2_2_G1_MINI_ALU_OperationResult_2, 
         L1_0_L2_2_G1_MINI_ALU_OperationResult_1, 
         L1_0_L2_2_G1_MINI_ALU_OperationResult_0, 
         L1_0_L2_2_G1_MINI_ALU_BoothXORCheck, 
         L1_0_L2_2_G1_MINI_ALU_BoothOperand_16, 
         L1_0_L2_2_G1_MINI_ALU_BoothOperand_15, 
         L1_0_L2_2_G1_MINI_ALU_BoothOperand_14, 
         L1_0_L2_2_G1_MINI_ALU_BoothOperand_13, 
         L1_0_L2_2_G1_MINI_ALU_BoothOperand_12, 
         L1_0_L2_2_G1_MINI_ALU_BoothOperand_11, 
         L1_0_L2_2_G1_MINI_ALU_BoothOperand_10, 
         L1_0_L2_2_G1_MINI_ALU_BoothOperand_9, L1_0_L2_2_G1_MINI_ALU_BoothP_16, 
         L1_0_L2_2_G1_MINI_ALU_BoothP_15, L1_0_L2_2_G1_MINI_ALU_BoothP_14, 
         L1_0_L2_2_G1_MINI_ALU_BoothP_13, L1_0_L2_2_G1_MINI_ALU_BoothP_12, 
         L1_0_L2_2_G1_MINI_ALU_BoothP_11, L1_0_L2_2_G1_MINI_ALU_BoothP_10, 
         L1_0_L2_2_G1_MINI_ALU_BoothP_9, L1_0_L2_2_G1_MINI_ALU_BoothP_8, 
         L1_0_L2_2_G1_MINI_ALU_BoothP_7, L1_0_L2_2_G1_MINI_ALU_BoothP_6, 
         L1_0_L2_2_G1_MINI_ALU_BoothP_5, L1_0_L2_2_G1_MINI_ALU_BoothP_4, 
         L1_0_L2_2_G1_MINI_ALU_BoothP_3, L1_0_L2_2_G1_MINI_ALU_BoothP_2, 
         L1_0_L2_2_G1_MINI_ALU_BoothP_1, L1_0_L2_2_G1_MINI_ALU_BoothP_0, 
         L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_15, 
         L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_14, 
         L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_13, 
         L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_12, 
         L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_11, 
         L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_10, 
         L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_9, 
         L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_8, 
         L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_7, 
         L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_6, 
         L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_5, 
         L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_4, 
         L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_3, 
         L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_2, 
         L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_1, 
         L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_0, 
         L1_0_L2_3_G1_MINI_ALU_OperationResult_15, 
         L1_0_L2_3_G1_MINI_ALU_OperationResult_14, 
         L1_0_L2_3_G1_MINI_ALU_OperationResult_13, 
         L1_0_L2_3_G1_MINI_ALU_OperationResult_12, 
         L1_0_L2_3_G1_MINI_ALU_OperationResult_11, 
         L1_0_L2_3_G1_MINI_ALU_OperationResult_10, 
         L1_0_L2_3_G1_MINI_ALU_OperationResult_9, 
         L1_0_L2_3_G1_MINI_ALU_OperationResult_8, 
         L1_0_L2_3_G1_MINI_ALU_OperationResult_7, 
         L1_0_L2_3_G1_MINI_ALU_OperationResult_6, 
         L1_0_L2_3_G1_MINI_ALU_OperationResult_5, 
         L1_0_L2_3_G1_MINI_ALU_OperationResult_4, 
         L1_0_L2_3_G1_MINI_ALU_OperationResult_3, 
         L1_0_L2_3_G1_MINI_ALU_OperationResult_2, 
         L1_0_L2_3_G1_MINI_ALU_OperationResult_1, 
         L1_0_L2_3_G1_MINI_ALU_OperationResult_0, 
         L1_0_L2_3_G1_MINI_ALU_BoothXORCheck, 
         L1_0_L2_3_G1_MINI_ALU_BoothOperand_16, 
         L1_0_L2_3_G1_MINI_ALU_BoothOperand_15, 
         L1_0_L2_3_G1_MINI_ALU_BoothOperand_14, 
         L1_0_L2_3_G1_MINI_ALU_BoothOperand_13, 
         L1_0_L2_3_G1_MINI_ALU_BoothOperand_12, 
         L1_0_L2_3_G1_MINI_ALU_BoothOperand_11, 
         L1_0_L2_3_G1_MINI_ALU_BoothOperand_10, 
         L1_0_L2_3_G1_MINI_ALU_BoothOperand_9, L1_0_L2_3_G1_MINI_ALU_BoothP_16, 
         L1_0_L2_3_G1_MINI_ALU_BoothP_15, L1_0_L2_3_G1_MINI_ALU_BoothP_14, 
         L1_0_L2_3_G1_MINI_ALU_BoothP_13, L1_0_L2_3_G1_MINI_ALU_BoothP_12, 
         L1_0_L2_3_G1_MINI_ALU_BoothP_11, L1_0_L2_3_G1_MINI_ALU_BoothP_10, 
         L1_0_L2_3_G1_MINI_ALU_BoothP_9, L1_0_L2_3_G1_MINI_ALU_BoothP_8, 
         L1_0_L2_3_G1_MINI_ALU_BoothP_7, L1_0_L2_3_G1_MINI_ALU_BoothP_6, 
         L1_0_L2_3_G1_MINI_ALU_BoothP_5, L1_0_L2_3_G1_MINI_ALU_BoothP_4, 
         L1_0_L2_3_G1_MINI_ALU_BoothP_3, L1_0_L2_3_G1_MINI_ALU_BoothP_2, 
         L1_0_L2_3_G1_MINI_ALU_BoothP_1, L1_0_L2_3_G1_MINI_ALU_BoothP_0, 
         L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_15, 
         L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_14, 
         L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_13, 
         L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_12, 
         L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_11, 
         L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_10, 
         L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_9, 
         L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_8, 
         L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_7, 
         L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_6, 
         L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_5, 
         L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_4, 
         L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_3, 
         L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_2, 
         L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_1, 
         L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_0, 
         L1_0_L2_4_G1_MINI_ALU_OperationResult_15, 
         L1_0_L2_4_G1_MINI_ALU_OperationResult_14, 
         L1_0_L2_4_G1_MINI_ALU_OperationResult_13, 
         L1_0_L2_4_G1_MINI_ALU_OperationResult_12, 
         L1_0_L2_4_G1_MINI_ALU_OperationResult_11, 
         L1_0_L2_4_G1_MINI_ALU_OperationResult_10, 
         L1_0_L2_4_G1_MINI_ALU_OperationResult_9, 
         L1_0_L2_4_G1_MINI_ALU_OperationResult_8, 
         L1_0_L2_4_G1_MINI_ALU_OperationResult_7, 
         L1_0_L2_4_G1_MINI_ALU_OperationResult_6, 
         L1_0_L2_4_G1_MINI_ALU_OperationResult_5, 
         L1_0_L2_4_G1_MINI_ALU_OperationResult_4, 
         L1_0_L2_4_G1_MINI_ALU_OperationResult_3, 
         L1_0_L2_4_G1_MINI_ALU_OperationResult_2, 
         L1_0_L2_4_G1_MINI_ALU_OperationResult_1, 
         L1_0_L2_4_G1_MINI_ALU_OperationResult_0, 
         L1_0_L2_4_G1_MINI_ALU_BoothXORCheck, 
         L1_0_L2_4_G1_MINI_ALU_BoothOperand_16, 
         L1_0_L2_4_G1_MINI_ALU_BoothOperand_15, 
         L1_0_L2_4_G1_MINI_ALU_BoothOperand_14, 
         L1_0_L2_4_G1_MINI_ALU_BoothOperand_13, 
         L1_0_L2_4_G1_MINI_ALU_BoothOperand_12, 
         L1_0_L2_4_G1_MINI_ALU_BoothOperand_11, 
         L1_0_L2_4_G1_MINI_ALU_BoothOperand_10, 
         L1_0_L2_4_G1_MINI_ALU_BoothOperand_9, L1_0_L2_4_G1_MINI_ALU_BoothP_16, 
         L1_0_L2_4_G1_MINI_ALU_BoothP_15, L1_0_L2_4_G1_MINI_ALU_BoothP_14, 
         L1_0_L2_4_G1_MINI_ALU_BoothP_13, L1_0_L2_4_G1_MINI_ALU_BoothP_12, 
         L1_0_L2_4_G1_MINI_ALU_BoothP_11, L1_0_L2_4_G1_MINI_ALU_BoothP_10, 
         L1_0_L2_4_G1_MINI_ALU_BoothP_9, L1_0_L2_4_G1_MINI_ALU_BoothP_8, 
         L1_0_L2_4_G1_MINI_ALU_BoothP_7, L1_0_L2_4_G1_MINI_ALU_BoothP_6, 
         L1_0_L2_4_G1_MINI_ALU_BoothP_5, L1_0_L2_4_G1_MINI_ALU_BoothP_4, 
         L1_0_L2_4_G1_MINI_ALU_BoothP_3, L1_0_L2_4_G1_MINI_ALU_BoothP_2, 
         L1_0_L2_4_G1_MINI_ALU_BoothP_1, L1_0_L2_4_G1_MINI_ALU_BoothP_0, 
         L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_15, 
         L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_14, 
         L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_13, 
         L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_12, 
         L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_11, 
         L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_10, 
         L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_9, 
         L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_8, 
         L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_7, 
         L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_6, 
         L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_5, 
         L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_4, 
         L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_3, 
         L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_2, 
         L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_1, 
         L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_0, 
         L1_1_L2_0_G1_MINI_ALU_OperationResult_15, 
         L1_1_L2_0_G1_MINI_ALU_OperationResult_14, 
         L1_1_L2_0_G1_MINI_ALU_OperationResult_13, 
         L1_1_L2_0_G1_MINI_ALU_OperationResult_12, 
         L1_1_L2_0_G1_MINI_ALU_OperationResult_11, 
         L1_1_L2_0_G1_MINI_ALU_OperationResult_10, 
         L1_1_L2_0_G1_MINI_ALU_OperationResult_9, 
         L1_1_L2_0_G1_MINI_ALU_OperationResult_8, 
         L1_1_L2_0_G1_MINI_ALU_OperationResult_7, 
         L1_1_L2_0_G1_MINI_ALU_OperationResult_6, 
         L1_1_L2_0_G1_MINI_ALU_OperationResult_5, 
         L1_1_L2_0_G1_MINI_ALU_OperationResult_4, 
         L1_1_L2_0_G1_MINI_ALU_OperationResult_3, 
         L1_1_L2_0_G1_MINI_ALU_OperationResult_2, 
         L1_1_L2_0_G1_MINI_ALU_OperationResult_1, 
         L1_1_L2_0_G1_MINI_ALU_OperationResult_0, 
         L1_1_L2_0_G1_MINI_ALU_BoothXORCheck, 
         L1_1_L2_0_G1_MINI_ALU_BoothOperand_16, 
         L1_1_L2_0_G1_MINI_ALU_BoothOperand_15, 
         L1_1_L2_0_G1_MINI_ALU_BoothOperand_14, 
         L1_1_L2_0_G1_MINI_ALU_BoothOperand_13, 
         L1_1_L2_0_G1_MINI_ALU_BoothOperand_12, 
         L1_1_L2_0_G1_MINI_ALU_BoothOperand_11, 
         L1_1_L2_0_G1_MINI_ALU_BoothOperand_10, 
         L1_1_L2_0_G1_MINI_ALU_BoothOperand_9, L1_1_L2_0_G1_MINI_ALU_BoothP_16, 
         L1_1_L2_0_G1_MINI_ALU_BoothP_15, L1_1_L2_0_G1_MINI_ALU_BoothP_14, 
         L1_1_L2_0_G1_MINI_ALU_BoothP_13, L1_1_L2_0_G1_MINI_ALU_BoothP_12, 
         L1_1_L2_0_G1_MINI_ALU_BoothP_11, L1_1_L2_0_G1_MINI_ALU_BoothP_10, 
         L1_1_L2_0_G1_MINI_ALU_BoothP_9, L1_1_L2_0_G1_MINI_ALU_BoothP_8, 
         L1_1_L2_0_G1_MINI_ALU_BoothP_7, L1_1_L2_0_G1_MINI_ALU_BoothP_6, 
         L1_1_L2_0_G1_MINI_ALU_BoothP_5, L1_1_L2_0_G1_MINI_ALU_BoothP_4, 
         L1_1_L2_0_G1_MINI_ALU_BoothP_3, L1_1_L2_0_G1_MINI_ALU_BoothP_2, 
         L1_1_L2_0_G1_MINI_ALU_BoothP_1, L1_1_L2_0_G1_MINI_ALU_BoothP_0, 
         L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_15, 
         L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_14, 
         L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_13, 
         L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_12, 
         L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_11, 
         L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_10, 
         L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_9, 
         L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_8, 
         L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_7, 
         L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_6, 
         L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_5, 
         L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_4, 
         L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_3, 
         L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_2, 
         L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_1, 
         L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_0, 
         L1_1_L2_1_G1_MINI_ALU_OperationResult_15, 
         L1_1_L2_1_G1_MINI_ALU_OperationResult_14, 
         L1_1_L2_1_G1_MINI_ALU_OperationResult_13, 
         L1_1_L2_1_G1_MINI_ALU_OperationResult_12, 
         L1_1_L2_1_G1_MINI_ALU_OperationResult_11, 
         L1_1_L2_1_G1_MINI_ALU_OperationResult_10, 
         L1_1_L2_1_G1_MINI_ALU_OperationResult_9, 
         L1_1_L2_1_G1_MINI_ALU_OperationResult_8, 
         L1_1_L2_1_G1_MINI_ALU_OperationResult_7, 
         L1_1_L2_1_G1_MINI_ALU_OperationResult_6, 
         L1_1_L2_1_G1_MINI_ALU_OperationResult_5, 
         L1_1_L2_1_G1_MINI_ALU_OperationResult_4, 
         L1_1_L2_1_G1_MINI_ALU_OperationResult_3, 
         L1_1_L2_1_G1_MINI_ALU_OperationResult_2, 
         L1_1_L2_1_G1_MINI_ALU_OperationResult_1, 
         L1_1_L2_1_G1_MINI_ALU_OperationResult_0, 
         L1_1_L2_1_G1_MINI_ALU_BoothXORCheck, 
         L1_1_L2_1_G1_MINI_ALU_BoothOperand_16, 
         L1_1_L2_1_G1_MINI_ALU_BoothOperand_15, 
         L1_1_L2_1_G1_MINI_ALU_BoothOperand_14, 
         L1_1_L2_1_G1_MINI_ALU_BoothOperand_13, 
         L1_1_L2_1_G1_MINI_ALU_BoothOperand_12, 
         L1_1_L2_1_G1_MINI_ALU_BoothOperand_11, 
         L1_1_L2_1_G1_MINI_ALU_BoothOperand_10, 
         L1_1_L2_1_G1_MINI_ALU_BoothOperand_9, L1_1_L2_1_G1_MINI_ALU_BoothP_16, 
         L1_1_L2_1_G1_MINI_ALU_BoothP_15, L1_1_L2_1_G1_MINI_ALU_BoothP_14, 
         L1_1_L2_1_G1_MINI_ALU_BoothP_13, L1_1_L2_1_G1_MINI_ALU_BoothP_12, 
         L1_1_L2_1_G1_MINI_ALU_BoothP_11, L1_1_L2_1_G1_MINI_ALU_BoothP_10, 
         L1_1_L2_1_G1_MINI_ALU_BoothP_9, L1_1_L2_1_G1_MINI_ALU_BoothP_8, 
         L1_1_L2_1_G1_MINI_ALU_BoothP_7, L1_1_L2_1_G1_MINI_ALU_BoothP_6, 
         L1_1_L2_1_G1_MINI_ALU_BoothP_5, L1_1_L2_1_G1_MINI_ALU_BoothP_4, 
         L1_1_L2_1_G1_MINI_ALU_BoothP_3, L1_1_L2_1_G1_MINI_ALU_BoothP_2, 
         L1_1_L2_1_G1_MINI_ALU_BoothP_1, L1_1_L2_1_G1_MINI_ALU_BoothP_0, 
         L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_15, 
         L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_14, 
         L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_13, 
         L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_12, 
         L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_11, 
         L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_10, 
         L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_9, 
         L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_8, 
         L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_7, 
         L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_6, 
         L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_5, 
         L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_4, 
         L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_3, 
         L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_2, 
         L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_1, 
         L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_0, 
         L1_1_L2_2_G1_MINI_ALU_OperationResult_15, 
         L1_1_L2_2_G1_MINI_ALU_OperationResult_14, 
         L1_1_L2_2_G1_MINI_ALU_OperationResult_13, 
         L1_1_L2_2_G1_MINI_ALU_OperationResult_12, 
         L1_1_L2_2_G1_MINI_ALU_OperationResult_11, 
         L1_1_L2_2_G1_MINI_ALU_OperationResult_10, 
         L1_1_L2_2_G1_MINI_ALU_OperationResult_9, 
         L1_1_L2_2_G1_MINI_ALU_OperationResult_8, 
         L1_1_L2_2_G1_MINI_ALU_OperationResult_7, 
         L1_1_L2_2_G1_MINI_ALU_OperationResult_6, 
         L1_1_L2_2_G1_MINI_ALU_OperationResult_5, 
         L1_1_L2_2_G1_MINI_ALU_OperationResult_4, 
         L1_1_L2_2_G1_MINI_ALU_OperationResult_3, 
         L1_1_L2_2_G1_MINI_ALU_OperationResult_2, 
         L1_1_L2_2_G1_MINI_ALU_OperationResult_1, 
         L1_1_L2_2_G1_MINI_ALU_OperationResult_0, 
         L1_1_L2_2_G1_MINI_ALU_BoothXORCheck, 
         L1_1_L2_2_G1_MINI_ALU_BoothOperand_16, 
         L1_1_L2_2_G1_MINI_ALU_BoothOperand_15, 
         L1_1_L2_2_G1_MINI_ALU_BoothOperand_14, 
         L1_1_L2_2_G1_MINI_ALU_BoothOperand_13, 
         L1_1_L2_2_G1_MINI_ALU_BoothOperand_12, 
         L1_1_L2_2_G1_MINI_ALU_BoothOperand_11, 
         L1_1_L2_2_G1_MINI_ALU_BoothOperand_10, 
         L1_1_L2_2_G1_MINI_ALU_BoothOperand_9, L1_1_L2_2_G1_MINI_ALU_BoothP_16, 
         L1_1_L2_2_G1_MINI_ALU_BoothP_15, L1_1_L2_2_G1_MINI_ALU_BoothP_14, 
         L1_1_L2_2_G1_MINI_ALU_BoothP_13, L1_1_L2_2_G1_MINI_ALU_BoothP_12, 
         L1_1_L2_2_G1_MINI_ALU_BoothP_11, L1_1_L2_2_G1_MINI_ALU_BoothP_10, 
         L1_1_L2_2_G1_MINI_ALU_BoothP_9, L1_1_L2_2_G1_MINI_ALU_BoothP_8, 
         L1_1_L2_2_G1_MINI_ALU_BoothP_7, L1_1_L2_2_G1_MINI_ALU_BoothP_6, 
         L1_1_L2_2_G1_MINI_ALU_BoothP_5, L1_1_L2_2_G1_MINI_ALU_BoothP_4, 
         L1_1_L2_2_G1_MINI_ALU_BoothP_3, L1_1_L2_2_G1_MINI_ALU_BoothP_2, 
         L1_1_L2_2_G1_MINI_ALU_BoothP_1, L1_1_L2_2_G1_MINI_ALU_BoothP_0, 
         L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_15, 
         L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_14, 
         L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_13, 
         L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_12, 
         L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_11, 
         L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_10, 
         L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_9, 
         L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_8, 
         L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_7, 
         L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_6, 
         L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_5, 
         L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_4, 
         L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_3, 
         L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_2, 
         L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_1, 
         L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_0, 
         L1_1_L2_3_G1_MINI_ALU_OperationResult_15, 
         L1_1_L2_3_G1_MINI_ALU_OperationResult_14, 
         L1_1_L2_3_G1_MINI_ALU_OperationResult_13, 
         L1_1_L2_3_G1_MINI_ALU_OperationResult_12, 
         L1_1_L2_3_G1_MINI_ALU_OperationResult_11, 
         L1_1_L2_3_G1_MINI_ALU_OperationResult_10, 
         L1_1_L2_3_G1_MINI_ALU_OperationResult_9, 
         L1_1_L2_3_G1_MINI_ALU_OperationResult_8, 
         L1_1_L2_3_G1_MINI_ALU_OperationResult_7, 
         L1_1_L2_3_G1_MINI_ALU_OperationResult_6, 
         L1_1_L2_3_G1_MINI_ALU_OperationResult_5, 
         L1_1_L2_3_G1_MINI_ALU_OperationResult_4, 
         L1_1_L2_3_G1_MINI_ALU_OperationResult_3, 
         L1_1_L2_3_G1_MINI_ALU_OperationResult_2, 
         L1_1_L2_3_G1_MINI_ALU_OperationResult_1, 
         L1_1_L2_3_G1_MINI_ALU_OperationResult_0, 
         L1_1_L2_3_G1_MINI_ALU_BoothXORCheck, 
         L1_1_L2_3_G1_MINI_ALU_BoothOperand_16, 
         L1_1_L2_3_G1_MINI_ALU_BoothOperand_15, 
         L1_1_L2_3_G1_MINI_ALU_BoothOperand_14, 
         L1_1_L2_3_G1_MINI_ALU_BoothOperand_13, 
         L1_1_L2_3_G1_MINI_ALU_BoothOperand_12, 
         L1_1_L2_3_G1_MINI_ALU_BoothOperand_11, 
         L1_1_L2_3_G1_MINI_ALU_BoothOperand_10, 
         L1_1_L2_3_G1_MINI_ALU_BoothOperand_9, L1_1_L2_3_G1_MINI_ALU_BoothP_16, 
         L1_1_L2_3_G1_MINI_ALU_BoothP_15, L1_1_L2_3_G1_MINI_ALU_BoothP_14, 
         L1_1_L2_3_G1_MINI_ALU_BoothP_13, L1_1_L2_3_G1_MINI_ALU_BoothP_12, 
         L1_1_L2_3_G1_MINI_ALU_BoothP_11, L1_1_L2_3_G1_MINI_ALU_BoothP_10, 
         L1_1_L2_3_G1_MINI_ALU_BoothP_9, L1_1_L2_3_G1_MINI_ALU_BoothP_8, 
         L1_1_L2_3_G1_MINI_ALU_BoothP_7, L1_1_L2_3_G1_MINI_ALU_BoothP_6, 
         L1_1_L2_3_G1_MINI_ALU_BoothP_5, L1_1_L2_3_G1_MINI_ALU_BoothP_4, 
         L1_1_L2_3_G1_MINI_ALU_BoothP_3, L1_1_L2_3_G1_MINI_ALU_BoothP_2, 
         L1_1_L2_3_G1_MINI_ALU_BoothP_1, L1_1_L2_3_G1_MINI_ALU_BoothP_0, 
         L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_15, 
         L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_14, 
         L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_13, 
         L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_12, 
         L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_11, 
         L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_10, 
         L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_9, 
         L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_8, 
         L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_7, 
         L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_6, 
         L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_5, 
         L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_4, 
         L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_3, 
         L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_2, 
         L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_1, 
         L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_0, 
         L1_1_L2_4_G1_MINI_ALU_OperationResult_15, 
         L1_1_L2_4_G1_MINI_ALU_OperationResult_14, 
         L1_1_L2_4_G1_MINI_ALU_OperationResult_13, 
         L1_1_L2_4_G1_MINI_ALU_OperationResult_12, 
         L1_1_L2_4_G1_MINI_ALU_OperationResult_11, 
         L1_1_L2_4_G1_MINI_ALU_OperationResult_10, 
         L1_1_L2_4_G1_MINI_ALU_OperationResult_9, 
         L1_1_L2_4_G1_MINI_ALU_OperationResult_8, 
         L1_1_L2_4_G1_MINI_ALU_OperationResult_7, 
         L1_1_L2_4_G1_MINI_ALU_OperationResult_6, 
         L1_1_L2_4_G1_MINI_ALU_OperationResult_5, 
         L1_1_L2_4_G1_MINI_ALU_OperationResult_4, 
         L1_1_L2_4_G1_MINI_ALU_OperationResult_3, 
         L1_1_L2_4_G1_MINI_ALU_OperationResult_2, 
         L1_1_L2_4_G1_MINI_ALU_OperationResult_1, 
         L1_1_L2_4_G1_MINI_ALU_OperationResult_0, 
         L1_1_L2_4_G1_MINI_ALU_BoothXORCheck, 
         L1_1_L2_4_G1_MINI_ALU_BoothOperand_16, 
         L1_1_L2_4_G1_MINI_ALU_BoothOperand_15, 
         L1_1_L2_4_G1_MINI_ALU_BoothOperand_14, 
         L1_1_L2_4_G1_MINI_ALU_BoothOperand_13, 
         L1_1_L2_4_G1_MINI_ALU_BoothOperand_12, 
         L1_1_L2_4_G1_MINI_ALU_BoothOperand_11, 
         L1_1_L2_4_G1_MINI_ALU_BoothOperand_10, 
         L1_1_L2_4_G1_MINI_ALU_BoothOperand_9, L1_1_L2_4_G1_MINI_ALU_BoothP_16, 
         L1_1_L2_4_G1_MINI_ALU_BoothP_15, L1_1_L2_4_G1_MINI_ALU_BoothP_14, 
         L1_1_L2_4_G1_MINI_ALU_BoothP_13, L1_1_L2_4_G1_MINI_ALU_BoothP_12, 
         L1_1_L2_4_G1_MINI_ALU_BoothP_11, L1_1_L2_4_G1_MINI_ALU_BoothP_10, 
         L1_1_L2_4_G1_MINI_ALU_BoothP_9, L1_1_L2_4_G1_MINI_ALU_BoothP_8, 
         L1_1_L2_4_G1_MINI_ALU_BoothP_7, L1_1_L2_4_G1_MINI_ALU_BoothP_6, 
         L1_1_L2_4_G1_MINI_ALU_BoothP_5, L1_1_L2_4_G1_MINI_ALU_BoothP_4, 
         L1_1_L2_4_G1_MINI_ALU_BoothP_3, L1_1_L2_4_G1_MINI_ALU_BoothP_2, 
         L1_1_L2_4_G1_MINI_ALU_BoothP_1, L1_1_L2_4_G1_MINI_ALU_BoothP_0, 
         L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_15, 
         L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_14, 
         L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_13, 
         L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_12, 
         L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_11, 
         L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_10, 
         L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_9, 
         L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_8, 
         L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_7, 
         L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_6, 
         L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_5, 
         L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_4, 
         L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_3, 
         L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_2, 
         L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_1, 
         L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_0, 
         L1_2_L2_0_G1_MINI_ALU_OperationResult_15, 
         L1_2_L2_0_G1_MINI_ALU_OperationResult_14, 
         L1_2_L2_0_G1_MINI_ALU_OperationResult_13, 
         L1_2_L2_0_G1_MINI_ALU_OperationResult_12, 
         L1_2_L2_0_G1_MINI_ALU_OperationResult_11, 
         L1_2_L2_0_G1_MINI_ALU_OperationResult_10, 
         L1_2_L2_0_G1_MINI_ALU_OperationResult_9, 
         L1_2_L2_0_G1_MINI_ALU_OperationResult_8, 
         L1_2_L2_0_G1_MINI_ALU_OperationResult_7, 
         L1_2_L2_0_G1_MINI_ALU_OperationResult_6, 
         L1_2_L2_0_G1_MINI_ALU_OperationResult_5, 
         L1_2_L2_0_G1_MINI_ALU_OperationResult_4, 
         L1_2_L2_0_G1_MINI_ALU_OperationResult_3, 
         L1_2_L2_0_G1_MINI_ALU_OperationResult_2, 
         L1_2_L2_0_G1_MINI_ALU_OperationResult_1, 
         L1_2_L2_0_G1_MINI_ALU_OperationResult_0, 
         L1_2_L2_0_G1_MINI_ALU_BoothXORCheck, 
         L1_2_L2_0_G1_MINI_ALU_BoothOperand_16, 
         L1_2_L2_0_G1_MINI_ALU_BoothOperand_15, 
         L1_2_L2_0_G1_MINI_ALU_BoothOperand_14, 
         L1_2_L2_0_G1_MINI_ALU_BoothOperand_13, 
         L1_2_L2_0_G1_MINI_ALU_BoothOperand_12, 
         L1_2_L2_0_G1_MINI_ALU_BoothOperand_11, 
         L1_2_L2_0_G1_MINI_ALU_BoothOperand_10, 
         L1_2_L2_0_G1_MINI_ALU_BoothOperand_9, L1_2_L2_0_G1_MINI_ALU_BoothP_16, 
         L1_2_L2_0_G1_MINI_ALU_BoothP_15, L1_2_L2_0_G1_MINI_ALU_BoothP_14, 
         L1_2_L2_0_G1_MINI_ALU_BoothP_13, L1_2_L2_0_G1_MINI_ALU_BoothP_12, 
         L1_2_L2_0_G1_MINI_ALU_BoothP_11, L1_2_L2_0_G1_MINI_ALU_BoothP_10, 
         L1_2_L2_0_G1_MINI_ALU_BoothP_9, L1_2_L2_0_G1_MINI_ALU_BoothP_8, 
         L1_2_L2_0_G1_MINI_ALU_BoothP_7, L1_2_L2_0_G1_MINI_ALU_BoothP_6, 
         L1_2_L2_0_G1_MINI_ALU_BoothP_5, L1_2_L2_0_G1_MINI_ALU_BoothP_4, 
         L1_2_L2_0_G1_MINI_ALU_BoothP_3, L1_2_L2_0_G1_MINI_ALU_BoothP_2, 
         L1_2_L2_0_G1_MINI_ALU_BoothP_1, L1_2_L2_0_G1_MINI_ALU_BoothP_0, 
         L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_15, 
         L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_14, 
         L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_13, 
         L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_12, 
         L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_11, 
         L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_10, 
         L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_9, 
         L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_8, 
         L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_7, 
         L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_6, 
         L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_5, 
         L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_4, 
         L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_3, 
         L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_2, 
         L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_1, 
         L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_0, 
         L1_2_L2_1_G1_MINI_ALU_OperationResult_15, 
         L1_2_L2_1_G1_MINI_ALU_OperationResult_14, 
         L1_2_L2_1_G1_MINI_ALU_OperationResult_13, 
         L1_2_L2_1_G1_MINI_ALU_OperationResult_12, 
         L1_2_L2_1_G1_MINI_ALU_OperationResult_11, 
         L1_2_L2_1_G1_MINI_ALU_OperationResult_10, 
         L1_2_L2_1_G1_MINI_ALU_OperationResult_9, 
         L1_2_L2_1_G1_MINI_ALU_OperationResult_8, 
         L1_2_L2_1_G1_MINI_ALU_OperationResult_7, 
         L1_2_L2_1_G1_MINI_ALU_OperationResult_6, 
         L1_2_L2_1_G1_MINI_ALU_OperationResult_5, 
         L1_2_L2_1_G1_MINI_ALU_OperationResult_4, 
         L1_2_L2_1_G1_MINI_ALU_OperationResult_3, 
         L1_2_L2_1_G1_MINI_ALU_OperationResult_2, 
         L1_2_L2_1_G1_MINI_ALU_OperationResult_1, 
         L1_2_L2_1_G1_MINI_ALU_OperationResult_0, 
         L1_2_L2_1_G1_MINI_ALU_BoothXORCheck, 
         L1_2_L2_1_G1_MINI_ALU_BoothOperand_16, 
         L1_2_L2_1_G1_MINI_ALU_BoothOperand_15, 
         L1_2_L2_1_G1_MINI_ALU_BoothOperand_14, 
         L1_2_L2_1_G1_MINI_ALU_BoothOperand_13, 
         L1_2_L2_1_G1_MINI_ALU_BoothOperand_12, 
         L1_2_L2_1_G1_MINI_ALU_BoothOperand_11, 
         L1_2_L2_1_G1_MINI_ALU_BoothOperand_10, 
         L1_2_L2_1_G1_MINI_ALU_BoothOperand_9, L1_2_L2_1_G1_MINI_ALU_BoothP_16, 
         L1_2_L2_1_G1_MINI_ALU_BoothP_15, L1_2_L2_1_G1_MINI_ALU_BoothP_14, 
         L1_2_L2_1_G1_MINI_ALU_BoothP_13, L1_2_L2_1_G1_MINI_ALU_BoothP_12, 
         L1_2_L2_1_G1_MINI_ALU_BoothP_11, L1_2_L2_1_G1_MINI_ALU_BoothP_10, 
         L1_2_L2_1_G1_MINI_ALU_BoothP_9, L1_2_L2_1_G1_MINI_ALU_BoothP_8, 
         L1_2_L2_1_G1_MINI_ALU_BoothP_7, L1_2_L2_1_G1_MINI_ALU_BoothP_6, 
         L1_2_L2_1_G1_MINI_ALU_BoothP_5, L1_2_L2_1_G1_MINI_ALU_BoothP_4, 
         L1_2_L2_1_G1_MINI_ALU_BoothP_3, L1_2_L2_1_G1_MINI_ALU_BoothP_2, 
         L1_2_L2_1_G1_MINI_ALU_BoothP_1, L1_2_L2_1_G1_MINI_ALU_BoothP_0, 
         L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_15, 
         L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_14, 
         L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_13, 
         L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_12, 
         L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_11, 
         L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_10, 
         L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_9, 
         L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_8, 
         L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_7, 
         L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_6, 
         L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_5, 
         L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_4, 
         L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_3, 
         L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_2, 
         L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_1, 
         L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_0, 
         L1_2_L2_2_G1_MINI_ALU_BoothXORCheck, 
         L1_2_L2_2_G1_MINI_ALU_BoothOperand_16, 
         L1_2_L2_2_G1_MINI_ALU_BoothOperand_15, 
         L1_2_L2_2_G1_MINI_ALU_BoothOperand_14, 
         L1_2_L2_2_G1_MINI_ALU_BoothOperand_13, 
         L1_2_L2_2_G1_MINI_ALU_BoothOperand_12, 
         L1_2_L2_2_G1_MINI_ALU_BoothOperand_11, 
         L1_2_L2_2_G1_MINI_ALU_BoothOperand_10, 
         L1_2_L2_2_G1_MINI_ALU_BoothOperand_9, L1_2_L2_2_G1_MINI_ALU_BoothP_16, 
         L1_2_L2_2_G1_MINI_ALU_BoothP_15, L1_2_L2_2_G1_MINI_ALU_BoothP_14, 
         L1_2_L2_2_G1_MINI_ALU_BoothP_13, L1_2_L2_2_G1_MINI_ALU_BoothP_12, 
         L1_2_L2_2_G1_MINI_ALU_BoothP_11, L1_2_L2_2_G1_MINI_ALU_BoothP_10, 
         L1_2_L2_2_G1_MINI_ALU_BoothP_9, L1_2_L2_2_G1_MINI_ALU_BoothP_8, 
         L1_2_L2_2_G1_MINI_ALU_BoothP_7, L1_2_L2_2_G1_MINI_ALU_BoothP_6, 
         L1_2_L2_2_G1_MINI_ALU_BoothP_5, L1_2_L2_2_G1_MINI_ALU_BoothP_4, 
         L1_2_L2_2_G1_MINI_ALU_BoothP_3, L1_2_L2_2_G1_MINI_ALU_BoothP_2, 
         L1_2_L2_2_G1_MINI_ALU_BoothP_1, 
         L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_15, 
         L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_14, 
         L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_13, 
         L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_12, 
         L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_11, 
         L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_10, 
         L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_9, 
         L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_8, 
         L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_7, 
         L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_6, 
         L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_5, 
         L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_4, 
         L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_3, 
         L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_2, 
         L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_1, 
         L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_0, 
         L1_2_L2_3_G2_MINI_ALU_BoothXORCheck, 
         L1_2_L2_3_G2_MINI_ALU_BoothOperand_16, 
         L1_2_L2_3_G2_MINI_ALU_BoothOperand_15, 
         L1_2_L2_3_G2_MINI_ALU_BoothOperand_14, 
         L1_2_L2_3_G2_MINI_ALU_BoothOperand_13, 
         L1_2_L2_3_G2_MINI_ALU_BoothOperand_12, 
         L1_2_L2_3_G2_MINI_ALU_BoothOperand_11, 
         L1_2_L2_3_G2_MINI_ALU_BoothOperand_10, 
         L1_2_L2_3_G2_MINI_ALU_BoothOperand_9, L1_2_L2_3_G2_MINI_ALU_BoothP_16, 
         L1_2_L2_3_G2_MINI_ALU_BoothP_15, L1_2_L2_3_G2_MINI_ALU_BoothP_14, 
         L1_2_L2_3_G2_MINI_ALU_BoothP_13, L1_2_L2_3_G2_MINI_ALU_BoothP_12, 
         L1_2_L2_3_G2_MINI_ALU_BoothP_11, L1_2_L2_3_G2_MINI_ALU_BoothP_10, 
         L1_2_L2_3_G2_MINI_ALU_BoothP_9, L1_2_L2_3_G2_MINI_ALU_BoothP_8, 
         L1_2_L2_3_G2_MINI_ALU_BoothP_7, L1_2_L2_3_G2_MINI_ALU_BoothP_6, 
         L1_2_L2_3_G2_MINI_ALU_BoothP_5, L1_2_L2_3_G2_MINI_ALU_BoothP_4, 
         L1_2_L2_3_G2_MINI_ALU_BoothP_3, L1_2_L2_3_G2_MINI_ALU_BoothP_2, 
         L1_2_L2_3_G2_MINI_ALU_BoothP_1, L1_2_L2_3_G2_MINI_ALU_BoothP_0, 
         L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_15, 
         L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_14, 
         L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_13, 
         L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_12, 
         L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_11, 
         L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_10, 
         L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_9, 
         L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_8, 
         L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_7, 
         L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_6, 
         L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_5, 
         L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_4, 
         L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_3, 
         L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_2, 
         L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_1, 
         L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_0, 
         L1_2_L2_4_G2_MINI_ALU_BoothXORCheck, 
         L1_2_L2_4_G2_MINI_ALU_BoothOperand_16, 
         L1_2_L2_4_G2_MINI_ALU_BoothOperand_15, 
         L1_2_L2_4_G2_MINI_ALU_BoothOperand_14, 
         L1_2_L2_4_G2_MINI_ALU_BoothOperand_13, 
         L1_2_L2_4_G2_MINI_ALU_BoothOperand_12, 
         L1_2_L2_4_G2_MINI_ALU_BoothOperand_11, 
         L1_2_L2_4_G2_MINI_ALU_BoothOperand_10, 
         L1_2_L2_4_G2_MINI_ALU_BoothOperand_9, L1_2_L2_4_G2_MINI_ALU_BoothP_16, 
         L1_2_L2_4_G2_MINI_ALU_BoothP_15, L1_2_L2_4_G2_MINI_ALU_BoothP_14, 
         L1_2_L2_4_G2_MINI_ALU_BoothP_13, L1_2_L2_4_G2_MINI_ALU_BoothP_12, 
         L1_2_L2_4_G2_MINI_ALU_BoothP_11, L1_2_L2_4_G2_MINI_ALU_BoothP_10, 
         L1_2_L2_4_G2_MINI_ALU_BoothP_9, L1_2_L2_4_G2_MINI_ALU_BoothP_8, 
         L1_2_L2_4_G2_MINI_ALU_BoothP_7, L1_2_L2_4_G2_MINI_ALU_BoothP_6, 
         L1_2_L2_4_G2_MINI_ALU_BoothP_5, L1_2_L2_4_G2_MINI_ALU_BoothP_4, 
         L1_2_L2_4_G2_MINI_ALU_BoothP_3, L1_2_L2_4_G2_MINI_ALU_BoothP_2, 
         L1_2_L2_4_G2_MINI_ALU_BoothP_1, L1_2_L2_4_G2_MINI_ALU_BoothP_0, 
         L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_15, 
         L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_14, 
         L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_13, 
         L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_12, 
         L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_11, 
         L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_10, 
         L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_9, 
         L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_8, 
         L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_7, 
         L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_6, 
         L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_5, 
         L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_4, 
         L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_3, 
         L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_2, 
         L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_1, 
         L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_0, 
         L1_3_L2_0_G2_MINI_ALU_BoothXORCheck, 
         L1_3_L2_0_G2_MINI_ALU_BoothOperand_16, 
         L1_3_L2_0_G2_MINI_ALU_BoothOperand_15, 
         L1_3_L2_0_G2_MINI_ALU_BoothOperand_14, 
         L1_3_L2_0_G2_MINI_ALU_BoothOperand_13, 
         L1_3_L2_0_G2_MINI_ALU_BoothOperand_12, 
         L1_3_L2_0_G2_MINI_ALU_BoothOperand_11, 
         L1_3_L2_0_G2_MINI_ALU_BoothOperand_10, 
         L1_3_L2_0_G2_MINI_ALU_BoothOperand_9, L1_3_L2_0_G2_MINI_ALU_BoothP_16, 
         L1_3_L2_0_G2_MINI_ALU_BoothP_15, L1_3_L2_0_G2_MINI_ALU_BoothP_14, 
         L1_3_L2_0_G2_MINI_ALU_BoothP_13, L1_3_L2_0_G2_MINI_ALU_BoothP_12, 
         L1_3_L2_0_G2_MINI_ALU_BoothP_11, L1_3_L2_0_G2_MINI_ALU_BoothP_10, 
         L1_3_L2_0_G2_MINI_ALU_BoothP_9, L1_3_L2_0_G2_MINI_ALU_BoothP_8, 
         L1_3_L2_0_G2_MINI_ALU_BoothP_7, L1_3_L2_0_G2_MINI_ALU_BoothP_6, 
         L1_3_L2_0_G2_MINI_ALU_BoothP_5, L1_3_L2_0_G2_MINI_ALU_BoothP_4, 
         L1_3_L2_0_G2_MINI_ALU_BoothP_3, L1_3_L2_0_G2_MINI_ALU_BoothP_2, 
         L1_3_L2_0_G2_MINI_ALU_BoothP_1, L1_3_L2_0_G2_MINI_ALU_BoothP_0, 
         L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_15, 
         L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_14, 
         L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_13, 
         L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_12, 
         L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_11, 
         L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_10, 
         L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_9, 
         L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_8, 
         L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_7, 
         L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_6, 
         L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_5, 
         L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_4, 
         L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_3, 
         L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_2, 
         L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_1, 
         L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_0, 
         L1_3_L2_1_G2_MINI_ALU_BoothXORCheck, 
         L1_3_L2_1_G2_MINI_ALU_BoothOperand_16, 
         L1_3_L2_1_G2_MINI_ALU_BoothOperand_15, 
         L1_3_L2_1_G2_MINI_ALU_BoothOperand_14, 
         L1_3_L2_1_G2_MINI_ALU_BoothOperand_13, 
         L1_3_L2_1_G2_MINI_ALU_BoothOperand_12, 
         L1_3_L2_1_G2_MINI_ALU_BoothOperand_11, 
         L1_3_L2_1_G2_MINI_ALU_BoothOperand_10, 
         L1_3_L2_1_G2_MINI_ALU_BoothOperand_9, L1_3_L2_1_G2_MINI_ALU_BoothP_16, 
         L1_3_L2_1_G2_MINI_ALU_BoothP_15, L1_3_L2_1_G2_MINI_ALU_BoothP_14, 
         L1_3_L2_1_G2_MINI_ALU_BoothP_13, L1_3_L2_1_G2_MINI_ALU_BoothP_12, 
         L1_3_L2_1_G2_MINI_ALU_BoothP_11, L1_3_L2_1_G2_MINI_ALU_BoothP_10, 
         L1_3_L2_1_G2_MINI_ALU_BoothP_9, L1_3_L2_1_G2_MINI_ALU_BoothP_8, 
         L1_3_L2_1_G2_MINI_ALU_BoothP_7, L1_3_L2_1_G2_MINI_ALU_BoothP_6, 
         L1_3_L2_1_G2_MINI_ALU_BoothP_5, L1_3_L2_1_G2_MINI_ALU_BoothP_4, 
         L1_3_L2_1_G2_MINI_ALU_BoothP_3, L1_3_L2_1_G2_MINI_ALU_BoothP_2, 
         L1_3_L2_1_G2_MINI_ALU_BoothP_1, L1_3_L2_1_G2_MINI_ALU_BoothP_0, 
         L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_15, 
         L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_14, 
         L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_13, 
         L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_12, 
         L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_11, 
         L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_10, 
         L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_9, 
         L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_8, 
         L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_7, 
         L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_6, 
         L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_5, 
         L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_4, 
         L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_3, 
         L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_2, 
         L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_1, 
         L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_0, 
         L1_3_L2_2_G2_MINI_ALU_BoothXORCheck, 
         L1_3_L2_2_G2_MINI_ALU_BoothOperand_16, 
         L1_3_L2_2_G2_MINI_ALU_BoothOperand_15, 
         L1_3_L2_2_G2_MINI_ALU_BoothOperand_14, 
         L1_3_L2_2_G2_MINI_ALU_BoothOperand_13, 
         L1_3_L2_2_G2_MINI_ALU_BoothOperand_12, 
         L1_3_L2_2_G2_MINI_ALU_BoothOperand_11, 
         L1_3_L2_2_G2_MINI_ALU_BoothOperand_10, 
         L1_3_L2_2_G2_MINI_ALU_BoothOperand_9, L1_3_L2_2_G2_MINI_ALU_BoothP_16, 
         L1_3_L2_2_G2_MINI_ALU_BoothP_15, L1_3_L2_2_G2_MINI_ALU_BoothP_14, 
         L1_3_L2_2_G2_MINI_ALU_BoothP_13, L1_3_L2_2_G2_MINI_ALU_BoothP_12, 
         L1_3_L2_2_G2_MINI_ALU_BoothP_11, L1_3_L2_2_G2_MINI_ALU_BoothP_10, 
         L1_3_L2_2_G2_MINI_ALU_BoothP_9, L1_3_L2_2_G2_MINI_ALU_BoothP_8, 
         L1_3_L2_2_G2_MINI_ALU_BoothP_7, L1_3_L2_2_G2_MINI_ALU_BoothP_6, 
         L1_3_L2_2_G2_MINI_ALU_BoothP_5, L1_3_L2_2_G2_MINI_ALU_BoothP_4, 
         L1_3_L2_2_G2_MINI_ALU_BoothP_3, L1_3_L2_2_G2_MINI_ALU_BoothP_2, 
         L1_3_L2_2_G2_MINI_ALU_BoothP_1, L1_3_L2_2_G2_MINI_ALU_BoothP_0, 
         L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_15, 
         L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_14, 
         L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_13, 
         L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_12, 
         L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_11, 
         L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_10, 
         L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_9, 
         L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_8, 
         L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_7, 
         L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_6, 
         L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_5, 
         L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_4, 
         L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_3, 
         L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_2, 
         L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_1, 
         L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_0, 
         L1_3_L2_3_G2_MINI_ALU_BoothXORCheck, 
         L1_3_L2_3_G2_MINI_ALU_BoothOperand_16, 
         L1_3_L2_3_G2_MINI_ALU_BoothOperand_15, 
         L1_3_L2_3_G2_MINI_ALU_BoothOperand_14, 
         L1_3_L2_3_G2_MINI_ALU_BoothOperand_13, 
         L1_3_L2_3_G2_MINI_ALU_BoothOperand_12, 
         L1_3_L2_3_G2_MINI_ALU_BoothOperand_11, 
         L1_3_L2_3_G2_MINI_ALU_BoothOperand_10, 
         L1_3_L2_3_G2_MINI_ALU_BoothOperand_9, L1_3_L2_3_G2_MINI_ALU_BoothP_16, 
         L1_3_L2_3_G2_MINI_ALU_BoothP_15, L1_3_L2_3_G2_MINI_ALU_BoothP_14, 
         L1_3_L2_3_G2_MINI_ALU_BoothP_13, L1_3_L2_3_G2_MINI_ALU_BoothP_12, 
         L1_3_L2_3_G2_MINI_ALU_BoothP_11, L1_3_L2_3_G2_MINI_ALU_BoothP_10, 
         L1_3_L2_3_G2_MINI_ALU_BoothP_9, L1_3_L2_3_G2_MINI_ALU_BoothP_8, 
         L1_3_L2_3_G2_MINI_ALU_BoothP_7, L1_3_L2_3_G2_MINI_ALU_BoothP_6, 
         L1_3_L2_3_G2_MINI_ALU_BoothP_5, L1_3_L2_3_G2_MINI_ALU_BoothP_4, 
         L1_3_L2_3_G2_MINI_ALU_BoothP_3, L1_3_L2_3_G2_MINI_ALU_BoothP_2, 
         L1_3_L2_3_G2_MINI_ALU_BoothP_1, L1_3_L2_3_G2_MINI_ALU_BoothP_0, 
         L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_15, 
         L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_14, 
         L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_13, 
         L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_12, 
         L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_11, 
         L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_10, 
         L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_9, 
         L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_8, 
         L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_7, 
         L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_6, 
         L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_5, 
         L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_4, 
         L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_3, 
         L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_2, 
         L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_1, 
         L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_0, 
         L1_3_L2_4_G3_MINI_ALU_BoothXORCheck, 
         L1_3_L2_4_G3_MINI_ALU_BoothOperand_16, 
         L1_3_L2_4_G3_MINI_ALU_BoothOperand_15, 
         L1_3_L2_4_G3_MINI_ALU_BoothOperand_14, 
         L1_3_L2_4_G3_MINI_ALU_BoothOperand_13, 
         L1_3_L2_4_G3_MINI_ALU_BoothOperand_12, 
         L1_3_L2_4_G3_MINI_ALU_BoothOperand_11, 
         L1_3_L2_4_G3_MINI_ALU_BoothOperand_10, 
         L1_3_L2_4_G3_MINI_ALU_BoothOperand_9, L1_3_L2_4_G3_MINI_ALU_BoothP_16, 
         L1_3_L2_4_G3_MINI_ALU_BoothP_15, L1_3_L2_4_G3_MINI_ALU_BoothP_14, 
         L1_3_L2_4_G3_MINI_ALU_BoothP_13, L1_3_L2_4_G3_MINI_ALU_BoothP_12, 
         L1_3_L2_4_G3_MINI_ALU_BoothP_11, L1_3_L2_4_G3_MINI_ALU_BoothP_10, 
         L1_3_L2_4_G3_MINI_ALU_BoothP_9, L1_3_L2_4_G3_MINI_ALU_BoothP_8, 
         L1_3_L2_4_G3_MINI_ALU_BoothP_7, L1_3_L2_4_G3_MINI_ALU_BoothP_6, 
         L1_3_L2_4_G3_MINI_ALU_BoothP_5, L1_3_L2_4_G3_MINI_ALU_BoothP_4, 
         L1_3_L2_4_G3_MINI_ALU_BoothP_3, L1_3_L2_4_G3_MINI_ALU_BoothP_2, 
         L1_3_L2_4_G3_MINI_ALU_BoothP_1, L1_3_L2_4_G3_MINI_ALU_BoothP_0, 
         L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_15, 
         L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_14, 
         L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_13, 
         L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_12, 
         L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_11, 
         L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_10, 
         L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_9, 
         L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_8, 
         L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_7, 
         L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_6, 
         L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_5, 
         L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_4, 
         L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_3, 
         L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_2, 
         L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_1, 
         L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_0, 
         L1_4_L2_0_G3_MINI_ALU_BoothXORCheck, 
         L1_4_L2_0_G3_MINI_ALU_BoothOperand_16, 
         L1_4_L2_0_G3_MINI_ALU_BoothOperand_15, 
         L1_4_L2_0_G3_MINI_ALU_BoothOperand_14, 
         L1_4_L2_0_G3_MINI_ALU_BoothOperand_13, 
         L1_4_L2_0_G3_MINI_ALU_BoothOperand_12, 
         L1_4_L2_0_G3_MINI_ALU_BoothOperand_11, 
         L1_4_L2_0_G3_MINI_ALU_BoothOperand_10, 
         L1_4_L2_0_G3_MINI_ALU_BoothOperand_9, L1_4_L2_0_G3_MINI_ALU_BoothP_16, 
         L1_4_L2_0_G3_MINI_ALU_BoothP_15, L1_4_L2_0_G3_MINI_ALU_BoothP_14, 
         L1_4_L2_0_G3_MINI_ALU_BoothP_13, L1_4_L2_0_G3_MINI_ALU_BoothP_12, 
         L1_4_L2_0_G3_MINI_ALU_BoothP_11, L1_4_L2_0_G3_MINI_ALU_BoothP_10, 
         L1_4_L2_0_G3_MINI_ALU_BoothP_9, L1_4_L2_0_G3_MINI_ALU_BoothP_8, 
         L1_4_L2_0_G3_MINI_ALU_BoothP_7, L1_4_L2_0_G3_MINI_ALU_BoothP_6, 
         L1_4_L2_0_G3_MINI_ALU_BoothP_5, L1_4_L2_0_G3_MINI_ALU_BoothP_4, 
         L1_4_L2_0_G3_MINI_ALU_BoothP_3, L1_4_L2_0_G3_MINI_ALU_BoothP_2, 
         L1_4_L2_0_G3_MINI_ALU_BoothP_1, L1_4_L2_0_G3_MINI_ALU_BoothP_0, 
         L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_15, 
         L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_14, 
         L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_13, 
         L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_12, 
         L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_11, 
         L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_10, 
         L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_9, 
         L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_8, 
         L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_7, 
         L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_6, 
         L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_5, 
         L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_4, 
         L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_3, 
         L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_2, 
         L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_1, 
         L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_0, 
         L1_4_L2_1_G3_MINI_ALU_BoothXORCheck, 
         L1_4_L2_1_G3_MINI_ALU_BoothOperand_16, 
         L1_4_L2_1_G3_MINI_ALU_BoothOperand_15, 
         L1_4_L2_1_G3_MINI_ALU_BoothOperand_14, 
         L1_4_L2_1_G3_MINI_ALU_BoothOperand_13, 
         L1_4_L2_1_G3_MINI_ALU_BoothOperand_12, 
         L1_4_L2_1_G3_MINI_ALU_BoothOperand_11, 
         L1_4_L2_1_G3_MINI_ALU_BoothOperand_10, 
         L1_4_L2_1_G3_MINI_ALU_BoothOperand_9, L1_4_L2_1_G3_MINI_ALU_BoothP_16, 
         L1_4_L2_1_G3_MINI_ALU_BoothP_15, L1_4_L2_1_G3_MINI_ALU_BoothP_14, 
         L1_4_L2_1_G3_MINI_ALU_BoothP_13, L1_4_L2_1_G3_MINI_ALU_BoothP_12, 
         L1_4_L2_1_G3_MINI_ALU_BoothP_11, L1_4_L2_1_G3_MINI_ALU_BoothP_10, 
         L1_4_L2_1_G3_MINI_ALU_BoothP_9, L1_4_L2_1_G3_MINI_ALU_BoothP_8, 
         L1_4_L2_1_G3_MINI_ALU_BoothP_7, L1_4_L2_1_G3_MINI_ALU_BoothP_6, 
         L1_4_L2_1_G3_MINI_ALU_BoothP_5, L1_4_L2_1_G3_MINI_ALU_BoothP_4, 
         L1_4_L2_1_G3_MINI_ALU_BoothP_3, L1_4_L2_1_G3_MINI_ALU_BoothP_2, 
         L1_4_L2_1_G3_MINI_ALU_BoothP_1, L1_4_L2_1_G3_MINI_ALU_BoothP_0, 
         L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_15, 
         L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_14, 
         L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_13, 
         L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_12, 
         L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_11, 
         L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_10, 
         L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_9, 
         L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_8, 
         L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_7, 
         L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_6, 
         L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_5, 
         L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_4, 
         L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_3, 
         L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_2, 
         L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_1, 
         L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_0, 
         L1_4_L2_2_G4_MINI_ALU_BoothXORCheck, 
         L1_4_L2_2_G4_MINI_ALU_BoothOperand_16, 
         L1_4_L2_2_G4_MINI_ALU_BoothOperand_15, 
         L1_4_L2_2_G4_MINI_ALU_BoothOperand_14, 
         L1_4_L2_2_G4_MINI_ALU_BoothOperand_13, 
         L1_4_L2_2_G4_MINI_ALU_BoothOperand_12, 
         L1_4_L2_2_G4_MINI_ALU_BoothOperand_11, 
         L1_4_L2_2_G4_MINI_ALU_BoothOperand_10, 
         L1_4_L2_2_G4_MINI_ALU_BoothOperand_9, L1_4_L2_2_G4_MINI_ALU_BoothP_16, 
         L1_4_L2_2_G4_MINI_ALU_BoothP_15, L1_4_L2_2_G4_MINI_ALU_BoothP_14, 
         L1_4_L2_2_G4_MINI_ALU_BoothP_13, L1_4_L2_2_G4_MINI_ALU_BoothP_12, 
         L1_4_L2_2_G4_MINI_ALU_BoothP_11, L1_4_L2_2_G4_MINI_ALU_BoothP_10, 
         L1_4_L2_2_G4_MINI_ALU_BoothP_9, L1_4_L2_2_G4_MINI_ALU_BoothP_8, 
         L1_4_L2_2_G4_MINI_ALU_BoothP_7, L1_4_L2_2_G4_MINI_ALU_BoothP_6, 
         L1_4_L2_2_G4_MINI_ALU_BoothP_5, L1_4_L2_2_G4_MINI_ALU_BoothP_4, 
         L1_4_L2_2_G4_MINI_ALU_BoothP_3, L1_4_L2_2_G4_MINI_ALU_BoothP_2, 
         L1_4_L2_2_G4_MINI_ALU_BoothP_1, L1_4_L2_2_G4_MINI_ALU_BoothP_0, 
         L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_15, 
         L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_14, 
         L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_13, 
         L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_12, 
         L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_11, 
         L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_10, 
         L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_9, 
         L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_8, 
         L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_7, 
         L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_6, 
         L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_5, 
         L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_4, 
         L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_3, 
         L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_2, 
         L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_1, 
         L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_0, 
         L1_4_L2_3_G5_MINI_ALU_BoothXORCheck, 
         L1_4_L2_3_G5_MINI_ALU_BoothOperand_16, 
         L1_4_L2_3_G5_MINI_ALU_BoothOperand_15, 
         L1_4_L2_3_G5_MINI_ALU_BoothOperand_14, 
         L1_4_L2_3_G5_MINI_ALU_BoothOperand_13, 
         L1_4_L2_3_G5_MINI_ALU_BoothOperand_12, 
         L1_4_L2_3_G5_MINI_ALU_BoothOperand_11, 
         L1_4_L2_3_G5_MINI_ALU_BoothOperand_10, 
         L1_4_L2_3_G5_MINI_ALU_BoothOperand_9, L1_4_L2_3_G5_MINI_ALU_BoothP_16, 
         L1_4_L2_3_G5_MINI_ALU_BoothP_15, L1_4_L2_3_G5_MINI_ALU_BoothP_14, 
         L1_4_L2_3_G5_MINI_ALU_BoothP_13, L1_4_L2_3_G5_MINI_ALU_BoothP_12, 
         L1_4_L2_3_G5_MINI_ALU_BoothP_11, L1_4_L2_3_G5_MINI_ALU_BoothP_10, 
         L1_4_L2_3_G5_MINI_ALU_BoothP_9, L1_4_L2_3_G5_MINI_ALU_BoothP_8, 
         L1_4_L2_3_G5_MINI_ALU_BoothP_7, L1_4_L2_3_G5_MINI_ALU_BoothP_6, 
         L1_4_L2_3_G5_MINI_ALU_BoothP_5, L1_4_L2_3_G5_MINI_ALU_BoothP_4, 
         L1_4_L2_3_G5_MINI_ALU_BoothP_3, L1_4_L2_3_G5_MINI_ALU_BoothP_2, 
         L1_4_L2_3_G5_MINI_ALU_BoothP_1, L1_4_L2_3_G5_MINI_ALU_BoothP_0, 
         L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_15, 
         L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_14, 
         L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_13, 
         L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_12, 
         L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_11, 
         L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_10, 
         L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_9, 
         L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_8, 
         L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_7, 
         L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_6, 
         L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_5, 
         L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_4, 
         L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_3, 
         L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_2, 
         L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_1, 
         L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_0, 
         L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_7, 
         L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_6, 
         L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_5, 
         L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_4, 
         L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_3, 
         L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_2, 
         L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_1, 
         L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_0, 
         L1_4_L2_4_G5_MINI_ALU_OperationResult_15, 
         L1_4_L2_4_G5_MINI_ALU_OperationResult_14, 
         L1_4_L2_4_G5_MINI_ALU_OperationResult_13, 
         L1_4_L2_4_G5_MINI_ALU_OperationResult_12, 
         L1_4_L2_4_G5_MINI_ALU_OperationResult_11, 
         L1_4_L2_4_G5_MINI_ALU_OperationResult_10, 
         L1_4_L2_4_G5_MINI_ALU_OperationResult_9, 
         L1_4_L2_4_G5_MINI_ALU_OperationResult_8, 
         L1_4_L2_4_G5_MINI_ALU_OperationResult_7, 
         L1_4_L2_4_G5_MINI_ALU_OperationResult_6, 
         L1_4_L2_4_G5_MINI_ALU_OperationResult_5, 
         L1_4_L2_4_G5_MINI_ALU_OperationResult_4, 
         L1_4_L2_4_G5_MINI_ALU_OperationResult_3, 
         L1_4_L2_4_G5_MINI_ALU_OperationResult_2, 
         L1_4_L2_4_G5_MINI_ALU_OperationResult_1, 
         L1_4_L2_4_G5_MINI_ALU_OperationResult_0, 
         L1_4_L2_4_G5_MINI_ALU_BoothXORCheck, 
         L1_4_L2_4_G5_MINI_ALU_BoothOperand_16, 
         L1_4_L2_4_G5_MINI_ALU_BoothOperand_15, 
         L1_4_L2_4_G5_MINI_ALU_BoothOperand_14, 
         L1_4_L2_4_G5_MINI_ALU_BoothOperand_13, 
         L1_4_L2_4_G5_MINI_ALU_BoothOperand_12, 
         L1_4_L2_4_G5_MINI_ALU_BoothOperand_11, 
         L1_4_L2_4_G5_MINI_ALU_BoothOperand_10, 
         L1_4_L2_4_G5_MINI_ALU_BoothOperand_9, L1_4_L2_4_G5_MINI_ALU_BoothP_16, 
         L1_4_L2_4_G5_MINI_ALU_BoothP_15, L1_4_L2_4_G5_MINI_ALU_BoothP_14, 
         L1_4_L2_4_G5_MINI_ALU_BoothP_13, L1_4_L2_4_G5_MINI_ALU_BoothP_12, 
         L1_4_L2_4_G5_MINI_ALU_BoothP_11, L1_4_L2_4_G5_MINI_ALU_BoothP_10, 
         L1_4_L2_4_G5_MINI_ALU_BoothP_9, L1_4_L2_4_G5_MINI_ALU_BoothP_8, 
         L1_4_L2_4_G5_MINI_ALU_BoothP_7, L1_4_L2_4_G5_MINI_ALU_BoothP_6, 
         L1_4_L2_4_G5_MINI_ALU_BoothP_5, L1_4_L2_4_G5_MINI_ALU_BoothP_4, 
         L1_4_L2_4_G5_MINI_ALU_BoothP_3, L1_4_L2_4_G5_MINI_ALU_BoothP_2, 
         L1_4_L2_4_G5_MINI_ALU_BoothP_1, L1_4_L2_4_G5_MINI_ALU_BoothP_0, 
         L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_15, 
         L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_14, 
         L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_13, 
         L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_12, 
         L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_11, 
         L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_10, 
         L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_9, 
         L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_8, 
         L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_7, 
         L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_6, 
         L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_5, 
         L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_4, 
         L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_3, 
         L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_2, 
         L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_1, 
         L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_0, L1FirstOperands_12__16, nx22, 
         CounterOut_0, NOT__13497, nx1032, NOT_CounterOut_0, nx1036, 
         CounterOut_3, CounterOut_2, CounterOut_1, nx1046, nx1058, nx1066, 
         nx2856, nx2868, nx2872, nx2876, nx3233, nx3236, nx3238, nx3242, nx3244, 
         nx3247, nx3249, nx3273, nx3275, nx3277, nx3279, nx3281, nx3283, nx3285, 
         nx3287, nx3289, nx3303, nx5, nx1, nx3304, nx3305, nx3306, nx3308;
    wire [901:0] \$dummy ;




    booth_adder_17 L1_0_L2_0_G1_MINI_ALU_BOOTH_ADDER (.AdderFirstOperand ({
                   L1FirstOperands_12__16,L1FirstOperands_0__15,
                   L1FirstOperands_0__14,L1FirstOperands_0__13,
                   L1FirstOperands_0__12,L1FirstOperands_0__11,
                   L1FirstOperands_0__10,L1FirstOperands_0__9,
                   L1FirstOperands_0__8,L1FirstOperands_0__7,
                   L1FirstOperands_0__6,L1FirstOperands_0__5,
                   L1FirstOperands_0__4,L1FirstOperands_0__3,
                   L1FirstOperands_0__2,L1FirstOperands_0__1,
                   L1FirstOperands_0__0}), .AdderSecondOperand ({
                   L1FirstOperands_12__16,
                   L1_0_L2_0_G1_MINI_ALU_OperationResult_15,
                   L1_0_L2_0_G1_MINI_ALU_OperationResult_14,
                   L1_0_L2_0_G1_MINI_ALU_OperationResult_13,
                   L1_0_L2_0_G1_MINI_ALU_OperationResult_12,
                   L1_0_L2_0_G1_MINI_ALU_OperationResult_11,
                   L1_0_L2_0_G1_MINI_ALU_OperationResult_10,
                   L1_0_L2_0_G1_MINI_ALU_OperationResult_9,
                   L1_0_L2_0_G1_MINI_ALU_OperationResult_8,
                   L1_0_L2_0_G1_MINI_ALU_OperationResult_7,
                   L1_0_L2_0_G1_MINI_ALU_OperationResult_6,
                   L1_0_L2_0_G1_MINI_ALU_OperationResult_5,
                   L1_0_L2_0_G1_MINI_ALU_OperationResult_4,
                   L1_0_L2_0_G1_MINI_ALU_OperationResult_3,
                   L1_0_L2_0_G1_MINI_ALU_OperationResult_2,
                   L1_0_L2_0_G1_MINI_ALU_OperationResult_1,
                   L1_0_L2_0_G1_MINI_ALU_OperationResult_0}), .BoothOperand ({
                   L1_0_L2_0_G1_MINI_ALU_BoothOperand_16,
                   L1_0_L2_0_G1_MINI_ALU_BoothOperand_15,
                   L1_0_L2_0_G1_MINI_ALU_BoothOperand_14,
                   L1_0_L2_0_G1_MINI_ALU_BoothOperand_13,
                   L1_0_L2_0_G1_MINI_ALU_BoothOperand_12,
                   L1_0_L2_0_G1_MINI_ALU_BoothOperand_11,
                   L1_0_L2_0_G1_MINI_ALU_BoothOperand_10,
                   L1_0_L2_0_G1_MINI_ALU_BoothOperand_9,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16}), .BoothP ({
                   L1_0_L2_0_G1_MINI_ALU_BoothP_16,
                   L1_0_L2_0_G1_MINI_ALU_BoothP_15,
                   L1_0_L2_0_G1_MINI_ALU_BoothP_14,
                   L1_0_L2_0_G1_MINI_ALU_BoothP_13,
                   L1_0_L2_0_G1_MINI_ALU_BoothP_12,
                   L1_0_L2_0_G1_MINI_ALU_BoothP_11,
                   L1_0_L2_0_G1_MINI_ALU_BoothP_10,
                   L1_0_L2_0_G1_MINI_ALU_BoothP_9,L1_0_L2_0_G1_MINI_ALU_BoothP_8
                   ,L1_0_L2_0_G1_MINI_ALU_BoothP_7,
                   L1_0_L2_0_G1_MINI_ALU_BoothP_6,L1_0_L2_0_G1_MINI_ALU_BoothP_5
                   ,L1_0_L2_0_G1_MINI_ALU_BoothP_4,
                   L1_0_L2_0_G1_MINI_ALU_BoothP_3,L1_0_L2_0_G1_MINI_ALU_BoothP_2
                   ,L1_0_L2_0_G1_MINI_ALU_BoothP_1,
                   L1_0_L2_0_G1_MINI_ALU_BoothP_0}), .SelOperand (nx3285), .Operation (
                   L1_0_L2_0_G1_MINI_ALU_BoothXORCheck), .AdderResult ({
                   L1ResultsLarge_0__16,L1ResultsLarge_0__15,
                   L1ResultsLarge_0__14,L1ResultsLarge_0__13,
                   L1ResultsLarge_0__12,L1ResultsLarge_0__11,
                   L1ResultsLarge_0__10,L1ResultsLarge_0__9,L1ResultsLarge_0__8,
                   L1ResultsLarge_0__7,L1ResultsLarge_0__6,L1ResultsLarge_0__5,
                   L1ResultsLarge_0__4,L1ResultsLarge_0__3,L1ResultsLarge_0__2,
                   L1ResultsLarge_0__1,L1ResultsLarge_0__0}), .AdderBoothResult (
                   {\$dummy [0],L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_15,
                   L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_14,
                   L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_13,
                   L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_12,
                   L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_11,
                   L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_10,
                   L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_9,
                   L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_8,
                   L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_7,
                   L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_6,
                   L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_5,
                   L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_4,
                   L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_3,
                   L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_2,
                   L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_1,
                   L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_0})) ;
    booth_unit_17 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT (.CLK (CLK), .RST (RST), .Start (
                  Start), .Instr (Instr), .LoopingAndResultNotReady (nx3275), .Filter (
                  {FilterDin_0__0__7,FilterDin_0__0__6,FilterDin_0__0__5,
                  FilterDin_0__0__4,FilterDin_0__0__3,FilterDin_0__0__2,
                  FilterDin_0__0__1,FilterDin_0__0__0}), .Window ({
                  WindowDin_0__0__7,WindowDin_0__0__6,WindowDin_0__0__5,
                  WindowDin_0__0__4,WindowDin_0__0__3,WindowDin_0__0__2,
                  WindowDin_0__0__1,WindowDin_0__0__0}), .AdderBoothResult ({
                  L1FirstOperands_12__16,
                  L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_15,
                  L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_14,
                  L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_13,
                  L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_12,
                  L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_11,
                  L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_10,
                  L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_9,
                  L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_8,
                  L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_7,
                  L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_6,
                  L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_5,
                  L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_4,
                  L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_3,
                  L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_2,
                  L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_1,
                  L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_0}), .BoothXORCheck (
                  L1_0_L2_0_G1_MINI_ALU_BoothXORCheck), .BoothResult ({
                  \$dummy [1],\$dummy [2],\$dummy [3],\$dummy [4],\$dummy [5],
                  \$dummy [6],\$dummy [7],\$dummy [8]}), .BoothAddingOperand ({
                  L1_0_L2_0_G1_MINI_ALU_BoothOperand_16,
                  L1_0_L2_0_G1_MINI_ALU_BoothOperand_15,
                  L1_0_L2_0_G1_MINI_ALU_BoothOperand_14,
                  L1_0_L2_0_G1_MINI_ALU_BoothOperand_13,
                  L1_0_L2_0_G1_MINI_ALU_BoothOperand_12,
                  L1_0_L2_0_G1_MINI_ALU_BoothOperand_11,
                  L1_0_L2_0_G1_MINI_ALU_BoothOperand_10,
                  L1_0_L2_0_G1_MINI_ALU_BoothOperand_9,\$dummy [9],\$dummy [10],
                  \$dummy [11],\$dummy [12],\$dummy [13],\$dummy [14],
                  \$dummy [15],\$dummy [16],\$dummy [17]}), .BoothP ({
                  L1_0_L2_0_G1_MINI_ALU_BoothP_16,
                  L1_0_L2_0_G1_MINI_ALU_BoothP_15,
                  L1_0_L2_0_G1_MINI_ALU_BoothP_14,
                  L1_0_L2_0_G1_MINI_ALU_BoothP_13,
                  L1_0_L2_0_G1_MINI_ALU_BoothP_12,
                  L1_0_L2_0_G1_MINI_ALU_BoothP_11,
                  L1_0_L2_0_G1_MINI_ALU_BoothP_10,L1_0_L2_0_G1_MINI_ALU_BoothP_9
                  ,L1_0_L2_0_G1_MINI_ALU_BoothP_8,L1_0_L2_0_G1_MINI_ALU_BoothP_7
                  ,L1_0_L2_0_G1_MINI_ALU_BoothP_6,L1_0_L2_0_G1_MINI_ALU_BoothP_5
                  ,L1_0_L2_0_G1_MINI_ALU_BoothP_4,L1_0_L2_0_G1_MINI_ALU_BoothP_3
                  ,L1_0_L2_0_G1_MINI_ALU_BoothP_2,L1_0_L2_0_G1_MINI_ALU_BoothP_1
                  ,L1_0_L2_0_G1_MINI_ALU_BoothP_0}), .LargeWindowShifted ({
                  \$dummy [18],\$dummy [19],\$dummy [20],\$dummy [21],
                  \$dummy [22],\$dummy [23],\$dummy [24],\$dummy [25],
                  \$dummy [26],\$dummy [27],\$dummy [28],\$dummy [29],
                  \$dummy [30],\$dummy [31],\$dummy [32],\$dummy [33],
                  \$dummy [34]})) ;
    booth_adder_17 L1_0_L2_1_G1_MINI_ALU_BOOTH_ADDER (.AdderFirstOperand ({
                   L1FirstOperands_12__16,L1FirstOperands_0__15,
                   L1FirstOperands_0__14,L1FirstOperands_0__13,
                   L1FirstOperands_0__12,L1FirstOperands_0__11,
                   L1FirstOperands_0__10,L1FirstOperands_0__9,
                   L1FirstOperands_0__8,L1FirstOperands_0__7,
                   L1FirstOperands_0__6,L1FirstOperands_0__5,
                   L1FirstOperands_0__4,L1FirstOperands_0__3,
                   L1FirstOperands_0__2,L1FirstOperands_0__1,
                   L1FirstOperands_0__0}), .AdderSecondOperand ({
                   L1FirstOperands_12__16,
                   L1_0_L2_1_G1_MINI_ALU_OperationResult_15,
                   L1_0_L2_1_G1_MINI_ALU_OperationResult_14,
                   L1_0_L2_1_G1_MINI_ALU_OperationResult_13,
                   L1_0_L2_1_G1_MINI_ALU_OperationResult_12,
                   L1_0_L2_1_G1_MINI_ALU_OperationResult_11,
                   L1_0_L2_1_G1_MINI_ALU_OperationResult_10,
                   L1_0_L2_1_G1_MINI_ALU_OperationResult_9,
                   L1_0_L2_1_G1_MINI_ALU_OperationResult_8,
                   L1_0_L2_1_G1_MINI_ALU_OperationResult_7,
                   L1_0_L2_1_G1_MINI_ALU_OperationResult_6,
                   L1_0_L2_1_G1_MINI_ALU_OperationResult_5,
                   L1_0_L2_1_G1_MINI_ALU_OperationResult_4,
                   L1_0_L2_1_G1_MINI_ALU_OperationResult_3,
                   L1_0_L2_1_G1_MINI_ALU_OperationResult_2,
                   L1_0_L2_1_G1_MINI_ALU_OperationResult_1,
                   L1_0_L2_1_G1_MINI_ALU_OperationResult_0}), .BoothOperand ({
                   L1_0_L2_1_G1_MINI_ALU_BoothOperand_16,
                   L1_0_L2_1_G1_MINI_ALU_BoothOperand_15,
                   L1_0_L2_1_G1_MINI_ALU_BoothOperand_14,
                   L1_0_L2_1_G1_MINI_ALU_BoothOperand_13,
                   L1_0_L2_1_G1_MINI_ALU_BoothOperand_12,
                   L1_0_L2_1_G1_MINI_ALU_BoothOperand_11,
                   L1_0_L2_1_G1_MINI_ALU_BoothOperand_10,
                   L1_0_L2_1_G1_MINI_ALU_BoothOperand_9,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16}), .BoothP ({
                   L1_0_L2_1_G1_MINI_ALU_BoothP_16,
                   L1_0_L2_1_G1_MINI_ALU_BoothP_15,
                   L1_0_L2_1_G1_MINI_ALU_BoothP_14,
                   L1_0_L2_1_G1_MINI_ALU_BoothP_13,
                   L1_0_L2_1_G1_MINI_ALU_BoothP_12,
                   L1_0_L2_1_G1_MINI_ALU_BoothP_11,
                   L1_0_L2_1_G1_MINI_ALU_BoothP_10,
                   L1_0_L2_1_G1_MINI_ALU_BoothP_9,L1_0_L2_1_G1_MINI_ALU_BoothP_8
                   ,L1_0_L2_1_G1_MINI_ALU_BoothP_7,
                   L1_0_L2_1_G1_MINI_ALU_BoothP_6,L1_0_L2_1_G1_MINI_ALU_BoothP_5
                   ,L1_0_L2_1_G1_MINI_ALU_BoothP_4,
                   L1_0_L2_1_G1_MINI_ALU_BoothP_3,L1_0_L2_1_G1_MINI_ALU_BoothP_2
                   ,L1_0_L2_1_G1_MINI_ALU_BoothP_1,
                   L1_0_L2_1_G1_MINI_ALU_BoothP_0}), .SelOperand (nx3285), .Operation (
                   L1_0_L2_1_G1_MINI_ALU_BoothXORCheck), .AdderResult ({
                   L1ResultsLarge_1__16,L1ResultsLarge_1__15,
                   L1ResultsLarge_1__14,L1ResultsLarge_1__13,
                   L1ResultsLarge_1__12,L1ResultsLarge_1__11,
                   L1ResultsLarge_1__10,L1ResultsLarge_1__9,L1ResultsLarge_1__8,
                   L1ResultsLarge_1__7,L1ResultsLarge_1__6,L1ResultsLarge_1__5,
                   L1ResultsLarge_1__4,L1ResultsLarge_1__3,L1ResultsLarge_1__2,
                   L1ResultsLarge_1__1,L1ResultsLarge_1__0}), .AdderBoothResult (
                   {\$dummy [35],L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_15,
                   L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_14,
                   L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_13,
                   L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_12,
                   L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_11,
                   L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_10,
                   L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_9,
                   L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_8,
                   L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_7,
                   L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_6,
                   L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_5,
                   L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_4,
                   L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_3,
                   L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_2,
                   L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_1,
                   L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_0})) ;
    booth_unit_17 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT (.CLK (CLK), .RST (RST), .Start (
                  Start), .Instr (Instr), .LoopingAndResultNotReady (nx3275), .Filter (
                  {FilterDin_0__1__7,FilterDin_0__1__6,FilterDin_0__1__5,
                  FilterDin_0__1__4,FilterDin_0__1__3,FilterDin_0__1__2,
                  FilterDin_0__1__1,FilterDin_0__1__0}), .Window ({
                  WindowDin_0__1__7,WindowDin_0__1__6,WindowDin_0__1__5,
                  WindowDin_0__1__4,WindowDin_0__1__3,WindowDin_0__1__2,
                  WindowDin_0__1__1,WindowDin_0__1__0}), .AdderBoothResult ({
                  L1FirstOperands_12__16,
                  L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_15,
                  L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_14,
                  L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_13,
                  L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_12,
                  L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_11,
                  L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_10,
                  L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_9,
                  L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_8,
                  L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_7,
                  L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_6,
                  L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_5,
                  L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_4,
                  L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_3,
                  L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_2,
                  L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_1,
                  L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_0}), .BoothXORCheck (
                  L1_0_L2_1_G1_MINI_ALU_BoothXORCheck), .BoothResult ({
                  \$dummy [36],\$dummy [37],\$dummy [38],\$dummy [39],
                  \$dummy [40],\$dummy [41],\$dummy [42],\$dummy [43]}), .BoothAddingOperand (
                  {L1_0_L2_1_G1_MINI_ALU_BoothOperand_16,
                  L1_0_L2_1_G1_MINI_ALU_BoothOperand_15,
                  L1_0_L2_1_G1_MINI_ALU_BoothOperand_14,
                  L1_0_L2_1_G1_MINI_ALU_BoothOperand_13,
                  L1_0_L2_1_G1_MINI_ALU_BoothOperand_12,
                  L1_0_L2_1_G1_MINI_ALU_BoothOperand_11,
                  L1_0_L2_1_G1_MINI_ALU_BoothOperand_10,
                  L1_0_L2_1_G1_MINI_ALU_BoothOperand_9,\$dummy [44],\$dummy [45]
                  ,\$dummy [46],\$dummy [47],\$dummy [48],\$dummy [49],
                  \$dummy [50],\$dummy [51],\$dummy [52]}), .BoothP ({
                  L1_0_L2_1_G1_MINI_ALU_BoothP_16,
                  L1_0_L2_1_G1_MINI_ALU_BoothP_15,
                  L1_0_L2_1_G1_MINI_ALU_BoothP_14,
                  L1_0_L2_1_G1_MINI_ALU_BoothP_13,
                  L1_0_L2_1_G1_MINI_ALU_BoothP_12,
                  L1_0_L2_1_G1_MINI_ALU_BoothP_11,
                  L1_0_L2_1_G1_MINI_ALU_BoothP_10,L1_0_L2_1_G1_MINI_ALU_BoothP_9
                  ,L1_0_L2_1_G1_MINI_ALU_BoothP_8,L1_0_L2_1_G1_MINI_ALU_BoothP_7
                  ,L1_0_L2_1_G1_MINI_ALU_BoothP_6,L1_0_L2_1_G1_MINI_ALU_BoothP_5
                  ,L1_0_L2_1_G1_MINI_ALU_BoothP_4,L1_0_L2_1_G1_MINI_ALU_BoothP_3
                  ,L1_0_L2_1_G1_MINI_ALU_BoothP_2,L1_0_L2_1_G1_MINI_ALU_BoothP_1
                  ,L1_0_L2_1_G1_MINI_ALU_BoothP_0}), .LargeWindowShifted ({
                  \$dummy [53],\$dummy [54],\$dummy [55],\$dummy [56],
                  \$dummy [57],\$dummy [58],\$dummy [59],\$dummy [60],
                  \$dummy [61],\$dummy [62],\$dummy [63],\$dummy [64],
                  \$dummy [65],\$dummy [66],\$dummy [67],\$dummy [68],
                  \$dummy [69]})) ;
    booth_adder_17 L1_0_L2_2_G1_MINI_ALU_BOOTH_ADDER (.AdderFirstOperand ({
                   L1FirstOperands_12__16,L1FirstOperands_2__15,
                   L1FirstOperands_2__14,L1FirstOperands_2__13,
                   L1FirstOperands_2__12,L1FirstOperands_2__11,
                   L1FirstOperands_2__10,L1FirstOperands_2__9,
                   L1FirstOperands_2__8,L1FirstOperands_2__7,
                   L1FirstOperands_2__6,L1FirstOperands_2__5,
                   L1FirstOperands_2__4,L1FirstOperands_2__3,
                   L1FirstOperands_2__2,L1FirstOperands_2__1,
                   L1FirstOperands_2__0}), .AdderSecondOperand ({
                   L1FirstOperands_12__16,
                   L1_0_L2_2_G1_MINI_ALU_OperationResult_15,
                   L1_0_L2_2_G1_MINI_ALU_OperationResult_14,
                   L1_0_L2_2_G1_MINI_ALU_OperationResult_13,
                   L1_0_L2_2_G1_MINI_ALU_OperationResult_12,
                   L1_0_L2_2_G1_MINI_ALU_OperationResult_11,
                   L1_0_L2_2_G1_MINI_ALU_OperationResult_10,
                   L1_0_L2_2_G1_MINI_ALU_OperationResult_9,
                   L1_0_L2_2_G1_MINI_ALU_OperationResult_8,
                   L1_0_L2_2_G1_MINI_ALU_OperationResult_7,
                   L1_0_L2_2_G1_MINI_ALU_OperationResult_6,
                   L1_0_L2_2_G1_MINI_ALU_OperationResult_5,
                   L1_0_L2_2_G1_MINI_ALU_OperationResult_4,
                   L1_0_L2_2_G1_MINI_ALU_OperationResult_3,
                   L1_0_L2_2_G1_MINI_ALU_OperationResult_2,
                   L1_0_L2_2_G1_MINI_ALU_OperationResult_1,
                   L1_0_L2_2_G1_MINI_ALU_OperationResult_0}), .BoothOperand ({
                   L1_0_L2_2_G1_MINI_ALU_BoothOperand_16,
                   L1_0_L2_2_G1_MINI_ALU_BoothOperand_15,
                   L1_0_L2_2_G1_MINI_ALU_BoothOperand_14,
                   L1_0_L2_2_G1_MINI_ALU_BoothOperand_13,
                   L1_0_L2_2_G1_MINI_ALU_BoothOperand_12,
                   L1_0_L2_2_G1_MINI_ALU_BoothOperand_11,
                   L1_0_L2_2_G1_MINI_ALU_BoothOperand_10,
                   L1_0_L2_2_G1_MINI_ALU_BoothOperand_9,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16}), .BoothP ({
                   L1_0_L2_2_G1_MINI_ALU_BoothP_16,
                   L1_0_L2_2_G1_MINI_ALU_BoothP_15,
                   L1_0_L2_2_G1_MINI_ALU_BoothP_14,
                   L1_0_L2_2_G1_MINI_ALU_BoothP_13,
                   L1_0_L2_2_G1_MINI_ALU_BoothP_12,
                   L1_0_L2_2_G1_MINI_ALU_BoothP_11,
                   L1_0_L2_2_G1_MINI_ALU_BoothP_10,
                   L1_0_L2_2_G1_MINI_ALU_BoothP_9,L1_0_L2_2_G1_MINI_ALU_BoothP_8
                   ,L1_0_L2_2_G1_MINI_ALU_BoothP_7,
                   L1_0_L2_2_G1_MINI_ALU_BoothP_6,L1_0_L2_2_G1_MINI_ALU_BoothP_5
                   ,L1_0_L2_2_G1_MINI_ALU_BoothP_4,
                   L1_0_L2_2_G1_MINI_ALU_BoothP_3,L1_0_L2_2_G1_MINI_ALU_BoothP_2
                   ,L1_0_L2_2_G1_MINI_ALU_BoothP_1,
                   L1_0_L2_2_G1_MINI_ALU_BoothP_0}), .SelOperand (nx3283), .Operation (
                   L1_0_L2_2_G1_MINI_ALU_BoothXORCheck), .AdderResult ({
                   L1ResultsLarge_2__16,L1ResultsLarge_2__15,
                   L1ResultsLarge_2__14,L1ResultsLarge_2__13,
                   L1ResultsLarge_2__12,L1ResultsLarge_2__11,
                   L1ResultsLarge_2__10,L1ResultsLarge_2__9,L1ResultsLarge_2__8,
                   L1ResultsLarge_2__7,L1ResultsLarge_2__6,L1ResultsLarge_2__5,
                   L1ResultsLarge_2__4,L1ResultsLarge_2__3,L1ResultsLarge_2__2,
                   L1ResultsLarge_2__1,L1ResultsLarge_2__0}), .AdderBoothResult (
                   {\$dummy [70],L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_15,
                   L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_14,
                   L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_13,
                   L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_12,
                   L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_11,
                   L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_10,
                   L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_9,
                   L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_8,
                   L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_7,
                   L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_6,
                   L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_5,
                   L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_4,
                   L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_3,
                   L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_2,
                   L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_1,
                   L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_0})) ;
    booth_unit_17 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT (.CLK (CLK), .RST (RST), .Start (
                  Start), .Instr (Instr), .LoopingAndResultNotReady (nx3275), .Filter (
                  {FilterDin_0__2__7,FilterDin_0__2__6,FilterDin_0__2__5,
                  FilterDin_0__2__4,FilterDin_0__2__3,FilterDin_0__2__2,
                  FilterDin_0__2__1,FilterDin_0__2__0}), .Window ({
                  WindowDin_0__2__7,WindowDin_0__2__6,WindowDin_0__2__5,
                  WindowDin_0__2__4,WindowDin_0__2__3,WindowDin_0__2__2,
                  WindowDin_0__2__1,WindowDin_0__2__0}), .AdderBoothResult ({
                  L1FirstOperands_12__16,
                  L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_15,
                  L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_14,
                  L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_13,
                  L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_12,
                  L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_11,
                  L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_10,
                  L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_9,
                  L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_8,
                  L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_7,
                  L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_6,
                  L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_5,
                  L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_4,
                  L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_3,
                  L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_2,
                  L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_1,
                  L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_0}), .BoothXORCheck (
                  L1_0_L2_2_G1_MINI_ALU_BoothXORCheck), .BoothResult ({
                  \$dummy [71],\$dummy [72],\$dummy [73],\$dummy [74],
                  \$dummy [75],\$dummy [76],\$dummy [77],\$dummy [78]}), .BoothAddingOperand (
                  {L1_0_L2_2_G1_MINI_ALU_BoothOperand_16,
                  L1_0_L2_2_G1_MINI_ALU_BoothOperand_15,
                  L1_0_L2_2_G1_MINI_ALU_BoothOperand_14,
                  L1_0_L2_2_G1_MINI_ALU_BoothOperand_13,
                  L1_0_L2_2_G1_MINI_ALU_BoothOperand_12,
                  L1_0_L2_2_G1_MINI_ALU_BoothOperand_11,
                  L1_0_L2_2_G1_MINI_ALU_BoothOperand_10,
                  L1_0_L2_2_G1_MINI_ALU_BoothOperand_9,\$dummy [79],\$dummy [80]
                  ,\$dummy [81],\$dummy [82],\$dummy [83],\$dummy [84],
                  \$dummy [85],\$dummy [86],\$dummy [87]}), .BoothP ({
                  L1_0_L2_2_G1_MINI_ALU_BoothP_16,
                  L1_0_L2_2_G1_MINI_ALU_BoothP_15,
                  L1_0_L2_2_G1_MINI_ALU_BoothP_14,
                  L1_0_L2_2_G1_MINI_ALU_BoothP_13,
                  L1_0_L2_2_G1_MINI_ALU_BoothP_12,
                  L1_0_L2_2_G1_MINI_ALU_BoothP_11,
                  L1_0_L2_2_G1_MINI_ALU_BoothP_10,L1_0_L2_2_G1_MINI_ALU_BoothP_9
                  ,L1_0_L2_2_G1_MINI_ALU_BoothP_8,L1_0_L2_2_G1_MINI_ALU_BoothP_7
                  ,L1_0_L2_2_G1_MINI_ALU_BoothP_6,L1_0_L2_2_G1_MINI_ALU_BoothP_5
                  ,L1_0_L2_2_G1_MINI_ALU_BoothP_4,L1_0_L2_2_G1_MINI_ALU_BoothP_3
                  ,L1_0_L2_2_G1_MINI_ALU_BoothP_2,L1_0_L2_2_G1_MINI_ALU_BoothP_1
                  ,L1_0_L2_2_G1_MINI_ALU_BoothP_0}), .LargeWindowShifted ({
                  \$dummy [88],\$dummy [89],\$dummy [90],\$dummy [91],
                  \$dummy [92],\$dummy [93],\$dummy [94],\$dummy [95],
                  \$dummy [96],\$dummy [97],\$dummy [98],\$dummy [99],
                  \$dummy [100],\$dummy [101],\$dummy [102],\$dummy [103],
                  \$dummy [104]})) ;
    booth_adder_17 L1_0_L2_3_G1_MINI_ALU_BOOTH_ADDER (.AdderFirstOperand ({
                   L1FirstOperands_12__16,L1FirstOperands_3__15,
                   L1FirstOperands_3__14,L1FirstOperands_3__13,
                   L1FirstOperands_3__12,L1FirstOperands_3__11,
                   L1FirstOperands_3__10,L1FirstOperands_3__9,
                   L1FirstOperands_3__8,L1FirstOperands_3__7,
                   L1FirstOperands_3__6,L1FirstOperands_3__5,
                   L1FirstOperands_3__4,L1FirstOperands_3__3,
                   L1FirstOperands_3__2,L1FirstOperands_3__1,
                   L1FirstOperands_3__0}), .AdderSecondOperand ({
                   L1FirstOperands_12__16,
                   L1_0_L2_3_G1_MINI_ALU_OperationResult_15,
                   L1_0_L2_3_G1_MINI_ALU_OperationResult_14,
                   L1_0_L2_3_G1_MINI_ALU_OperationResult_13,
                   L1_0_L2_3_G1_MINI_ALU_OperationResult_12,
                   L1_0_L2_3_G1_MINI_ALU_OperationResult_11,
                   L1_0_L2_3_G1_MINI_ALU_OperationResult_10,
                   L1_0_L2_3_G1_MINI_ALU_OperationResult_9,
                   L1_0_L2_3_G1_MINI_ALU_OperationResult_8,
                   L1_0_L2_3_G1_MINI_ALU_OperationResult_7,
                   L1_0_L2_3_G1_MINI_ALU_OperationResult_6,
                   L1_0_L2_3_G1_MINI_ALU_OperationResult_5,
                   L1_0_L2_3_G1_MINI_ALU_OperationResult_4,
                   L1_0_L2_3_G1_MINI_ALU_OperationResult_3,
                   L1_0_L2_3_G1_MINI_ALU_OperationResult_2,
                   L1_0_L2_3_G1_MINI_ALU_OperationResult_1,
                   L1_0_L2_3_G1_MINI_ALU_OperationResult_0}), .BoothOperand ({
                   L1_0_L2_3_G1_MINI_ALU_BoothOperand_16,
                   L1_0_L2_3_G1_MINI_ALU_BoothOperand_15,
                   L1_0_L2_3_G1_MINI_ALU_BoothOperand_14,
                   L1_0_L2_3_G1_MINI_ALU_BoothOperand_13,
                   L1_0_L2_3_G1_MINI_ALU_BoothOperand_12,
                   L1_0_L2_3_G1_MINI_ALU_BoothOperand_11,
                   L1_0_L2_3_G1_MINI_ALU_BoothOperand_10,
                   L1_0_L2_3_G1_MINI_ALU_BoothOperand_9,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16}), .BoothP ({
                   L1_0_L2_3_G1_MINI_ALU_BoothP_16,
                   L1_0_L2_3_G1_MINI_ALU_BoothP_15,
                   L1_0_L2_3_G1_MINI_ALU_BoothP_14,
                   L1_0_L2_3_G1_MINI_ALU_BoothP_13,
                   L1_0_L2_3_G1_MINI_ALU_BoothP_12,
                   L1_0_L2_3_G1_MINI_ALU_BoothP_11,
                   L1_0_L2_3_G1_MINI_ALU_BoothP_10,
                   L1_0_L2_3_G1_MINI_ALU_BoothP_9,L1_0_L2_3_G1_MINI_ALU_BoothP_8
                   ,L1_0_L2_3_G1_MINI_ALU_BoothP_7,
                   L1_0_L2_3_G1_MINI_ALU_BoothP_6,L1_0_L2_3_G1_MINI_ALU_BoothP_5
                   ,L1_0_L2_3_G1_MINI_ALU_BoothP_4,
                   L1_0_L2_3_G1_MINI_ALU_BoothP_3,L1_0_L2_3_G1_MINI_ALU_BoothP_2
                   ,L1_0_L2_3_G1_MINI_ALU_BoothP_1,
                   L1_0_L2_3_G1_MINI_ALU_BoothP_0}), .SelOperand (nx3283), .Operation (
                   L1_0_L2_3_G1_MINI_ALU_BoothXORCheck), .AdderResult ({
                   L1ResultsLarge_3__16,L1ResultsLarge_3__15,
                   L1ResultsLarge_3__14,L1ResultsLarge_3__13,
                   L1ResultsLarge_3__12,L1ResultsLarge_3__11,
                   L1ResultsLarge_3__10,L1ResultsLarge_3__9,L1ResultsLarge_3__8,
                   L1ResultsLarge_3__7,L1ResultsLarge_3__6,L1ResultsLarge_3__5,
                   L1ResultsLarge_3__4,L1ResultsLarge_3__3,L1ResultsLarge_3__2,
                   L1ResultsLarge_3__1,L1ResultsLarge_3__0}), .AdderBoothResult (
                   {\$dummy [105],L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_15,
                   L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_14,
                   L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_13,
                   L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_12,
                   L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_11,
                   L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_10,
                   L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_9,
                   L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_8,
                   L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_7,
                   L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_6,
                   L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_5,
                   L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_4,
                   L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_3,
                   L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_2,
                   L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_1,
                   L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_0})) ;
    booth_unit_17 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT (.CLK (CLK), .RST (RST), .Start (
                  Start), .Instr (Instr), .LoopingAndResultNotReady (nx3275), .Filter (
                  {FilterDin_0__3__7,FilterDin_0__3__6,FilterDin_0__3__5,
                  FilterDin_0__3__4,FilterDin_0__3__3,FilterDin_0__3__2,
                  FilterDin_0__3__1,FilterDin_0__3__0}), .Window ({
                  WindowDin_0__3__7,WindowDin_0__3__6,WindowDin_0__3__5,
                  WindowDin_0__3__4,WindowDin_0__3__3,WindowDin_0__3__2,
                  WindowDin_0__3__1,WindowDin_0__3__0}), .AdderBoothResult ({
                  L1FirstOperands_12__16,
                  L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_15,
                  L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_14,
                  L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_13,
                  L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_12,
                  L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_11,
                  L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_10,
                  L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_9,
                  L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_8,
                  L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_7,
                  L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_6,
                  L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_5,
                  L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_4,
                  L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_3,
                  L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_2,
                  L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_1,
                  L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_0}), .BoothXORCheck (
                  L1_0_L2_3_G1_MINI_ALU_BoothXORCheck), .BoothResult ({
                  \$dummy [106],\$dummy [107],\$dummy [108],\$dummy [109],
                  \$dummy [110],\$dummy [111],\$dummy [112],\$dummy [113]}), .BoothAddingOperand (
                  {L1_0_L2_3_G1_MINI_ALU_BoothOperand_16,
                  L1_0_L2_3_G1_MINI_ALU_BoothOperand_15,
                  L1_0_L2_3_G1_MINI_ALU_BoothOperand_14,
                  L1_0_L2_3_G1_MINI_ALU_BoothOperand_13,
                  L1_0_L2_3_G1_MINI_ALU_BoothOperand_12,
                  L1_0_L2_3_G1_MINI_ALU_BoothOperand_11,
                  L1_0_L2_3_G1_MINI_ALU_BoothOperand_10,
                  L1_0_L2_3_G1_MINI_ALU_BoothOperand_9,\$dummy [114],
                  \$dummy [115],\$dummy [116],\$dummy [117],\$dummy [118],
                  \$dummy [119],\$dummy [120],\$dummy [121],\$dummy [122]}), .BoothP (
                  {L1_0_L2_3_G1_MINI_ALU_BoothP_16,
                  L1_0_L2_3_G1_MINI_ALU_BoothP_15,
                  L1_0_L2_3_G1_MINI_ALU_BoothP_14,
                  L1_0_L2_3_G1_MINI_ALU_BoothP_13,
                  L1_0_L2_3_G1_MINI_ALU_BoothP_12,
                  L1_0_L2_3_G1_MINI_ALU_BoothP_11,
                  L1_0_L2_3_G1_MINI_ALU_BoothP_10,L1_0_L2_3_G1_MINI_ALU_BoothP_9
                  ,L1_0_L2_3_G1_MINI_ALU_BoothP_8,L1_0_L2_3_G1_MINI_ALU_BoothP_7
                  ,L1_0_L2_3_G1_MINI_ALU_BoothP_6,L1_0_L2_3_G1_MINI_ALU_BoothP_5
                  ,L1_0_L2_3_G1_MINI_ALU_BoothP_4,L1_0_L2_3_G1_MINI_ALU_BoothP_3
                  ,L1_0_L2_3_G1_MINI_ALU_BoothP_2,L1_0_L2_3_G1_MINI_ALU_BoothP_1
                  ,L1_0_L2_3_G1_MINI_ALU_BoothP_0}), .LargeWindowShifted ({
                  \$dummy [123],\$dummy [124],\$dummy [125],\$dummy [126],
                  \$dummy [127],\$dummy [128],\$dummy [129],\$dummy [130],
                  \$dummy [131],\$dummy [132],\$dummy [133],\$dummy [134],
                  \$dummy [135],\$dummy [136],\$dummy [137],\$dummy [138],
                  \$dummy [139]})) ;
    booth_adder_17 L1_0_L2_4_G1_MINI_ALU_BOOTH_ADDER (.AdderFirstOperand ({
                   L1FirstOperands_12__16,L1FirstOperands_4__15,
                   L1FirstOperands_4__14,L1FirstOperands_4__13,
                   L1FirstOperands_4__12,L1FirstOperands_4__11,
                   L1FirstOperands_4__10,L1FirstOperands_4__9,
                   L1FirstOperands_4__8,L1FirstOperands_4__7,
                   L1FirstOperands_4__6,L1FirstOperands_4__5,
                   L1FirstOperands_4__4,L1FirstOperands_4__3,
                   L1FirstOperands_4__2,L1FirstOperands_4__1,
                   L1FirstOperands_4__0}), .AdderSecondOperand ({
                   L1FirstOperands_12__16,
                   L1_0_L2_4_G1_MINI_ALU_OperationResult_15,
                   L1_0_L2_4_G1_MINI_ALU_OperationResult_14,
                   L1_0_L2_4_G1_MINI_ALU_OperationResult_13,
                   L1_0_L2_4_G1_MINI_ALU_OperationResult_12,
                   L1_0_L2_4_G1_MINI_ALU_OperationResult_11,
                   L1_0_L2_4_G1_MINI_ALU_OperationResult_10,
                   L1_0_L2_4_G1_MINI_ALU_OperationResult_9,
                   L1_0_L2_4_G1_MINI_ALU_OperationResult_8,
                   L1_0_L2_4_G1_MINI_ALU_OperationResult_7,
                   L1_0_L2_4_G1_MINI_ALU_OperationResult_6,
                   L1_0_L2_4_G1_MINI_ALU_OperationResult_5,
                   L1_0_L2_4_G1_MINI_ALU_OperationResult_4,
                   L1_0_L2_4_G1_MINI_ALU_OperationResult_3,
                   L1_0_L2_4_G1_MINI_ALU_OperationResult_2,
                   L1_0_L2_4_G1_MINI_ALU_OperationResult_1,
                   L1_0_L2_4_G1_MINI_ALU_OperationResult_0}), .BoothOperand ({
                   L1_0_L2_4_G1_MINI_ALU_BoothOperand_16,
                   L1_0_L2_4_G1_MINI_ALU_BoothOperand_15,
                   L1_0_L2_4_G1_MINI_ALU_BoothOperand_14,
                   L1_0_L2_4_G1_MINI_ALU_BoothOperand_13,
                   L1_0_L2_4_G1_MINI_ALU_BoothOperand_12,
                   L1_0_L2_4_G1_MINI_ALU_BoothOperand_11,
                   L1_0_L2_4_G1_MINI_ALU_BoothOperand_10,
                   L1_0_L2_4_G1_MINI_ALU_BoothOperand_9,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16}), .BoothP ({
                   L1_0_L2_4_G1_MINI_ALU_BoothP_16,
                   L1_0_L2_4_G1_MINI_ALU_BoothP_15,
                   L1_0_L2_4_G1_MINI_ALU_BoothP_14,
                   L1_0_L2_4_G1_MINI_ALU_BoothP_13,
                   L1_0_L2_4_G1_MINI_ALU_BoothP_12,
                   L1_0_L2_4_G1_MINI_ALU_BoothP_11,
                   L1_0_L2_4_G1_MINI_ALU_BoothP_10,
                   L1_0_L2_4_G1_MINI_ALU_BoothP_9,L1_0_L2_4_G1_MINI_ALU_BoothP_8
                   ,L1_0_L2_4_G1_MINI_ALU_BoothP_7,
                   L1_0_L2_4_G1_MINI_ALU_BoothP_6,L1_0_L2_4_G1_MINI_ALU_BoothP_5
                   ,L1_0_L2_4_G1_MINI_ALU_BoothP_4,
                   L1_0_L2_4_G1_MINI_ALU_BoothP_3,L1_0_L2_4_G1_MINI_ALU_BoothP_2
                   ,L1_0_L2_4_G1_MINI_ALU_BoothP_1,
                   L1_0_L2_4_G1_MINI_ALU_BoothP_0}), .SelOperand (nx3283), .Operation (
                   L1_0_L2_4_G1_MINI_ALU_BoothXORCheck), .AdderResult ({
                   L1ResultsLarge_4__16,L1ResultsLarge_4__15,
                   L1ResultsLarge_4__14,L1ResultsLarge_4__13,
                   L1ResultsLarge_4__12,L1ResultsLarge_4__11,
                   L1ResultsLarge_4__10,L1ResultsLarge_4__9,L1ResultsLarge_4__8,
                   L1ResultsLarge_4__7,L1ResultsLarge_4__6,L1ResultsLarge_4__5,
                   L1ResultsLarge_4__4,L1ResultsLarge_4__3,L1ResultsLarge_4__2,
                   L1ResultsLarge_4__1,L1ResultsLarge_4__0}), .AdderBoothResult (
                   {\$dummy [140],L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_15,
                   L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_14,
                   L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_13,
                   L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_12,
                   L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_11,
                   L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_10,
                   L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_9,
                   L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_8,
                   L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_7,
                   L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_6,
                   L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_5,
                   L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_4,
                   L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_3,
                   L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_2,
                   L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_1,
                   L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_0})) ;
    booth_unit_17 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT (.CLK (CLK), .RST (RST), .Start (
                  Start), .Instr (Instr), .LoopingAndResultNotReady (nx3275), .Filter (
                  {FilterDin_0__4__7,FilterDin_0__4__6,FilterDin_0__4__5,
                  FilterDin_0__4__4,FilterDin_0__4__3,FilterDin_0__4__2,
                  FilterDin_0__4__1,FilterDin_0__4__0}), .Window ({
                  WindowDin_0__4__7,WindowDin_0__4__6,WindowDin_0__4__5,
                  WindowDin_0__4__4,WindowDin_0__4__3,WindowDin_0__4__2,
                  WindowDin_0__4__1,WindowDin_0__4__0}), .AdderBoothResult ({
                  L1FirstOperands_12__16,
                  L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_15,
                  L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_14,
                  L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_13,
                  L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_12,
                  L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_11,
                  L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_10,
                  L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_9,
                  L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_8,
                  L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_7,
                  L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_6,
                  L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_5,
                  L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_4,
                  L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_3,
                  L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_2,
                  L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_1,
                  L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_0}), .BoothXORCheck (
                  L1_0_L2_4_G1_MINI_ALU_BoothXORCheck), .BoothResult ({
                  \$dummy [141],\$dummy [142],\$dummy [143],\$dummy [144],
                  \$dummy [145],\$dummy [146],\$dummy [147],\$dummy [148]}), .BoothAddingOperand (
                  {L1_0_L2_4_G1_MINI_ALU_BoothOperand_16,
                  L1_0_L2_4_G1_MINI_ALU_BoothOperand_15,
                  L1_0_L2_4_G1_MINI_ALU_BoothOperand_14,
                  L1_0_L2_4_G1_MINI_ALU_BoothOperand_13,
                  L1_0_L2_4_G1_MINI_ALU_BoothOperand_12,
                  L1_0_L2_4_G1_MINI_ALU_BoothOperand_11,
                  L1_0_L2_4_G1_MINI_ALU_BoothOperand_10,
                  L1_0_L2_4_G1_MINI_ALU_BoothOperand_9,\$dummy [149],
                  \$dummy [150],\$dummy [151],\$dummy [152],\$dummy [153],
                  \$dummy [154],\$dummy [155],\$dummy [156],\$dummy [157]}), .BoothP (
                  {L1_0_L2_4_G1_MINI_ALU_BoothP_16,
                  L1_0_L2_4_G1_MINI_ALU_BoothP_15,
                  L1_0_L2_4_G1_MINI_ALU_BoothP_14,
                  L1_0_L2_4_G1_MINI_ALU_BoothP_13,
                  L1_0_L2_4_G1_MINI_ALU_BoothP_12,
                  L1_0_L2_4_G1_MINI_ALU_BoothP_11,
                  L1_0_L2_4_G1_MINI_ALU_BoothP_10,L1_0_L2_4_G1_MINI_ALU_BoothP_9
                  ,L1_0_L2_4_G1_MINI_ALU_BoothP_8,L1_0_L2_4_G1_MINI_ALU_BoothP_7
                  ,L1_0_L2_4_G1_MINI_ALU_BoothP_6,L1_0_L2_4_G1_MINI_ALU_BoothP_5
                  ,L1_0_L2_4_G1_MINI_ALU_BoothP_4,L1_0_L2_4_G1_MINI_ALU_BoothP_3
                  ,L1_0_L2_4_G1_MINI_ALU_BoothP_2,L1_0_L2_4_G1_MINI_ALU_BoothP_1
                  ,L1_0_L2_4_G1_MINI_ALU_BoothP_0}), .LargeWindowShifted ({
                  \$dummy [158],\$dummy [159],\$dummy [160],\$dummy [161],
                  \$dummy [162],\$dummy [163],\$dummy [164],\$dummy [165],
                  \$dummy [166],\$dummy [167],\$dummy [168],\$dummy [169],
                  \$dummy [170],\$dummy [171],\$dummy [172],\$dummy [173],
                  \$dummy [174]})) ;
    booth_adder_17 L1_1_L2_0_G1_MINI_ALU_BOOTH_ADDER (.AdderFirstOperand ({
                   L1FirstOperands_12__16,L1FirstOperands_2__15,
                   L1FirstOperands_2__14,L1FirstOperands_2__13,
                   L1FirstOperands_2__12,L1FirstOperands_2__11,
                   L1FirstOperands_2__10,L1FirstOperands_2__9,
                   L1FirstOperands_2__8,L1FirstOperands_2__7,
                   L1FirstOperands_2__6,L1FirstOperands_2__5,
                   L1FirstOperands_2__4,L1FirstOperands_2__3,
                   L1FirstOperands_2__2,L1FirstOperands_2__1,
                   L1FirstOperands_2__0}), .AdderSecondOperand ({
                   L1FirstOperands_12__16,
                   L1_1_L2_0_G1_MINI_ALU_OperationResult_15,
                   L1_1_L2_0_G1_MINI_ALU_OperationResult_14,
                   L1_1_L2_0_G1_MINI_ALU_OperationResult_13,
                   L1_1_L2_0_G1_MINI_ALU_OperationResult_12,
                   L1_1_L2_0_G1_MINI_ALU_OperationResult_11,
                   L1_1_L2_0_G1_MINI_ALU_OperationResult_10,
                   L1_1_L2_0_G1_MINI_ALU_OperationResult_9,
                   L1_1_L2_0_G1_MINI_ALU_OperationResult_8,
                   L1_1_L2_0_G1_MINI_ALU_OperationResult_7,
                   L1_1_L2_0_G1_MINI_ALU_OperationResult_6,
                   L1_1_L2_0_G1_MINI_ALU_OperationResult_5,
                   L1_1_L2_0_G1_MINI_ALU_OperationResult_4,
                   L1_1_L2_0_G1_MINI_ALU_OperationResult_3,
                   L1_1_L2_0_G1_MINI_ALU_OperationResult_2,
                   L1_1_L2_0_G1_MINI_ALU_OperationResult_1,
                   L1_1_L2_0_G1_MINI_ALU_OperationResult_0}), .BoothOperand ({
                   L1_1_L2_0_G1_MINI_ALU_BoothOperand_16,
                   L1_1_L2_0_G1_MINI_ALU_BoothOperand_15,
                   L1_1_L2_0_G1_MINI_ALU_BoothOperand_14,
                   L1_1_L2_0_G1_MINI_ALU_BoothOperand_13,
                   L1_1_L2_0_G1_MINI_ALU_BoothOperand_12,
                   L1_1_L2_0_G1_MINI_ALU_BoothOperand_11,
                   L1_1_L2_0_G1_MINI_ALU_BoothOperand_10,
                   L1_1_L2_0_G1_MINI_ALU_BoothOperand_9,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16}), .BoothP ({
                   L1_1_L2_0_G1_MINI_ALU_BoothP_16,
                   L1_1_L2_0_G1_MINI_ALU_BoothP_15,
                   L1_1_L2_0_G1_MINI_ALU_BoothP_14,
                   L1_1_L2_0_G1_MINI_ALU_BoothP_13,
                   L1_1_L2_0_G1_MINI_ALU_BoothP_12,
                   L1_1_L2_0_G1_MINI_ALU_BoothP_11,
                   L1_1_L2_0_G1_MINI_ALU_BoothP_10,
                   L1_1_L2_0_G1_MINI_ALU_BoothP_9,L1_1_L2_0_G1_MINI_ALU_BoothP_8
                   ,L1_1_L2_0_G1_MINI_ALU_BoothP_7,
                   L1_1_L2_0_G1_MINI_ALU_BoothP_6,L1_1_L2_0_G1_MINI_ALU_BoothP_5
                   ,L1_1_L2_0_G1_MINI_ALU_BoothP_4,
                   L1_1_L2_0_G1_MINI_ALU_BoothP_3,L1_1_L2_0_G1_MINI_ALU_BoothP_2
                   ,L1_1_L2_0_G1_MINI_ALU_BoothP_1,
                   L1_1_L2_0_G1_MINI_ALU_BoothP_0}), .SelOperand (nx3283), .Operation (
                   L1_1_L2_0_G1_MINI_ALU_BoothXORCheck), .AdderResult ({
                   L1ResultsLarge_5__16,L1ResultsLarge_5__15,
                   L1ResultsLarge_5__14,L1ResultsLarge_5__13,
                   L1ResultsLarge_5__12,L1ResultsLarge_5__11,
                   L1ResultsLarge_5__10,L1ResultsLarge_5__9,L1ResultsLarge_5__8,
                   L1ResultsLarge_5__7,L1ResultsLarge_5__6,L1ResultsLarge_5__5,
                   L1ResultsLarge_5__4,L1ResultsLarge_5__3,L1ResultsLarge_5__2,
                   L1ResultsLarge_5__1,L1ResultsLarge_5__0}), .AdderBoothResult (
                   {\$dummy [175],L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_15,
                   L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_14,
                   L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_13,
                   L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_12,
                   L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_11,
                   L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_10,
                   L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_9,
                   L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_8,
                   L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_7,
                   L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_6,
                   L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_5,
                   L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_4,
                   L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_3,
                   L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_2,
                   L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_1,
                   L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_0})) ;
    booth_unit_17 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT (.CLK (CLK), .RST (RST), .Start (
                  Start), .Instr (Instr), .LoopingAndResultNotReady (nx3275), .Filter (
                  {FilterDin_1__0__7,FilterDin_1__0__6,FilterDin_1__0__5,
                  FilterDin_1__0__4,FilterDin_1__0__3,FilterDin_1__0__2,
                  FilterDin_1__0__1,FilterDin_1__0__0}), .Window ({
                  WindowDin_1__0__7,WindowDin_1__0__6,WindowDin_1__0__5,
                  WindowDin_1__0__4,WindowDin_1__0__3,WindowDin_1__0__2,
                  WindowDin_1__0__1,WindowDin_1__0__0}), .AdderBoothResult ({
                  L1FirstOperands_12__16,
                  L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_15,
                  L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_14,
                  L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_13,
                  L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_12,
                  L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_11,
                  L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_10,
                  L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_9,
                  L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_8,
                  L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_7,
                  L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_6,
                  L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_5,
                  L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_4,
                  L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_3,
                  L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_2,
                  L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_1,
                  L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_0}), .BoothXORCheck (
                  L1_1_L2_0_G1_MINI_ALU_BoothXORCheck), .BoothResult ({
                  \$dummy [176],\$dummy [177],\$dummy [178],\$dummy [179],
                  \$dummy [180],\$dummy [181],\$dummy [182],\$dummy [183]}), .BoothAddingOperand (
                  {L1_1_L2_0_G1_MINI_ALU_BoothOperand_16,
                  L1_1_L2_0_G1_MINI_ALU_BoothOperand_15,
                  L1_1_L2_0_G1_MINI_ALU_BoothOperand_14,
                  L1_1_L2_0_G1_MINI_ALU_BoothOperand_13,
                  L1_1_L2_0_G1_MINI_ALU_BoothOperand_12,
                  L1_1_L2_0_G1_MINI_ALU_BoothOperand_11,
                  L1_1_L2_0_G1_MINI_ALU_BoothOperand_10,
                  L1_1_L2_0_G1_MINI_ALU_BoothOperand_9,\$dummy [184],
                  \$dummy [185],\$dummy [186],\$dummy [187],\$dummy [188],
                  \$dummy [189],\$dummy [190],\$dummy [191],\$dummy [192]}), .BoothP (
                  {L1_1_L2_0_G1_MINI_ALU_BoothP_16,
                  L1_1_L2_0_G1_MINI_ALU_BoothP_15,
                  L1_1_L2_0_G1_MINI_ALU_BoothP_14,
                  L1_1_L2_0_G1_MINI_ALU_BoothP_13,
                  L1_1_L2_0_G1_MINI_ALU_BoothP_12,
                  L1_1_L2_0_G1_MINI_ALU_BoothP_11,
                  L1_1_L2_0_G1_MINI_ALU_BoothP_10,L1_1_L2_0_G1_MINI_ALU_BoothP_9
                  ,L1_1_L2_0_G1_MINI_ALU_BoothP_8,L1_1_L2_0_G1_MINI_ALU_BoothP_7
                  ,L1_1_L2_0_G1_MINI_ALU_BoothP_6,L1_1_L2_0_G1_MINI_ALU_BoothP_5
                  ,L1_1_L2_0_G1_MINI_ALU_BoothP_4,L1_1_L2_0_G1_MINI_ALU_BoothP_3
                  ,L1_1_L2_0_G1_MINI_ALU_BoothP_2,L1_1_L2_0_G1_MINI_ALU_BoothP_1
                  ,L1_1_L2_0_G1_MINI_ALU_BoothP_0}), .LargeWindowShifted ({
                  \$dummy [193],\$dummy [194],\$dummy [195],\$dummy [196],
                  \$dummy [197],\$dummy [198],\$dummy [199],\$dummy [200],
                  \$dummy [201],\$dummy [202],\$dummy [203],\$dummy [204],
                  \$dummy [205],\$dummy [206],\$dummy [207],\$dummy [208],
                  \$dummy [209]})) ;
    booth_adder_17 L1_1_L2_1_G1_MINI_ALU_BOOTH_ADDER (.AdderFirstOperand ({
                   L1FirstOperands_12__16,L1FirstOperands_6__15,
                   L1FirstOperands_6__14,L1FirstOperands_6__13,
                   L1FirstOperands_6__12,L1FirstOperands_6__11,
                   L1FirstOperands_6__10,L1FirstOperands_6__9,
                   L1FirstOperands_6__8,L1FirstOperands_6__7,
                   L1FirstOperands_6__6,L1FirstOperands_6__5,
                   L1FirstOperands_6__4,L1FirstOperands_6__3,
                   L1FirstOperands_6__2,L1FirstOperands_6__1,
                   L1FirstOperands_6__0}), .AdderSecondOperand ({
                   L1FirstOperands_12__16,
                   L1_1_L2_1_G1_MINI_ALU_OperationResult_15,
                   L1_1_L2_1_G1_MINI_ALU_OperationResult_14,
                   L1_1_L2_1_G1_MINI_ALU_OperationResult_13,
                   L1_1_L2_1_G1_MINI_ALU_OperationResult_12,
                   L1_1_L2_1_G1_MINI_ALU_OperationResult_11,
                   L1_1_L2_1_G1_MINI_ALU_OperationResult_10,
                   L1_1_L2_1_G1_MINI_ALU_OperationResult_9,
                   L1_1_L2_1_G1_MINI_ALU_OperationResult_8,
                   L1_1_L2_1_G1_MINI_ALU_OperationResult_7,
                   L1_1_L2_1_G1_MINI_ALU_OperationResult_6,
                   L1_1_L2_1_G1_MINI_ALU_OperationResult_5,
                   L1_1_L2_1_G1_MINI_ALU_OperationResult_4,
                   L1_1_L2_1_G1_MINI_ALU_OperationResult_3,
                   L1_1_L2_1_G1_MINI_ALU_OperationResult_2,
                   L1_1_L2_1_G1_MINI_ALU_OperationResult_1,
                   L1_1_L2_1_G1_MINI_ALU_OperationResult_0}), .BoothOperand ({
                   L1_1_L2_1_G1_MINI_ALU_BoothOperand_16,
                   L1_1_L2_1_G1_MINI_ALU_BoothOperand_15,
                   L1_1_L2_1_G1_MINI_ALU_BoothOperand_14,
                   L1_1_L2_1_G1_MINI_ALU_BoothOperand_13,
                   L1_1_L2_1_G1_MINI_ALU_BoothOperand_12,
                   L1_1_L2_1_G1_MINI_ALU_BoothOperand_11,
                   L1_1_L2_1_G1_MINI_ALU_BoothOperand_10,
                   L1_1_L2_1_G1_MINI_ALU_BoothOperand_9,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16}), .BoothP ({
                   L1_1_L2_1_G1_MINI_ALU_BoothP_16,
                   L1_1_L2_1_G1_MINI_ALU_BoothP_15,
                   L1_1_L2_1_G1_MINI_ALU_BoothP_14,
                   L1_1_L2_1_G1_MINI_ALU_BoothP_13,
                   L1_1_L2_1_G1_MINI_ALU_BoothP_12,
                   L1_1_L2_1_G1_MINI_ALU_BoothP_11,
                   L1_1_L2_1_G1_MINI_ALU_BoothP_10,
                   L1_1_L2_1_G1_MINI_ALU_BoothP_9,L1_1_L2_1_G1_MINI_ALU_BoothP_8
                   ,L1_1_L2_1_G1_MINI_ALU_BoothP_7,
                   L1_1_L2_1_G1_MINI_ALU_BoothP_6,L1_1_L2_1_G1_MINI_ALU_BoothP_5
                   ,L1_1_L2_1_G1_MINI_ALU_BoothP_4,
                   L1_1_L2_1_G1_MINI_ALU_BoothP_3,L1_1_L2_1_G1_MINI_ALU_BoothP_2
                   ,L1_1_L2_1_G1_MINI_ALU_BoothP_1,
                   L1_1_L2_1_G1_MINI_ALU_BoothP_0}), .SelOperand (nx3283), .Operation (
                   L1_1_L2_1_G1_MINI_ALU_BoothXORCheck), .AdderResult ({
                   L1ResultsLarge_6__16,L1ResultsLarge_6__15,
                   L1ResultsLarge_6__14,L1ResultsLarge_6__13,
                   L1ResultsLarge_6__12,L1ResultsLarge_6__11,
                   L1ResultsLarge_6__10,L1ResultsLarge_6__9,L1ResultsLarge_6__8,
                   L1ResultsLarge_6__7,L1ResultsLarge_6__6,L1ResultsLarge_6__5,
                   L1ResultsLarge_6__4,L1ResultsLarge_6__3,L1ResultsLarge_6__2,
                   L1ResultsLarge_6__1,L1ResultsLarge_6__0}), .AdderBoothResult (
                   {\$dummy [210],L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_15,
                   L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_14,
                   L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_13,
                   L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_12,
                   L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_11,
                   L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_10,
                   L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_9,
                   L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_8,
                   L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_7,
                   L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_6,
                   L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_5,
                   L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_4,
                   L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_3,
                   L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_2,
                   L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_1,
                   L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_0})) ;
    booth_unit_17 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT (.CLK (CLK), .RST (RST), .Start (
                  Start), .Instr (Instr), .LoopingAndResultNotReady (nx3275), .Filter (
                  {FilterDin_1__1__7,FilterDin_1__1__6,FilterDin_1__1__5,
                  FilterDin_1__1__4,FilterDin_1__1__3,FilterDin_1__1__2,
                  FilterDin_1__1__1,FilterDin_1__1__0}), .Window ({
                  WindowDin_1__1__7,WindowDin_1__1__6,WindowDin_1__1__5,
                  WindowDin_1__1__4,WindowDin_1__1__3,WindowDin_1__1__2,
                  WindowDin_1__1__1,WindowDin_1__1__0}), .AdderBoothResult ({
                  L1FirstOperands_12__16,
                  L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_15,
                  L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_14,
                  L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_13,
                  L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_12,
                  L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_11,
                  L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_10,
                  L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_9,
                  L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_8,
                  L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_7,
                  L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_6,
                  L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_5,
                  L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_4,
                  L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_3,
                  L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_2,
                  L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_1,
                  L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_0}), .BoothXORCheck (
                  L1_1_L2_1_G1_MINI_ALU_BoothXORCheck), .BoothResult ({
                  \$dummy [211],\$dummy [212],\$dummy [213],\$dummy [214],
                  \$dummy [215],\$dummy [216],\$dummy [217],\$dummy [218]}), .BoothAddingOperand (
                  {L1_1_L2_1_G1_MINI_ALU_BoothOperand_16,
                  L1_1_L2_1_G1_MINI_ALU_BoothOperand_15,
                  L1_1_L2_1_G1_MINI_ALU_BoothOperand_14,
                  L1_1_L2_1_G1_MINI_ALU_BoothOperand_13,
                  L1_1_L2_1_G1_MINI_ALU_BoothOperand_12,
                  L1_1_L2_1_G1_MINI_ALU_BoothOperand_11,
                  L1_1_L2_1_G1_MINI_ALU_BoothOperand_10,
                  L1_1_L2_1_G1_MINI_ALU_BoothOperand_9,\$dummy [219],
                  \$dummy [220],\$dummy [221],\$dummy [222],\$dummy [223],
                  \$dummy [224],\$dummy [225],\$dummy [226],\$dummy [227]}), .BoothP (
                  {L1_1_L2_1_G1_MINI_ALU_BoothP_16,
                  L1_1_L2_1_G1_MINI_ALU_BoothP_15,
                  L1_1_L2_1_G1_MINI_ALU_BoothP_14,
                  L1_1_L2_1_G1_MINI_ALU_BoothP_13,
                  L1_1_L2_1_G1_MINI_ALU_BoothP_12,
                  L1_1_L2_1_G1_MINI_ALU_BoothP_11,
                  L1_1_L2_1_G1_MINI_ALU_BoothP_10,L1_1_L2_1_G1_MINI_ALU_BoothP_9
                  ,L1_1_L2_1_G1_MINI_ALU_BoothP_8,L1_1_L2_1_G1_MINI_ALU_BoothP_7
                  ,L1_1_L2_1_G1_MINI_ALU_BoothP_6,L1_1_L2_1_G1_MINI_ALU_BoothP_5
                  ,L1_1_L2_1_G1_MINI_ALU_BoothP_4,L1_1_L2_1_G1_MINI_ALU_BoothP_3
                  ,L1_1_L2_1_G1_MINI_ALU_BoothP_2,L1_1_L2_1_G1_MINI_ALU_BoothP_1
                  ,L1_1_L2_1_G1_MINI_ALU_BoothP_0}), .LargeWindowShifted ({
                  \$dummy [228],\$dummy [229],\$dummy [230],\$dummy [231],
                  \$dummy [232],\$dummy [233],\$dummy [234],\$dummy [235],
                  \$dummy [236],\$dummy [237],\$dummy [238],\$dummy [239],
                  \$dummy [240],\$dummy [241],\$dummy [242],\$dummy [243],
                  \$dummy [244]})) ;
    booth_adder_17 L1_1_L2_2_G1_MINI_ALU_BOOTH_ADDER (.AdderFirstOperand ({
                   L1FirstOperands_12__16,L1FirstOperands_7__15,
                   L1FirstOperands_7__14,L1FirstOperands_7__13,
                   L1FirstOperands_7__12,L1FirstOperands_7__11,
                   L1FirstOperands_7__10,L1FirstOperands_7__9,
                   L1FirstOperands_7__8,L1FirstOperands_7__7,
                   L1FirstOperands_7__6,L1FirstOperands_7__5,
                   L1FirstOperands_7__4,L1FirstOperands_7__3,
                   L1FirstOperands_7__2,L1FirstOperands_7__1,
                   L1FirstOperands_7__0}), .AdderSecondOperand ({
                   L1FirstOperands_12__16,
                   L1_1_L2_2_G1_MINI_ALU_OperationResult_15,
                   L1_1_L2_2_G1_MINI_ALU_OperationResult_14,
                   L1_1_L2_2_G1_MINI_ALU_OperationResult_13,
                   L1_1_L2_2_G1_MINI_ALU_OperationResult_12,
                   L1_1_L2_2_G1_MINI_ALU_OperationResult_11,
                   L1_1_L2_2_G1_MINI_ALU_OperationResult_10,
                   L1_1_L2_2_G1_MINI_ALU_OperationResult_9,
                   L1_1_L2_2_G1_MINI_ALU_OperationResult_8,
                   L1_1_L2_2_G1_MINI_ALU_OperationResult_7,
                   L1_1_L2_2_G1_MINI_ALU_OperationResult_6,
                   L1_1_L2_2_G1_MINI_ALU_OperationResult_5,
                   L1_1_L2_2_G1_MINI_ALU_OperationResult_4,
                   L1_1_L2_2_G1_MINI_ALU_OperationResult_3,
                   L1_1_L2_2_G1_MINI_ALU_OperationResult_2,
                   L1_1_L2_2_G1_MINI_ALU_OperationResult_1,
                   L1_1_L2_2_G1_MINI_ALU_OperationResult_0}), .BoothOperand ({
                   L1_1_L2_2_G1_MINI_ALU_BoothOperand_16,
                   L1_1_L2_2_G1_MINI_ALU_BoothOperand_15,
                   L1_1_L2_2_G1_MINI_ALU_BoothOperand_14,
                   L1_1_L2_2_G1_MINI_ALU_BoothOperand_13,
                   L1_1_L2_2_G1_MINI_ALU_BoothOperand_12,
                   L1_1_L2_2_G1_MINI_ALU_BoothOperand_11,
                   L1_1_L2_2_G1_MINI_ALU_BoothOperand_10,
                   L1_1_L2_2_G1_MINI_ALU_BoothOperand_9,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16}), .BoothP ({
                   L1_1_L2_2_G1_MINI_ALU_BoothP_16,
                   L1_1_L2_2_G1_MINI_ALU_BoothP_15,
                   L1_1_L2_2_G1_MINI_ALU_BoothP_14,
                   L1_1_L2_2_G1_MINI_ALU_BoothP_13,
                   L1_1_L2_2_G1_MINI_ALU_BoothP_12,
                   L1_1_L2_2_G1_MINI_ALU_BoothP_11,
                   L1_1_L2_2_G1_MINI_ALU_BoothP_10,
                   L1_1_L2_2_G1_MINI_ALU_BoothP_9,L1_1_L2_2_G1_MINI_ALU_BoothP_8
                   ,L1_1_L2_2_G1_MINI_ALU_BoothP_7,
                   L1_1_L2_2_G1_MINI_ALU_BoothP_6,L1_1_L2_2_G1_MINI_ALU_BoothP_5
                   ,L1_1_L2_2_G1_MINI_ALU_BoothP_4,
                   L1_1_L2_2_G1_MINI_ALU_BoothP_3,L1_1_L2_2_G1_MINI_ALU_BoothP_2
                   ,L1_1_L2_2_G1_MINI_ALU_BoothP_1,
                   L1_1_L2_2_G1_MINI_ALU_BoothP_0}), .SelOperand (nx3283), .Operation (
                   L1_1_L2_2_G1_MINI_ALU_BoothXORCheck), .AdderResult ({
                   L1ResultsLarge_7__16,L1ResultsLarge_7__15,
                   L1ResultsLarge_7__14,L1ResultsLarge_7__13,
                   L1ResultsLarge_7__12,L1ResultsLarge_7__11,
                   L1ResultsLarge_7__10,L1ResultsLarge_7__9,L1ResultsLarge_7__8,
                   L1ResultsLarge_7__7,L1ResultsLarge_7__6,L1ResultsLarge_7__5,
                   L1ResultsLarge_7__4,L1ResultsLarge_7__3,L1ResultsLarge_7__2,
                   L1ResultsLarge_7__1,L1ResultsLarge_7__0}), .AdderBoothResult (
                   {\$dummy [245],L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_15,
                   L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_14,
                   L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_13,
                   L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_12,
                   L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_11,
                   L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_10,
                   L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_9,
                   L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_8,
                   L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_7,
                   L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_6,
                   L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_5,
                   L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_4,
                   L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_3,
                   L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_2,
                   L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_1,
                   L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_0})) ;
    booth_unit_17 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT (.CLK (CLK), .RST (RST), .Start (
                  Start), .Instr (Instr), .LoopingAndResultNotReady (nx3277), .Filter (
                  {FilterDin_1__2__7,FilterDin_1__2__6,FilterDin_1__2__5,
                  FilterDin_1__2__4,FilterDin_1__2__3,FilterDin_1__2__2,
                  FilterDin_1__2__1,FilterDin_1__2__0}), .Window ({
                  WindowDin_1__2__7,WindowDin_1__2__6,WindowDin_1__2__5,
                  WindowDin_1__2__4,WindowDin_1__2__3,WindowDin_1__2__2,
                  WindowDin_1__2__1,WindowDin_1__2__0}), .AdderBoothResult ({
                  L1FirstOperands_12__16,
                  L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_15,
                  L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_14,
                  L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_13,
                  L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_12,
                  L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_11,
                  L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_10,
                  L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_9,
                  L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_8,
                  L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_7,
                  L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_6,
                  L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_5,
                  L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_4,
                  L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_3,
                  L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_2,
                  L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_1,
                  L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_0}), .BoothXORCheck (
                  L1_1_L2_2_G1_MINI_ALU_BoothXORCheck), .BoothResult ({
                  \$dummy [246],\$dummy [247],\$dummy [248],\$dummy [249],
                  \$dummy [250],\$dummy [251],\$dummy [252],\$dummy [253]}), .BoothAddingOperand (
                  {L1_1_L2_2_G1_MINI_ALU_BoothOperand_16,
                  L1_1_L2_2_G1_MINI_ALU_BoothOperand_15,
                  L1_1_L2_2_G1_MINI_ALU_BoothOperand_14,
                  L1_1_L2_2_G1_MINI_ALU_BoothOperand_13,
                  L1_1_L2_2_G1_MINI_ALU_BoothOperand_12,
                  L1_1_L2_2_G1_MINI_ALU_BoothOperand_11,
                  L1_1_L2_2_G1_MINI_ALU_BoothOperand_10,
                  L1_1_L2_2_G1_MINI_ALU_BoothOperand_9,\$dummy [254],
                  \$dummy [255],\$dummy [256],\$dummy [257],\$dummy [258],
                  \$dummy [259],\$dummy [260],\$dummy [261],\$dummy [262]}), .BoothP (
                  {L1_1_L2_2_G1_MINI_ALU_BoothP_16,
                  L1_1_L2_2_G1_MINI_ALU_BoothP_15,
                  L1_1_L2_2_G1_MINI_ALU_BoothP_14,
                  L1_1_L2_2_G1_MINI_ALU_BoothP_13,
                  L1_1_L2_2_G1_MINI_ALU_BoothP_12,
                  L1_1_L2_2_G1_MINI_ALU_BoothP_11,
                  L1_1_L2_2_G1_MINI_ALU_BoothP_10,L1_1_L2_2_G1_MINI_ALU_BoothP_9
                  ,L1_1_L2_2_G1_MINI_ALU_BoothP_8,L1_1_L2_2_G1_MINI_ALU_BoothP_7
                  ,L1_1_L2_2_G1_MINI_ALU_BoothP_6,L1_1_L2_2_G1_MINI_ALU_BoothP_5
                  ,L1_1_L2_2_G1_MINI_ALU_BoothP_4,L1_1_L2_2_G1_MINI_ALU_BoothP_3
                  ,L1_1_L2_2_G1_MINI_ALU_BoothP_2,L1_1_L2_2_G1_MINI_ALU_BoothP_1
                  ,L1_1_L2_2_G1_MINI_ALU_BoothP_0}), .LargeWindowShifted ({
                  \$dummy [263],\$dummy [264],\$dummy [265],\$dummy [266],
                  \$dummy [267],\$dummy [268],\$dummy [269],\$dummy [270],
                  \$dummy [271],\$dummy [272],\$dummy [273],\$dummy [274],
                  \$dummy [275],\$dummy [276],\$dummy [277],\$dummy [278],
                  \$dummy [279]})) ;
    booth_adder_17 L1_1_L2_3_G1_MINI_ALU_BOOTH_ADDER (.AdderFirstOperand ({
                   L1FirstOperands_12__16,L1FirstOperands_8__15,
                   L1FirstOperands_8__14,L1FirstOperands_8__13,
                   L1FirstOperands_8__12,L1FirstOperands_8__11,
                   L1FirstOperands_8__10,L1FirstOperands_8__9,
                   L1FirstOperands_8__8,L1FirstOperands_8__7,
                   L1FirstOperands_8__6,L1FirstOperands_8__5,
                   L1FirstOperands_8__4,L1FirstOperands_8__3,
                   L1FirstOperands_8__2,L1FirstOperands_8__1,
                   L1FirstOperands_8__0}), .AdderSecondOperand ({
                   L1FirstOperands_12__16,
                   L1_1_L2_3_G1_MINI_ALU_OperationResult_15,
                   L1_1_L2_3_G1_MINI_ALU_OperationResult_14,
                   L1_1_L2_3_G1_MINI_ALU_OperationResult_13,
                   L1_1_L2_3_G1_MINI_ALU_OperationResult_12,
                   L1_1_L2_3_G1_MINI_ALU_OperationResult_11,
                   L1_1_L2_3_G1_MINI_ALU_OperationResult_10,
                   L1_1_L2_3_G1_MINI_ALU_OperationResult_9,
                   L1_1_L2_3_G1_MINI_ALU_OperationResult_8,
                   L1_1_L2_3_G1_MINI_ALU_OperationResult_7,
                   L1_1_L2_3_G1_MINI_ALU_OperationResult_6,
                   L1_1_L2_3_G1_MINI_ALU_OperationResult_5,
                   L1_1_L2_3_G1_MINI_ALU_OperationResult_4,
                   L1_1_L2_3_G1_MINI_ALU_OperationResult_3,
                   L1_1_L2_3_G1_MINI_ALU_OperationResult_2,
                   L1_1_L2_3_G1_MINI_ALU_OperationResult_1,
                   L1_1_L2_3_G1_MINI_ALU_OperationResult_0}), .BoothOperand ({
                   L1_1_L2_3_G1_MINI_ALU_BoothOperand_16,
                   L1_1_L2_3_G1_MINI_ALU_BoothOperand_15,
                   L1_1_L2_3_G1_MINI_ALU_BoothOperand_14,
                   L1_1_L2_3_G1_MINI_ALU_BoothOperand_13,
                   L1_1_L2_3_G1_MINI_ALU_BoothOperand_12,
                   L1_1_L2_3_G1_MINI_ALU_BoothOperand_11,
                   L1_1_L2_3_G1_MINI_ALU_BoothOperand_10,
                   L1_1_L2_3_G1_MINI_ALU_BoothOperand_9,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16}), .BoothP ({
                   L1_1_L2_3_G1_MINI_ALU_BoothP_16,
                   L1_1_L2_3_G1_MINI_ALU_BoothP_15,
                   L1_1_L2_3_G1_MINI_ALU_BoothP_14,
                   L1_1_L2_3_G1_MINI_ALU_BoothP_13,
                   L1_1_L2_3_G1_MINI_ALU_BoothP_12,
                   L1_1_L2_3_G1_MINI_ALU_BoothP_11,
                   L1_1_L2_3_G1_MINI_ALU_BoothP_10,
                   L1_1_L2_3_G1_MINI_ALU_BoothP_9,L1_1_L2_3_G1_MINI_ALU_BoothP_8
                   ,L1_1_L2_3_G1_MINI_ALU_BoothP_7,
                   L1_1_L2_3_G1_MINI_ALU_BoothP_6,L1_1_L2_3_G1_MINI_ALU_BoothP_5
                   ,L1_1_L2_3_G1_MINI_ALU_BoothP_4,
                   L1_1_L2_3_G1_MINI_ALU_BoothP_3,L1_1_L2_3_G1_MINI_ALU_BoothP_2
                   ,L1_1_L2_3_G1_MINI_ALU_BoothP_1,
                   L1_1_L2_3_G1_MINI_ALU_BoothP_0}), .SelOperand (nx3285), .Operation (
                   L1_1_L2_3_G1_MINI_ALU_BoothXORCheck), .AdderResult ({
                   L1ResultsLarge_8__16,L1ResultsLarge_8__15,
                   L1ResultsLarge_8__14,L1ResultsLarge_8__13,
                   L1ResultsLarge_8__12,L1ResultsLarge_8__11,
                   L1ResultsLarge_8__10,L1ResultsLarge_8__9,L1ResultsLarge_8__8,
                   L1ResultsLarge_8__7,L1ResultsLarge_8__6,L1ResultsLarge_8__5,
                   L1ResultsLarge_8__4,L1ResultsLarge_8__3,L1ResultsLarge_8__2,
                   L1ResultsLarge_8__1,L1ResultsLarge_8__0}), .AdderBoothResult (
                   {\$dummy [280],L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_15,
                   L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_14,
                   L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_13,
                   L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_12,
                   L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_11,
                   L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_10,
                   L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_9,
                   L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_8,
                   L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_7,
                   L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_6,
                   L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_5,
                   L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_4,
                   L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_3,
                   L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_2,
                   L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_1,
                   L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_0})) ;
    booth_unit_17 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT (.CLK (CLK), .RST (RST), .Start (
                  Start), .Instr (Instr), .LoopingAndResultNotReady (nx3277), .Filter (
                  {FilterDin_1__3__7,FilterDin_1__3__6,FilterDin_1__3__5,
                  FilterDin_1__3__4,FilterDin_1__3__3,FilterDin_1__3__2,
                  FilterDin_1__3__1,FilterDin_1__3__0}), .Window ({
                  WindowDin_1__3__7,WindowDin_1__3__6,WindowDin_1__3__5,
                  WindowDin_1__3__4,WindowDin_1__3__3,WindowDin_1__3__2,
                  WindowDin_1__3__1,WindowDin_1__3__0}), .AdderBoothResult ({
                  L1FirstOperands_12__16,
                  L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_15,
                  L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_14,
                  L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_13,
                  L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_12,
                  L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_11,
                  L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_10,
                  L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_9,
                  L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_8,
                  L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_7,
                  L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_6,
                  L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_5,
                  L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_4,
                  L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_3,
                  L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_2,
                  L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_1,
                  L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_0}), .BoothXORCheck (
                  L1_1_L2_3_G1_MINI_ALU_BoothXORCheck), .BoothResult ({
                  \$dummy [281],\$dummy [282],\$dummy [283],\$dummy [284],
                  \$dummy [285],\$dummy [286],\$dummy [287],\$dummy [288]}), .BoothAddingOperand (
                  {L1_1_L2_3_G1_MINI_ALU_BoothOperand_16,
                  L1_1_L2_3_G1_MINI_ALU_BoothOperand_15,
                  L1_1_L2_3_G1_MINI_ALU_BoothOperand_14,
                  L1_1_L2_3_G1_MINI_ALU_BoothOperand_13,
                  L1_1_L2_3_G1_MINI_ALU_BoothOperand_12,
                  L1_1_L2_3_G1_MINI_ALU_BoothOperand_11,
                  L1_1_L2_3_G1_MINI_ALU_BoothOperand_10,
                  L1_1_L2_3_G1_MINI_ALU_BoothOperand_9,\$dummy [289],
                  \$dummy [290],\$dummy [291],\$dummy [292],\$dummy [293],
                  \$dummy [294],\$dummy [295],\$dummy [296],\$dummy [297]}), .BoothP (
                  {L1_1_L2_3_G1_MINI_ALU_BoothP_16,
                  L1_1_L2_3_G1_MINI_ALU_BoothP_15,
                  L1_1_L2_3_G1_MINI_ALU_BoothP_14,
                  L1_1_L2_3_G1_MINI_ALU_BoothP_13,
                  L1_1_L2_3_G1_MINI_ALU_BoothP_12,
                  L1_1_L2_3_G1_MINI_ALU_BoothP_11,
                  L1_1_L2_3_G1_MINI_ALU_BoothP_10,L1_1_L2_3_G1_MINI_ALU_BoothP_9
                  ,L1_1_L2_3_G1_MINI_ALU_BoothP_8,L1_1_L2_3_G1_MINI_ALU_BoothP_7
                  ,L1_1_L2_3_G1_MINI_ALU_BoothP_6,L1_1_L2_3_G1_MINI_ALU_BoothP_5
                  ,L1_1_L2_3_G1_MINI_ALU_BoothP_4,L1_1_L2_3_G1_MINI_ALU_BoothP_3
                  ,L1_1_L2_3_G1_MINI_ALU_BoothP_2,L1_1_L2_3_G1_MINI_ALU_BoothP_1
                  ,L1_1_L2_3_G1_MINI_ALU_BoothP_0}), .LargeWindowShifted ({
                  \$dummy [298],\$dummy [299],\$dummy [300],\$dummy [301],
                  \$dummy [302],\$dummy [303],\$dummy [304],\$dummy [305],
                  \$dummy [306],\$dummy [307],\$dummy [308],\$dummy [309],
                  \$dummy [310],\$dummy [311],\$dummy [312],\$dummy [313],
                  \$dummy [314]})) ;
    booth_adder_17 L1_1_L2_4_G1_MINI_ALU_BOOTH_ADDER (.AdderFirstOperand ({
                   L1FirstOperands_12__16,L1FirstOperands_4__15,
                   L1FirstOperands_4__14,L1FirstOperands_4__13,
                   L1FirstOperands_4__12,L1FirstOperands_4__11,
                   L1FirstOperands_4__10,L1FirstOperands_4__9,
                   L1FirstOperands_4__8,L1FirstOperands_4__7,
                   L1FirstOperands_4__6,L1FirstOperands_4__5,
                   L1FirstOperands_4__4,L1FirstOperands_4__3,
                   L1FirstOperands_4__2,L1FirstOperands_4__1,
                   L1FirstOperands_4__0}), .AdderSecondOperand ({
                   L1FirstOperands_12__16,
                   L1_1_L2_4_G1_MINI_ALU_OperationResult_15,
                   L1_1_L2_4_G1_MINI_ALU_OperationResult_14,
                   L1_1_L2_4_G1_MINI_ALU_OperationResult_13,
                   L1_1_L2_4_G1_MINI_ALU_OperationResult_12,
                   L1_1_L2_4_G1_MINI_ALU_OperationResult_11,
                   L1_1_L2_4_G1_MINI_ALU_OperationResult_10,
                   L1_1_L2_4_G1_MINI_ALU_OperationResult_9,
                   L1_1_L2_4_G1_MINI_ALU_OperationResult_8,
                   L1_1_L2_4_G1_MINI_ALU_OperationResult_7,
                   L1_1_L2_4_G1_MINI_ALU_OperationResult_6,
                   L1_1_L2_4_G1_MINI_ALU_OperationResult_5,
                   L1_1_L2_4_G1_MINI_ALU_OperationResult_4,
                   L1_1_L2_4_G1_MINI_ALU_OperationResult_3,
                   L1_1_L2_4_G1_MINI_ALU_OperationResult_2,
                   L1_1_L2_4_G1_MINI_ALU_OperationResult_1,
                   L1_1_L2_4_G1_MINI_ALU_OperationResult_0}), .BoothOperand ({
                   L1_1_L2_4_G1_MINI_ALU_BoothOperand_16,
                   L1_1_L2_4_G1_MINI_ALU_BoothOperand_15,
                   L1_1_L2_4_G1_MINI_ALU_BoothOperand_14,
                   L1_1_L2_4_G1_MINI_ALU_BoothOperand_13,
                   L1_1_L2_4_G1_MINI_ALU_BoothOperand_12,
                   L1_1_L2_4_G1_MINI_ALU_BoothOperand_11,
                   L1_1_L2_4_G1_MINI_ALU_BoothOperand_10,
                   L1_1_L2_4_G1_MINI_ALU_BoothOperand_9,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16}), .BoothP ({
                   L1_1_L2_4_G1_MINI_ALU_BoothP_16,
                   L1_1_L2_4_G1_MINI_ALU_BoothP_15,
                   L1_1_L2_4_G1_MINI_ALU_BoothP_14,
                   L1_1_L2_4_G1_MINI_ALU_BoothP_13,
                   L1_1_L2_4_G1_MINI_ALU_BoothP_12,
                   L1_1_L2_4_G1_MINI_ALU_BoothP_11,
                   L1_1_L2_4_G1_MINI_ALU_BoothP_10,
                   L1_1_L2_4_G1_MINI_ALU_BoothP_9,L1_1_L2_4_G1_MINI_ALU_BoothP_8
                   ,L1_1_L2_4_G1_MINI_ALU_BoothP_7,
                   L1_1_L2_4_G1_MINI_ALU_BoothP_6,L1_1_L2_4_G1_MINI_ALU_BoothP_5
                   ,L1_1_L2_4_G1_MINI_ALU_BoothP_4,
                   L1_1_L2_4_G1_MINI_ALU_BoothP_3,L1_1_L2_4_G1_MINI_ALU_BoothP_2
                   ,L1_1_L2_4_G1_MINI_ALU_BoothP_1,
                   L1_1_L2_4_G1_MINI_ALU_BoothP_0}), .SelOperand (nx3285), .Operation (
                   L1_1_L2_4_G1_MINI_ALU_BoothXORCheck), .AdderResult ({
                   L1ResultsLarge_9__16,L1ResultsLarge_9__15,
                   L1ResultsLarge_9__14,L1ResultsLarge_9__13,
                   L1ResultsLarge_9__12,L1ResultsLarge_9__11,
                   L1ResultsLarge_9__10,L1ResultsLarge_9__9,L1ResultsLarge_9__8,
                   L1ResultsLarge_9__7,L1ResultsLarge_9__6,L1ResultsLarge_9__5,
                   L1ResultsLarge_9__4,L1ResultsLarge_9__3,L1ResultsLarge_9__2,
                   L1ResultsLarge_9__1,L1ResultsLarge_9__0}), .AdderBoothResult (
                   {\$dummy [315],L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_15,
                   L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_14,
                   L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_13,
                   L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_12,
                   L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_11,
                   L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_10,
                   L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_9,
                   L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_8,
                   L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_7,
                   L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_6,
                   L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_5,
                   L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_4,
                   L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_3,
                   L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_2,
                   L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_1,
                   L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_0})) ;
    booth_unit_17 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT (.CLK (CLK), .RST (RST), .Start (
                  Start), .Instr (Instr), .LoopingAndResultNotReady (nx3277), .Filter (
                  {FilterDin_1__4__7,FilterDin_1__4__6,FilterDin_1__4__5,
                  FilterDin_1__4__4,FilterDin_1__4__3,FilterDin_1__4__2,
                  FilterDin_1__4__1,FilterDin_1__4__0}), .Window ({
                  WindowDin_1__4__7,WindowDin_1__4__6,WindowDin_1__4__5,
                  WindowDin_1__4__4,WindowDin_1__4__3,WindowDin_1__4__2,
                  WindowDin_1__4__1,WindowDin_1__4__0}), .AdderBoothResult ({
                  L1FirstOperands_12__16,
                  L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_15,
                  L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_14,
                  L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_13,
                  L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_12,
                  L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_11,
                  L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_10,
                  L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_9,
                  L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_8,
                  L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_7,
                  L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_6,
                  L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_5,
                  L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_4,
                  L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_3,
                  L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_2,
                  L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_1,
                  L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_0}), .BoothXORCheck (
                  L1_1_L2_4_G1_MINI_ALU_BoothXORCheck), .BoothResult ({
                  \$dummy [316],\$dummy [317],\$dummy [318],\$dummy [319],
                  \$dummy [320],\$dummy [321],\$dummy [322],\$dummy [323]}), .BoothAddingOperand (
                  {L1_1_L2_4_G1_MINI_ALU_BoothOperand_16,
                  L1_1_L2_4_G1_MINI_ALU_BoothOperand_15,
                  L1_1_L2_4_G1_MINI_ALU_BoothOperand_14,
                  L1_1_L2_4_G1_MINI_ALU_BoothOperand_13,
                  L1_1_L2_4_G1_MINI_ALU_BoothOperand_12,
                  L1_1_L2_4_G1_MINI_ALU_BoothOperand_11,
                  L1_1_L2_4_G1_MINI_ALU_BoothOperand_10,
                  L1_1_L2_4_G1_MINI_ALU_BoothOperand_9,\$dummy [324],
                  \$dummy [325],\$dummy [326],\$dummy [327],\$dummy [328],
                  \$dummy [329],\$dummy [330],\$dummy [331],\$dummy [332]}), .BoothP (
                  {L1_1_L2_4_G1_MINI_ALU_BoothP_16,
                  L1_1_L2_4_G1_MINI_ALU_BoothP_15,
                  L1_1_L2_4_G1_MINI_ALU_BoothP_14,
                  L1_1_L2_4_G1_MINI_ALU_BoothP_13,
                  L1_1_L2_4_G1_MINI_ALU_BoothP_12,
                  L1_1_L2_4_G1_MINI_ALU_BoothP_11,
                  L1_1_L2_4_G1_MINI_ALU_BoothP_10,L1_1_L2_4_G1_MINI_ALU_BoothP_9
                  ,L1_1_L2_4_G1_MINI_ALU_BoothP_8,L1_1_L2_4_G1_MINI_ALU_BoothP_7
                  ,L1_1_L2_4_G1_MINI_ALU_BoothP_6,L1_1_L2_4_G1_MINI_ALU_BoothP_5
                  ,L1_1_L2_4_G1_MINI_ALU_BoothP_4,L1_1_L2_4_G1_MINI_ALU_BoothP_3
                  ,L1_1_L2_4_G1_MINI_ALU_BoothP_2,L1_1_L2_4_G1_MINI_ALU_BoothP_1
                  ,L1_1_L2_4_G1_MINI_ALU_BoothP_0}), .LargeWindowShifted ({
                  \$dummy [333],\$dummy [334],\$dummy [335],\$dummy [336],
                  \$dummy [337],\$dummy [338],\$dummy [339],\$dummy [340],
                  \$dummy [341],\$dummy [342],\$dummy [343],\$dummy [344],
                  \$dummy [345],\$dummy [346],\$dummy [347],\$dummy [348],
                  \$dummy [349]})) ;
    booth_adder_17 L1_2_L2_0_G1_MINI_ALU_BOOTH_ADDER (.AdderFirstOperand ({
                   L1FirstOperands_12__16,L1FirstOperands_10__15,
                   L1FirstOperands_10__14,L1FirstOperands_10__13,
                   L1FirstOperands_10__12,L1FirstOperands_10__11,
                   L1FirstOperands_10__10,L1FirstOperands_10__9,
                   L1FirstOperands_10__8,L1FirstOperands_10__7,
                   L1FirstOperands_10__6,L1FirstOperands_10__5,
                   L1FirstOperands_10__4,L1FirstOperands_10__3,
                   L1FirstOperands_10__2,L1FirstOperands_10__1,
                   L1FirstOperands_10__0}), .AdderSecondOperand ({
                   L1FirstOperands_12__16,
                   L1_2_L2_0_G1_MINI_ALU_OperationResult_15,
                   L1_2_L2_0_G1_MINI_ALU_OperationResult_14,
                   L1_2_L2_0_G1_MINI_ALU_OperationResult_13,
                   L1_2_L2_0_G1_MINI_ALU_OperationResult_12,
                   L1_2_L2_0_G1_MINI_ALU_OperationResult_11,
                   L1_2_L2_0_G1_MINI_ALU_OperationResult_10,
                   L1_2_L2_0_G1_MINI_ALU_OperationResult_9,
                   L1_2_L2_0_G1_MINI_ALU_OperationResult_8,
                   L1_2_L2_0_G1_MINI_ALU_OperationResult_7,
                   L1_2_L2_0_G1_MINI_ALU_OperationResult_6,
                   L1_2_L2_0_G1_MINI_ALU_OperationResult_5,
                   L1_2_L2_0_G1_MINI_ALU_OperationResult_4,
                   L1_2_L2_0_G1_MINI_ALU_OperationResult_3,
                   L1_2_L2_0_G1_MINI_ALU_OperationResult_2,
                   L1_2_L2_0_G1_MINI_ALU_OperationResult_1,
                   L1_2_L2_0_G1_MINI_ALU_OperationResult_0}), .BoothOperand ({
                   L1_2_L2_0_G1_MINI_ALU_BoothOperand_16,
                   L1_2_L2_0_G1_MINI_ALU_BoothOperand_15,
                   L1_2_L2_0_G1_MINI_ALU_BoothOperand_14,
                   L1_2_L2_0_G1_MINI_ALU_BoothOperand_13,
                   L1_2_L2_0_G1_MINI_ALU_BoothOperand_12,
                   L1_2_L2_0_G1_MINI_ALU_BoothOperand_11,
                   L1_2_L2_0_G1_MINI_ALU_BoothOperand_10,
                   L1_2_L2_0_G1_MINI_ALU_BoothOperand_9,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16}), .BoothP ({
                   L1_2_L2_0_G1_MINI_ALU_BoothP_16,
                   L1_2_L2_0_G1_MINI_ALU_BoothP_15,
                   L1_2_L2_0_G1_MINI_ALU_BoothP_14,
                   L1_2_L2_0_G1_MINI_ALU_BoothP_13,
                   L1_2_L2_0_G1_MINI_ALU_BoothP_12,
                   L1_2_L2_0_G1_MINI_ALU_BoothP_11,
                   L1_2_L2_0_G1_MINI_ALU_BoothP_10,
                   L1_2_L2_0_G1_MINI_ALU_BoothP_9,L1_2_L2_0_G1_MINI_ALU_BoothP_8
                   ,L1_2_L2_0_G1_MINI_ALU_BoothP_7,
                   L1_2_L2_0_G1_MINI_ALU_BoothP_6,L1_2_L2_0_G1_MINI_ALU_BoothP_5
                   ,L1_2_L2_0_G1_MINI_ALU_BoothP_4,
                   L1_2_L2_0_G1_MINI_ALU_BoothP_3,L1_2_L2_0_G1_MINI_ALU_BoothP_2
                   ,L1_2_L2_0_G1_MINI_ALU_BoothP_1,
                   L1_2_L2_0_G1_MINI_ALU_BoothP_0}), .SelOperand (nx3285), .Operation (
                   L1_2_L2_0_G1_MINI_ALU_BoothXORCheck), .AdderResult ({
                   L1ResultsLarge_10__16,L1ResultsLarge_10__15,
                   L1ResultsLarge_10__14,L1ResultsLarge_10__13,
                   L1ResultsLarge_10__12,L1ResultsLarge_10__11,
                   L1ResultsLarge_10__10,L1ResultsLarge_10__9,
                   L1ResultsLarge_10__8,L1ResultsLarge_10__7,
                   L1ResultsLarge_10__6,L1ResultsLarge_10__5,
                   L1ResultsLarge_10__4,L1ResultsLarge_10__3,
                   L1ResultsLarge_10__2,L1ResultsLarge_10__1,
                   L1ResultsLarge_10__0}), .AdderBoothResult ({\$dummy [350],
                   L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_15,
                   L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_14,
                   L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_13,
                   L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_12,
                   L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_11,
                   L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_10,
                   L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_9,
                   L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_8,
                   L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_7,
                   L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_6,
                   L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_5,
                   L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_4,
                   L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_3,
                   L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_2,
                   L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_1,
                   L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_0})) ;
    booth_unit_17 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT (.CLK (CLK), .RST (RST), .Start (
                  Start), .Instr (Instr), .LoopingAndResultNotReady (nx3277), .Filter (
                  {FilterDin_2__0__7,FilterDin_2__0__6,FilterDin_2__0__5,
                  FilterDin_2__0__4,FilterDin_2__0__3,FilterDin_2__0__2,
                  FilterDin_2__0__1,FilterDin_2__0__0}), .Window ({
                  WindowDin_2__0__7,WindowDin_2__0__6,WindowDin_2__0__5,
                  WindowDin_2__0__4,WindowDin_2__0__3,WindowDin_2__0__2,
                  WindowDin_2__0__1,WindowDin_2__0__0}), .AdderBoothResult ({
                  L1FirstOperands_12__16,
                  L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_15,
                  L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_14,
                  L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_13,
                  L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_12,
                  L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_11,
                  L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_10,
                  L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_9,
                  L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_8,
                  L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_7,
                  L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_6,
                  L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_5,
                  L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_4,
                  L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_3,
                  L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_2,
                  L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_1,
                  L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_0}), .BoothXORCheck (
                  L1_2_L2_0_G1_MINI_ALU_BoothXORCheck), .BoothResult ({
                  \$dummy [351],\$dummy [352],\$dummy [353],\$dummy [354],
                  \$dummy [355],\$dummy [356],\$dummy [357],\$dummy [358]}), .BoothAddingOperand (
                  {L1_2_L2_0_G1_MINI_ALU_BoothOperand_16,
                  L1_2_L2_0_G1_MINI_ALU_BoothOperand_15,
                  L1_2_L2_0_G1_MINI_ALU_BoothOperand_14,
                  L1_2_L2_0_G1_MINI_ALU_BoothOperand_13,
                  L1_2_L2_0_G1_MINI_ALU_BoothOperand_12,
                  L1_2_L2_0_G1_MINI_ALU_BoothOperand_11,
                  L1_2_L2_0_G1_MINI_ALU_BoothOperand_10,
                  L1_2_L2_0_G1_MINI_ALU_BoothOperand_9,\$dummy [359],
                  \$dummy [360],\$dummy [361],\$dummy [362],\$dummy [363],
                  \$dummy [364],\$dummy [365],\$dummy [366],\$dummy [367]}), .BoothP (
                  {L1_2_L2_0_G1_MINI_ALU_BoothP_16,
                  L1_2_L2_0_G1_MINI_ALU_BoothP_15,
                  L1_2_L2_0_G1_MINI_ALU_BoothP_14,
                  L1_2_L2_0_G1_MINI_ALU_BoothP_13,
                  L1_2_L2_0_G1_MINI_ALU_BoothP_12,
                  L1_2_L2_0_G1_MINI_ALU_BoothP_11,
                  L1_2_L2_0_G1_MINI_ALU_BoothP_10,L1_2_L2_0_G1_MINI_ALU_BoothP_9
                  ,L1_2_L2_0_G1_MINI_ALU_BoothP_8,L1_2_L2_0_G1_MINI_ALU_BoothP_7
                  ,L1_2_L2_0_G1_MINI_ALU_BoothP_6,L1_2_L2_0_G1_MINI_ALU_BoothP_5
                  ,L1_2_L2_0_G1_MINI_ALU_BoothP_4,L1_2_L2_0_G1_MINI_ALU_BoothP_3
                  ,L1_2_L2_0_G1_MINI_ALU_BoothP_2,L1_2_L2_0_G1_MINI_ALU_BoothP_1
                  ,L1_2_L2_0_G1_MINI_ALU_BoothP_0}), .LargeWindowShifted ({
                  \$dummy [368],\$dummy [369],\$dummy [370],\$dummy [371],
                  \$dummy [372],\$dummy [373],\$dummy [374],\$dummy [375],
                  \$dummy [376],\$dummy [377],\$dummy [378],\$dummy [379],
                  \$dummy [380],\$dummy [381],\$dummy [382],\$dummy [383],
                  \$dummy [384]})) ;
    booth_adder_17 L1_2_L2_1_G1_MINI_ALU_BOOTH_ADDER (.AdderFirstOperand ({
                   L1FirstOperands_12__16,L1FirstOperands_11__15,
                   L1FirstOperands_11__14,L1FirstOperands_11__13,
                   L1FirstOperands_11__12,L1FirstOperands_11__11,
                   L1FirstOperands_11__10,L1FirstOperands_11__9,
                   L1FirstOperands_11__8,L1FirstOperands_11__7,
                   L1FirstOperands_11__6,L1FirstOperands_11__5,
                   L1FirstOperands_11__4,L1FirstOperands_11__3,
                   L1FirstOperands_11__2,L1FirstOperands_11__1,
                   L1FirstOperands_11__0}), .AdderSecondOperand ({
                   L1FirstOperands_12__16,
                   L1_2_L2_1_G1_MINI_ALU_OperationResult_15,
                   L1_2_L2_1_G1_MINI_ALU_OperationResult_14,
                   L1_2_L2_1_G1_MINI_ALU_OperationResult_13,
                   L1_2_L2_1_G1_MINI_ALU_OperationResult_12,
                   L1_2_L2_1_G1_MINI_ALU_OperationResult_11,
                   L1_2_L2_1_G1_MINI_ALU_OperationResult_10,
                   L1_2_L2_1_G1_MINI_ALU_OperationResult_9,
                   L1_2_L2_1_G1_MINI_ALU_OperationResult_8,
                   L1_2_L2_1_G1_MINI_ALU_OperationResult_7,
                   L1_2_L2_1_G1_MINI_ALU_OperationResult_6,
                   L1_2_L2_1_G1_MINI_ALU_OperationResult_5,
                   L1_2_L2_1_G1_MINI_ALU_OperationResult_4,
                   L1_2_L2_1_G1_MINI_ALU_OperationResult_3,
                   L1_2_L2_1_G1_MINI_ALU_OperationResult_2,
                   L1_2_L2_1_G1_MINI_ALU_OperationResult_1,
                   L1_2_L2_1_G1_MINI_ALU_OperationResult_0}), .BoothOperand ({
                   L1_2_L2_1_G1_MINI_ALU_BoothOperand_16,
                   L1_2_L2_1_G1_MINI_ALU_BoothOperand_15,
                   L1_2_L2_1_G1_MINI_ALU_BoothOperand_14,
                   L1_2_L2_1_G1_MINI_ALU_BoothOperand_13,
                   L1_2_L2_1_G1_MINI_ALU_BoothOperand_12,
                   L1_2_L2_1_G1_MINI_ALU_BoothOperand_11,
                   L1_2_L2_1_G1_MINI_ALU_BoothOperand_10,
                   L1_2_L2_1_G1_MINI_ALU_BoothOperand_9,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16}), .BoothP ({
                   L1_2_L2_1_G1_MINI_ALU_BoothP_16,
                   L1_2_L2_1_G1_MINI_ALU_BoothP_15,
                   L1_2_L2_1_G1_MINI_ALU_BoothP_14,
                   L1_2_L2_1_G1_MINI_ALU_BoothP_13,
                   L1_2_L2_1_G1_MINI_ALU_BoothP_12,
                   L1_2_L2_1_G1_MINI_ALU_BoothP_11,
                   L1_2_L2_1_G1_MINI_ALU_BoothP_10,
                   L1_2_L2_1_G1_MINI_ALU_BoothP_9,L1_2_L2_1_G1_MINI_ALU_BoothP_8
                   ,L1_2_L2_1_G1_MINI_ALU_BoothP_7,
                   L1_2_L2_1_G1_MINI_ALU_BoothP_6,L1_2_L2_1_G1_MINI_ALU_BoothP_5
                   ,L1_2_L2_1_G1_MINI_ALU_BoothP_4,
                   L1_2_L2_1_G1_MINI_ALU_BoothP_3,L1_2_L2_1_G1_MINI_ALU_BoothP_2
                   ,L1_2_L2_1_G1_MINI_ALU_BoothP_1,
                   L1_2_L2_1_G1_MINI_ALU_BoothP_0}), .SelOperand (nx3285), .Operation (
                   L1_2_L2_1_G1_MINI_ALU_BoothXORCheck), .AdderResult ({
                   L1ResultsLarge_11__16,L1ResultsLarge_11__15,
                   L1ResultsLarge_11__14,L1ResultsLarge_11__13,
                   L1ResultsLarge_11__12,L1ResultsLarge_11__11,
                   L1ResultsLarge_11__10,L1ResultsLarge_11__9,
                   L1ResultsLarge_11__8,L1ResultsLarge_11__7,
                   L1ResultsLarge_11__6,L1ResultsLarge_11__5,
                   L1ResultsLarge_11__4,L1ResultsLarge_11__3,
                   L1ResultsLarge_11__2,L1ResultsLarge_11__1,
                   L1ResultsLarge_11__0}), .AdderBoothResult ({\$dummy [385],
                   L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_15,
                   L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_14,
                   L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_13,
                   L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_12,
                   L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_11,
                   L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_10,
                   L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_9,
                   L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_8,
                   L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_7,
                   L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_6,
                   L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_5,
                   L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_4,
                   L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_3,
                   L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_2,
                   L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_1,
                   L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_0})) ;
    booth_unit_17 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT (.CLK (CLK), .RST (RST), .Start (
                  Start), .Instr (Instr), .LoopingAndResultNotReady (nx3277), .Filter (
                  {FilterDin_2__1__7,FilterDin_2__1__6,FilterDin_2__1__5,
                  FilterDin_2__1__4,FilterDin_2__1__3,FilterDin_2__1__2,
                  FilterDin_2__1__1,FilterDin_2__1__0}), .Window ({
                  WindowDin_2__1__7,WindowDin_2__1__6,WindowDin_2__1__5,
                  WindowDin_2__1__4,WindowDin_2__1__3,WindowDin_2__1__2,
                  WindowDin_2__1__1,WindowDin_2__1__0}), .AdderBoothResult ({
                  L1FirstOperands_12__16,
                  L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_15,
                  L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_14,
                  L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_13,
                  L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_12,
                  L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_11,
                  L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_10,
                  L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_9,
                  L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_8,
                  L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_7,
                  L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_6,
                  L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_5,
                  L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_4,
                  L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_3,
                  L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_2,
                  L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_1,
                  L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_0}), .BoothXORCheck (
                  L1_2_L2_1_G1_MINI_ALU_BoothXORCheck), .BoothResult ({
                  \$dummy [386],\$dummy [387],\$dummy [388],\$dummy [389],
                  \$dummy [390],\$dummy [391],\$dummy [392],\$dummy [393]}), .BoothAddingOperand (
                  {L1_2_L2_1_G1_MINI_ALU_BoothOperand_16,
                  L1_2_L2_1_G1_MINI_ALU_BoothOperand_15,
                  L1_2_L2_1_G1_MINI_ALU_BoothOperand_14,
                  L1_2_L2_1_G1_MINI_ALU_BoothOperand_13,
                  L1_2_L2_1_G1_MINI_ALU_BoothOperand_12,
                  L1_2_L2_1_G1_MINI_ALU_BoothOperand_11,
                  L1_2_L2_1_G1_MINI_ALU_BoothOperand_10,
                  L1_2_L2_1_G1_MINI_ALU_BoothOperand_9,\$dummy [394],
                  \$dummy [395],\$dummy [396],\$dummy [397],\$dummy [398],
                  \$dummy [399],\$dummy [400],\$dummy [401],\$dummy [402]}), .BoothP (
                  {L1_2_L2_1_G1_MINI_ALU_BoothP_16,
                  L1_2_L2_1_G1_MINI_ALU_BoothP_15,
                  L1_2_L2_1_G1_MINI_ALU_BoothP_14,
                  L1_2_L2_1_G1_MINI_ALU_BoothP_13,
                  L1_2_L2_1_G1_MINI_ALU_BoothP_12,
                  L1_2_L2_1_G1_MINI_ALU_BoothP_11,
                  L1_2_L2_1_G1_MINI_ALU_BoothP_10,L1_2_L2_1_G1_MINI_ALU_BoothP_9
                  ,L1_2_L2_1_G1_MINI_ALU_BoothP_8,L1_2_L2_1_G1_MINI_ALU_BoothP_7
                  ,L1_2_L2_1_G1_MINI_ALU_BoothP_6,L1_2_L2_1_G1_MINI_ALU_BoothP_5
                  ,L1_2_L2_1_G1_MINI_ALU_BoothP_4,L1_2_L2_1_G1_MINI_ALU_BoothP_3
                  ,L1_2_L2_1_G1_MINI_ALU_BoothP_2,L1_2_L2_1_G1_MINI_ALU_BoothP_1
                  ,L1_2_L2_1_G1_MINI_ALU_BoothP_0}), .LargeWindowShifted ({
                  \$dummy [403],\$dummy [404],\$dummy [405],\$dummy [406],
                  \$dummy [407],\$dummy [408],\$dummy [409],\$dummy [410],
                  \$dummy [411],\$dummy [412],\$dummy [413],\$dummy [414],
                  \$dummy [415],\$dummy [416],\$dummy [417],\$dummy [418],
                  \$dummy [419]})) ;
    booth_adder_17_unfolded3 L1_2_L2_2_G1_MINI_ALU_BOOTH_ADDER (.AdderFirstOperand (
                             {L1FirstOperands_12__16,L1FirstOperands_12__16,
                             L1FirstOperands_12__16,L1FirstOperands_12__16,
                             L1FirstOperands_12__16,L1FirstOperands_12__16,
                             L1FirstOperands_12__16,L1FirstOperands_12__16,
                             L1FirstOperands_12__16,L1FirstOperands_12__16,
                             L1FirstOperands_12__16,L1FirstOperands_12__16,
                             L1FirstOperands_12__16,L1FirstOperands_12__16,
                             L1FirstOperands_12__16,L1FirstOperands_12__16,
                             L1FirstOperands_12__16}), .AdderSecondOperand ({
                             L1FirstOperands_12__16,L1FirstOperands_12__16,
                             L1FirstOperands_12__16,L1FirstOperands_12__16,
                             L1FirstOperands_12__16,L1FirstOperands_12__16,
                             L1FirstOperands_12__16,L1FirstOperands_12__16,
                             L1FirstOperands_12__16,L1FirstOperands_12__16,
                             L1FirstOperands_12__16,L1FirstOperands_12__16,
                             L1FirstOperands_12__16,L1FirstOperands_12__16,
                             L1FirstOperands_12__16,L1FirstOperands_12__16,
                             L1FirstOperands_12__16}), .BoothOperand ({
                             L1_2_L2_2_G1_MINI_ALU_BoothOperand_16,
                             L1_2_L2_2_G1_MINI_ALU_BoothOperand_15,
                             L1_2_L2_2_G1_MINI_ALU_BoothOperand_14,
                             L1_2_L2_2_G1_MINI_ALU_BoothOperand_13,
                             L1_2_L2_2_G1_MINI_ALU_BoothOperand_12,
                             L1_2_L2_2_G1_MINI_ALU_BoothOperand_11,
                             L1_2_L2_2_G1_MINI_ALU_BoothOperand_10,
                             L1_2_L2_2_G1_MINI_ALU_BoothOperand_9,
                             L1FirstOperands_12__16,L1FirstOperands_12__16,
                             L1FirstOperands_12__16,L1FirstOperands_12__16,
                             L1FirstOperands_12__16,L1FirstOperands_12__16,
                             L1FirstOperands_12__16,L1FirstOperands_12__16,
                             L1FirstOperands_12__16}), .BoothP ({
                             L1_2_L2_2_G1_MINI_ALU_BoothP_16,
                             L1_2_L2_2_G1_MINI_ALU_BoothP_15,
                             L1_2_L2_2_G1_MINI_ALU_BoothP_14,
                             L1_2_L2_2_G1_MINI_ALU_BoothP_13,
                             L1_2_L2_2_G1_MINI_ALU_BoothP_12,
                             L1_2_L2_2_G1_MINI_ALU_BoothP_11,
                             L1_2_L2_2_G1_MINI_ALU_BoothP_10,
                             L1_2_L2_2_G1_MINI_ALU_BoothP_9,
                             L1_2_L2_2_G1_MINI_ALU_BoothP_8,
                             L1_2_L2_2_G1_MINI_ALU_BoothP_7,
                             L1_2_L2_2_G1_MINI_ALU_BoothP_6,
                             L1_2_L2_2_G1_MINI_ALU_BoothP_5,
                             L1_2_L2_2_G1_MINI_ALU_BoothP_4,
                             L1_2_L2_2_G1_MINI_ALU_BoothP_3,
                             L1_2_L2_2_G1_MINI_ALU_BoothP_2,
                             L1_2_L2_2_G1_MINI_ALU_BoothP_1,
                             L1FirstOperands_12__16}), .SelOperand (nx3283), .Operation (
                             L1_2_L2_2_G1_MINI_ALU_BoothXORCheck), .AdderResult (
                             {\$dummy [420],\$dummy [421],\$dummy [422],
                             \$dummy [423],\$dummy [424],\$dummy [425],
                             \$dummy [426],\$dummy [427],\$dummy [428],
                             \$dummy [429],\$dummy [430],\$dummy [431],
                             \$dummy [432],\$dummy [433],\$dummy [434],
                             \$dummy [435],\$dummy [436]}), .AdderBoothResult ({
                             \$dummy [437],
                             L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_15,
                             L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_14,
                             L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_13,
                             L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_12,
                             L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_11,
                             L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_10,
                             L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_9,
                             L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_8,
                             L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_7,
                             L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_6,
                             L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_5,
                             L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_4,
                             L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_3,
                             L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_2,
                             L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_1,
                             L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_0})) ;
    booth_unit_17_unfolded1 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT (.CLK (CLK), .RST (
                            RST), .Start (Start), .Instr (Instr), .LoopingAndResultNotReady (
                            nx3277), .Filter ({FilterDin_2__2__7,
                            FilterDin_2__2__6,FilterDin_2__2__5,
                            FilterDin_2__2__4,FilterDin_2__2__3,
                            FilterDin_2__2__2,FilterDin_2__2__1,
                            FilterDin_2__2__0}), .Window ({WindowDin_2__2__7,
                            WindowDin_2__2__6,WindowDin_2__2__5,
                            WindowDin_2__2__4,WindowDin_2__2__3,
                            WindowDin_2__2__2,WindowDin_2__2__1,
                            WindowDin_2__2__0}), .AdderBoothResult ({
                            L1FirstOperands_12__16,
                            L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_15,
                            L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_14,
                            L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_13,
                            L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_12,
                            L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_11,
                            L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_10,
                            L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_9,
                            L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_8,
                            L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_7,
                            L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_6,
                            L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_5,
                            L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_4,
                            L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_3,
                            L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_2,
                            L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_1,
                            L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_0}), .BoothXORCheck (
                            L1_2_L2_2_G1_MINI_ALU_BoothXORCheck), .BoothResult (
                            {\$dummy [438],\$dummy [439],\$dummy [440],
                            \$dummy [441],\$dummy [442],\$dummy [443],
                            \$dummy [444],\$dummy [445]}), .BoothAddingOperand (
                            {L1_2_L2_2_G1_MINI_ALU_BoothOperand_16,
                            L1_2_L2_2_G1_MINI_ALU_BoothOperand_15,
                            L1_2_L2_2_G1_MINI_ALU_BoothOperand_14,
                            L1_2_L2_2_G1_MINI_ALU_BoothOperand_13,
                            L1_2_L2_2_G1_MINI_ALU_BoothOperand_12,
                            L1_2_L2_2_G1_MINI_ALU_BoothOperand_11,
                            L1_2_L2_2_G1_MINI_ALU_BoothOperand_10,
                            L1_2_L2_2_G1_MINI_ALU_BoothOperand_9,\$dummy [446],
                            \$dummy [447],\$dummy [448],\$dummy [449],
                            \$dummy [450],\$dummy [451],\$dummy [452],
                            \$dummy [453],\$dummy [454]}), .BoothP ({
                            L1_2_L2_2_G1_MINI_ALU_BoothP_16,
                            L1_2_L2_2_G1_MINI_ALU_BoothP_15,
                            L1_2_L2_2_G1_MINI_ALU_BoothP_14,
                            L1_2_L2_2_G1_MINI_ALU_BoothP_13,
                            L1_2_L2_2_G1_MINI_ALU_BoothP_12,
                            L1_2_L2_2_G1_MINI_ALU_BoothP_11,
                            L1_2_L2_2_G1_MINI_ALU_BoothP_10,
                            L1_2_L2_2_G1_MINI_ALU_BoothP_9,
                            L1_2_L2_2_G1_MINI_ALU_BoothP_8,
                            L1_2_L2_2_G1_MINI_ALU_BoothP_7,
                            L1_2_L2_2_G1_MINI_ALU_BoothP_6,
                            L1_2_L2_2_G1_MINI_ALU_BoothP_5,
                            L1_2_L2_2_G1_MINI_ALU_BoothP_4,
                            L1_2_L2_2_G1_MINI_ALU_BoothP_3,
                            L1_2_L2_2_G1_MINI_ALU_BoothP_2,
                            L1_2_L2_2_G1_MINI_ALU_BoothP_1,\$dummy [455]}), .LargeWindowShifted (
                            {\$dummy [456],\$dummy [457],\$dummy [458],
                            \$dummy [459],\$dummy [460],\$dummy [461],
                            \$dummy [462],\$dummy [463],\$dummy [464],
                            \$dummy [465],\$dummy [466],\$dummy [467],
                            \$dummy [468],\$dummy [469],\$dummy [470],
                            \$dummy [471],\$dummy [472]})) ;
    booth_adder_17_unfolded4 L1_2_L2_3_G2_MINI_ALU_BOOTH_ADDER (.AdderFirstOperand (
                             {L1ResultsLarge_0__16,L1ResultsLarge_0__15,
                             L1ResultsLarge_0__14,L1ResultsLarge_0__13,
                             L1ResultsLarge_0__12,L1ResultsLarge_0__11,
                             L1ResultsLarge_0__10,L1ResultsLarge_0__9,
                             L1ResultsLarge_0__8,L1ResultsLarge_0__7,
                             L1ResultsLarge_0__6,L1ResultsLarge_0__5,
                             L1ResultsLarge_0__4,L1ResultsLarge_0__3,
                             L1ResultsLarge_0__2,L1ResultsLarge_0__1,
                             L1ResultsLarge_0__0}), .AdderSecondOperand ({
                             L1ResultsLarge_1__16,L1ResultsLarge_1__15,
                             L1ResultsLarge_1__14,L1ResultsLarge_1__13,
                             L1ResultsLarge_1__12,L1ResultsLarge_1__11,
                             L1ResultsLarge_1__10,L1ResultsLarge_1__9,
                             L1ResultsLarge_1__8,L1ResultsLarge_1__7,
                             L1ResultsLarge_1__6,L1ResultsLarge_1__5,
                             L1ResultsLarge_1__4,L1ResultsLarge_1__3,
                             L1ResultsLarge_1__2,L1ResultsLarge_1__1,
                             L1ResultsLarge_1__0}), .BoothOperand ({
                             L1_2_L2_3_G2_MINI_ALU_BoothOperand_16,
                             L1_2_L2_3_G2_MINI_ALU_BoothOperand_15,
                             L1_2_L2_3_G2_MINI_ALU_BoothOperand_14,
                             L1_2_L2_3_G2_MINI_ALU_BoothOperand_13,
                             L1_2_L2_3_G2_MINI_ALU_BoothOperand_12,
                             L1_2_L2_3_G2_MINI_ALU_BoothOperand_11,
                             L1_2_L2_3_G2_MINI_ALU_BoothOperand_10,
                             L1_2_L2_3_G2_MINI_ALU_BoothOperand_9,
                             L1FirstOperands_12__16,L1FirstOperands_12__16,
                             L1FirstOperands_12__16,L1FirstOperands_12__16,
                             L1FirstOperands_12__16,L1FirstOperands_12__16,
                             L1FirstOperands_12__16,L1FirstOperands_12__16,
                             L1FirstOperands_12__16}), .BoothP ({
                             L1_2_L2_3_G2_MINI_ALU_BoothP_16,
                             L1_2_L2_3_G2_MINI_ALU_BoothP_15,
                             L1_2_L2_3_G2_MINI_ALU_BoothP_14,
                             L1_2_L2_3_G2_MINI_ALU_BoothP_13,
                             L1_2_L2_3_G2_MINI_ALU_BoothP_12,
                             L1_2_L2_3_G2_MINI_ALU_BoothP_11,
                             L1_2_L2_3_G2_MINI_ALU_BoothP_10,
                             L1_2_L2_3_G2_MINI_ALU_BoothP_9,
                             L1_2_L2_3_G2_MINI_ALU_BoothP_8,
                             L1_2_L2_3_G2_MINI_ALU_BoothP_7,
                             L1_2_L2_3_G2_MINI_ALU_BoothP_6,
                             L1_2_L2_3_G2_MINI_ALU_BoothP_5,
                             L1_2_L2_3_G2_MINI_ALU_BoothP_4,
                             L1_2_L2_3_G2_MINI_ALU_BoothP_3,
                             L1_2_L2_3_G2_MINI_ALU_BoothP_2,
                             L1_2_L2_3_G2_MINI_ALU_BoothP_1,
                             L1_2_L2_3_G2_MINI_ALU_BoothP_0}), .SelOperand (
                             nx3287), .Operation (
                             L1_2_L2_3_G2_MINI_ALU_BoothXORCheck), .AdderResult (
                             {L2ResultsLarge_0__16,L2ResultsLarge_0__15,
                             L2ResultsLarge_0__14,L2ResultsLarge_0__13,
                             L2ResultsLarge_0__12,L2ResultsLarge_0__11,
                             L2ResultsLarge_0__10,L2ResultsLarge_0__9,
                             L2ResultsLarge_0__8,L2ResultsLarge_0__7,
                             L2ResultsLarge_0__6,L2ResultsLarge_0__5,
                             L2ResultsLarge_0__4,L2ResultsLarge_0__3,
                             L2ResultsLarge_0__2,L2ResultsLarge_0__1,
                             L2ResultsLarge_0__0}), .AdderBoothResult ({
                             \$dummy [473],
                             L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_15,
                             L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_14,
                             L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_13,
                             L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_12,
                             L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_11,
                             L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_10,
                             L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_9,
                             L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_8,
                             L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_7,
                             L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_6,
                             L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_5,
                             L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_4,
                             L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_3,
                             L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_2,
                             L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_1,
                             L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_0})) ;
    booth_unit_17 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT (.CLK (CLK), .RST (RST), .Start (
                  Start), .Instr (Instr), .LoopingAndResultNotReady (nx3277), .Filter (
                  {FilterDin_2__3__7,FilterDin_2__3__6,FilterDin_2__3__5,
                  FilterDin_2__3__4,FilterDin_2__3__3,FilterDin_2__3__2,
                  FilterDin_2__3__1,FilterDin_2__3__0}), .Window ({
                  WindowDin_2__3__7,WindowDin_2__3__6,WindowDin_2__3__5,
                  WindowDin_2__3__4,WindowDin_2__3__3,WindowDin_2__3__2,
                  WindowDin_2__3__1,WindowDin_2__3__0}), .AdderBoothResult ({
                  L1FirstOperands_12__16,
                  L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_15,
                  L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_14,
                  L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_13,
                  L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_12,
                  L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_11,
                  L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_10,
                  L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_9,
                  L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_8,
                  L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_7,
                  L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_6,
                  L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_5,
                  L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_4,
                  L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_3,
                  L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_2,
                  L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_1,
                  L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_0}), .BoothXORCheck (
                  L1_2_L2_3_G2_MINI_ALU_BoothXORCheck), .BoothResult ({
                  \$dummy [474],\$dummy [475],\$dummy [476],\$dummy [477],
                  \$dummy [478],\$dummy [479],\$dummy [480],\$dummy [481]}), .BoothAddingOperand (
                  {L1_2_L2_3_G2_MINI_ALU_BoothOperand_16,
                  L1_2_L2_3_G2_MINI_ALU_BoothOperand_15,
                  L1_2_L2_3_G2_MINI_ALU_BoothOperand_14,
                  L1_2_L2_3_G2_MINI_ALU_BoothOperand_13,
                  L1_2_L2_3_G2_MINI_ALU_BoothOperand_12,
                  L1_2_L2_3_G2_MINI_ALU_BoothOperand_11,
                  L1_2_L2_3_G2_MINI_ALU_BoothOperand_10,
                  L1_2_L2_3_G2_MINI_ALU_BoothOperand_9,\$dummy [482],
                  \$dummy [483],\$dummy [484],\$dummy [485],\$dummy [486],
                  \$dummy [487],\$dummy [488],\$dummy [489],\$dummy [490]}), .BoothP (
                  {L1_2_L2_3_G2_MINI_ALU_BoothP_16,
                  L1_2_L2_3_G2_MINI_ALU_BoothP_15,
                  L1_2_L2_3_G2_MINI_ALU_BoothP_14,
                  L1_2_L2_3_G2_MINI_ALU_BoothP_13,
                  L1_2_L2_3_G2_MINI_ALU_BoothP_12,
                  L1_2_L2_3_G2_MINI_ALU_BoothP_11,
                  L1_2_L2_3_G2_MINI_ALU_BoothP_10,L1_2_L2_3_G2_MINI_ALU_BoothP_9
                  ,L1_2_L2_3_G2_MINI_ALU_BoothP_8,L1_2_L2_3_G2_MINI_ALU_BoothP_7
                  ,L1_2_L2_3_G2_MINI_ALU_BoothP_6,L1_2_L2_3_G2_MINI_ALU_BoothP_5
                  ,L1_2_L2_3_G2_MINI_ALU_BoothP_4,L1_2_L2_3_G2_MINI_ALU_BoothP_3
                  ,L1_2_L2_3_G2_MINI_ALU_BoothP_2,L1_2_L2_3_G2_MINI_ALU_BoothP_1
                  ,L1_2_L2_3_G2_MINI_ALU_BoothP_0}), .LargeWindowShifted ({
                  \$dummy [491],\$dummy [492],\$dummy [493],\$dummy [494],
                  \$dummy [495],\$dummy [496],\$dummy [497],\$dummy [498],
                  \$dummy [499],\$dummy [500],\$dummy [501],\$dummy [502],
                  \$dummy [503],\$dummy [504],\$dummy [505],\$dummy [506],
                  \$dummy [507]})) ;
    booth_adder_17_unfolded4 L1_2_L2_4_G2_MINI_ALU_BOOTH_ADDER (.AdderFirstOperand (
                             {L1ResultsLarge_2__16,L1ResultsLarge_2__15,
                             L1ResultsLarge_2__14,L1ResultsLarge_2__13,
                             L1ResultsLarge_2__12,L1ResultsLarge_2__11,
                             L1ResultsLarge_2__10,L1ResultsLarge_2__9,
                             L1ResultsLarge_2__8,L1ResultsLarge_2__7,
                             L1ResultsLarge_2__6,L1ResultsLarge_2__5,
                             L1ResultsLarge_2__4,L1ResultsLarge_2__3,
                             L1ResultsLarge_2__2,L1ResultsLarge_2__1,
                             L1ResultsLarge_2__0}), .AdderSecondOperand ({
                             L1ResultsLarge_3__16,L1ResultsLarge_3__15,
                             L1ResultsLarge_3__14,L1ResultsLarge_3__13,
                             L1ResultsLarge_3__12,L1ResultsLarge_3__11,
                             L1ResultsLarge_3__10,L1ResultsLarge_3__9,
                             L1ResultsLarge_3__8,L1ResultsLarge_3__7,
                             L1ResultsLarge_3__6,L1ResultsLarge_3__5,
                             L1ResultsLarge_3__4,L1ResultsLarge_3__3,
                             L1ResultsLarge_3__2,L1ResultsLarge_3__1,
                             L1ResultsLarge_3__0}), .BoothOperand ({
                             L1_2_L2_4_G2_MINI_ALU_BoothOperand_16,
                             L1_2_L2_4_G2_MINI_ALU_BoothOperand_15,
                             L1_2_L2_4_G2_MINI_ALU_BoothOperand_14,
                             L1_2_L2_4_G2_MINI_ALU_BoothOperand_13,
                             L1_2_L2_4_G2_MINI_ALU_BoothOperand_12,
                             L1_2_L2_4_G2_MINI_ALU_BoothOperand_11,
                             L1_2_L2_4_G2_MINI_ALU_BoothOperand_10,
                             L1_2_L2_4_G2_MINI_ALU_BoothOperand_9,
                             L1FirstOperands_12__16,L1FirstOperands_12__16,
                             L1FirstOperands_12__16,L1FirstOperands_12__16,
                             L1FirstOperands_12__16,L1FirstOperands_12__16,
                             L1FirstOperands_12__16,L1FirstOperands_12__16,
                             L1FirstOperands_12__16}), .BoothP ({
                             L1_2_L2_4_G2_MINI_ALU_BoothP_16,
                             L1_2_L2_4_G2_MINI_ALU_BoothP_15,
                             L1_2_L2_4_G2_MINI_ALU_BoothP_14,
                             L1_2_L2_4_G2_MINI_ALU_BoothP_13,
                             L1_2_L2_4_G2_MINI_ALU_BoothP_12,
                             L1_2_L2_4_G2_MINI_ALU_BoothP_11,
                             L1_2_L2_4_G2_MINI_ALU_BoothP_10,
                             L1_2_L2_4_G2_MINI_ALU_BoothP_9,
                             L1_2_L2_4_G2_MINI_ALU_BoothP_8,
                             L1_2_L2_4_G2_MINI_ALU_BoothP_7,
                             L1_2_L2_4_G2_MINI_ALU_BoothP_6,
                             L1_2_L2_4_G2_MINI_ALU_BoothP_5,
                             L1_2_L2_4_G2_MINI_ALU_BoothP_4,
                             L1_2_L2_4_G2_MINI_ALU_BoothP_3,
                             L1_2_L2_4_G2_MINI_ALU_BoothP_2,
                             L1_2_L2_4_G2_MINI_ALU_BoothP_1,
                             L1_2_L2_4_G2_MINI_ALU_BoothP_0}), .SelOperand (
                             nx3287), .Operation (
                             L1_2_L2_4_G2_MINI_ALU_BoothXORCheck), .AdderResult (
                             {L2ResultsLarge_1__16,L2ResultsLarge_1__15,
                             L2ResultsLarge_1__14,L2ResultsLarge_1__13,
                             L2ResultsLarge_1__12,L2ResultsLarge_1__11,
                             L2ResultsLarge_1__10,L2ResultsLarge_1__9,
                             L2ResultsLarge_1__8,L2ResultsLarge_1__7,
                             L2ResultsLarge_1__6,L2ResultsLarge_1__5,
                             L2ResultsLarge_1__4,L2ResultsLarge_1__3,
                             L2ResultsLarge_1__2,L2ResultsLarge_1__1,
                             L2ResultsLarge_1__0}), .AdderBoothResult ({
                             \$dummy [508],
                             L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_15,
                             L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_14,
                             L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_13,
                             L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_12,
                             L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_11,
                             L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_10,
                             L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_9,
                             L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_8,
                             L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_7,
                             L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_6,
                             L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_5,
                             L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_4,
                             L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_3,
                             L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_2,
                             L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_1,
                             L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_0})) ;
    booth_unit_17 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT (.CLK (CLK), .RST (RST), .Start (
                  Start), .Instr (Instr), .LoopingAndResultNotReady (nx3279), .Filter (
                  {FilterDin_2__4__7,FilterDin_2__4__6,FilterDin_2__4__5,
                  FilterDin_2__4__4,FilterDin_2__4__3,FilterDin_2__4__2,
                  FilterDin_2__4__1,FilterDin_2__4__0}), .Window ({
                  WindowDin_2__4__7,WindowDin_2__4__6,WindowDin_2__4__5,
                  WindowDin_2__4__4,WindowDin_2__4__3,WindowDin_2__4__2,
                  WindowDin_2__4__1,WindowDin_2__4__0}), .AdderBoothResult ({
                  L1FirstOperands_12__16,
                  L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_15,
                  L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_14,
                  L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_13,
                  L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_12,
                  L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_11,
                  L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_10,
                  L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_9,
                  L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_8,
                  L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_7,
                  L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_6,
                  L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_5,
                  L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_4,
                  L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_3,
                  L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_2,
                  L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_1,
                  L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_0}), .BoothXORCheck (
                  L1_2_L2_4_G2_MINI_ALU_BoothXORCheck), .BoothResult ({
                  \$dummy [509],\$dummy [510],\$dummy [511],\$dummy [512],
                  \$dummy [513],\$dummy [514],\$dummy [515],\$dummy [516]}), .BoothAddingOperand (
                  {L1_2_L2_4_G2_MINI_ALU_BoothOperand_16,
                  L1_2_L2_4_G2_MINI_ALU_BoothOperand_15,
                  L1_2_L2_4_G2_MINI_ALU_BoothOperand_14,
                  L1_2_L2_4_G2_MINI_ALU_BoothOperand_13,
                  L1_2_L2_4_G2_MINI_ALU_BoothOperand_12,
                  L1_2_L2_4_G2_MINI_ALU_BoothOperand_11,
                  L1_2_L2_4_G2_MINI_ALU_BoothOperand_10,
                  L1_2_L2_4_G2_MINI_ALU_BoothOperand_9,\$dummy [517],
                  \$dummy [518],\$dummy [519],\$dummy [520],\$dummy [521],
                  \$dummy [522],\$dummy [523],\$dummy [524],\$dummy [525]}), .BoothP (
                  {L1_2_L2_4_G2_MINI_ALU_BoothP_16,
                  L1_2_L2_4_G2_MINI_ALU_BoothP_15,
                  L1_2_L2_4_G2_MINI_ALU_BoothP_14,
                  L1_2_L2_4_G2_MINI_ALU_BoothP_13,
                  L1_2_L2_4_G2_MINI_ALU_BoothP_12,
                  L1_2_L2_4_G2_MINI_ALU_BoothP_11,
                  L1_2_L2_4_G2_MINI_ALU_BoothP_10,L1_2_L2_4_G2_MINI_ALU_BoothP_9
                  ,L1_2_L2_4_G2_MINI_ALU_BoothP_8,L1_2_L2_4_G2_MINI_ALU_BoothP_7
                  ,L1_2_L2_4_G2_MINI_ALU_BoothP_6,L1_2_L2_4_G2_MINI_ALU_BoothP_5
                  ,L1_2_L2_4_G2_MINI_ALU_BoothP_4,L1_2_L2_4_G2_MINI_ALU_BoothP_3
                  ,L1_2_L2_4_G2_MINI_ALU_BoothP_2,L1_2_L2_4_G2_MINI_ALU_BoothP_1
                  ,L1_2_L2_4_G2_MINI_ALU_BoothP_0}), .LargeWindowShifted ({
                  \$dummy [526],\$dummy [527],\$dummy [528],\$dummy [529],
                  \$dummy [530],\$dummy [531],\$dummy [532],\$dummy [533],
                  \$dummy [534],\$dummy [535],\$dummy [536],\$dummy [537],
                  \$dummy [538],\$dummy [539],\$dummy [540],\$dummy [541],
                  \$dummy [542]})) ;
    booth_adder_17_unfolded4 L1_3_L2_0_G2_MINI_ALU_BOOTH_ADDER (.AdderFirstOperand (
                             {L1ResultsLarge_4__16,L1ResultsLarge_4__15,
                             L1ResultsLarge_4__14,L1ResultsLarge_4__13,
                             L1ResultsLarge_4__12,L1ResultsLarge_4__11,
                             L1ResultsLarge_4__10,L1ResultsLarge_4__9,
                             L1ResultsLarge_4__8,L1ResultsLarge_4__7,
                             L1ResultsLarge_4__6,L1ResultsLarge_4__5,
                             L1ResultsLarge_4__4,L1ResultsLarge_4__3,
                             L1ResultsLarge_4__2,L1ResultsLarge_4__1,
                             L1ResultsLarge_4__0}), .AdderSecondOperand ({
                             L1ResultsLarge_5__16,L1ResultsLarge_5__15,
                             L1ResultsLarge_5__14,L1ResultsLarge_5__13,
                             L1ResultsLarge_5__12,L1ResultsLarge_5__11,
                             L1ResultsLarge_5__10,L1ResultsLarge_5__9,
                             L1ResultsLarge_5__8,L1ResultsLarge_5__7,
                             L1ResultsLarge_5__6,L1ResultsLarge_5__5,
                             L1ResultsLarge_5__4,L1ResultsLarge_5__3,
                             L1ResultsLarge_5__2,L1ResultsLarge_5__1,
                             L1ResultsLarge_5__0}), .BoothOperand ({
                             L1_3_L2_0_G2_MINI_ALU_BoothOperand_16,
                             L1_3_L2_0_G2_MINI_ALU_BoothOperand_15,
                             L1_3_L2_0_G2_MINI_ALU_BoothOperand_14,
                             L1_3_L2_0_G2_MINI_ALU_BoothOperand_13,
                             L1_3_L2_0_G2_MINI_ALU_BoothOperand_12,
                             L1_3_L2_0_G2_MINI_ALU_BoothOperand_11,
                             L1_3_L2_0_G2_MINI_ALU_BoothOperand_10,
                             L1_3_L2_0_G2_MINI_ALU_BoothOperand_9,
                             L1FirstOperands_12__16,L1FirstOperands_12__16,
                             L1FirstOperands_12__16,L1FirstOperands_12__16,
                             L1FirstOperands_12__16,L1FirstOperands_12__16,
                             L1FirstOperands_12__16,L1FirstOperands_12__16,
                             L1FirstOperands_12__16}), .BoothP ({
                             L1_3_L2_0_G2_MINI_ALU_BoothP_16,
                             L1_3_L2_0_G2_MINI_ALU_BoothP_15,
                             L1_3_L2_0_G2_MINI_ALU_BoothP_14,
                             L1_3_L2_0_G2_MINI_ALU_BoothP_13,
                             L1_3_L2_0_G2_MINI_ALU_BoothP_12,
                             L1_3_L2_0_G2_MINI_ALU_BoothP_11,
                             L1_3_L2_0_G2_MINI_ALU_BoothP_10,
                             L1_3_L2_0_G2_MINI_ALU_BoothP_9,
                             L1_3_L2_0_G2_MINI_ALU_BoothP_8,
                             L1_3_L2_0_G2_MINI_ALU_BoothP_7,
                             L1_3_L2_0_G2_MINI_ALU_BoothP_6,
                             L1_3_L2_0_G2_MINI_ALU_BoothP_5,
                             L1_3_L2_0_G2_MINI_ALU_BoothP_4,
                             L1_3_L2_0_G2_MINI_ALU_BoothP_3,
                             L1_3_L2_0_G2_MINI_ALU_BoothP_2,
                             L1_3_L2_0_G2_MINI_ALU_BoothP_1,
                             L1_3_L2_0_G2_MINI_ALU_BoothP_0}), .SelOperand (
                             nx3287), .Operation (
                             L1_3_L2_0_G2_MINI_ALU_BoothXORCheck), .AdderResult (
                             {L2ResultsLarge_2__16,L2ResultsLarge_2__15,
                             L2ResultsLarge_2__14,L2ResultsLarge_2__13,
                             L2ResultsLarge_2__12,L2ResultsLarge_2__11,
                             L2ResultsLarge_2__10,L2ResultsLarge_2__9,
                             L2ResultsLarge_2__8,L2ResultsLarge_2__7,
                             L2ResultsLarge_2__6,L2ResultsLarge_2__5,
                             L2ResultsLarge_2__4,L2ResultsLarge_2__3,
                             L2ResultsLarge_2__2,L2ResultsLarge_2__1,
                             L2ResultsLarge_2__0}), .AdderBoothResult ({
                             \$dummy [543],
                             L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_15,
                             L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_14,
                             L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_13,
                             L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_12,
                             L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_11,
                             L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_10,
                             L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_9,
                             L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_8,
                             L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_7,
                             L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_6,
                             L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_5,
                             L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_4,
                             L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_3,
                             L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_2,
                             L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_1,
                             L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_0})) ;
    booth_unit_17 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT (.CLK (CLK), .RST (RST), .Start (
                  Start), .Instr (Instr), .LoopingAndResultNotReady (nx3279), .Filter (
                  {FilterDin_3__0__7,FilterDin_3__0__6,FilterDin_3__0__5,
                  FilterDin_3__0__4,FilterDin_3__0__3,FilterDin_3__0__2,
                  FilterDin_3__0__1,FilterDin_3__0__0}), .Window ({
                  WindowDin_3__0__7,WindowDin_3__0__6,WindowDin_3__0__5,
                  WindowDin_3__0__4,WindowDin_3__0__3,WindowDin_3__0__2,
                  WindowDin_3__0__1,WindowDin_3__0__0}), .AdderBoothResult ({
                  L1FirstOperands_12__16,
                  L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_15,
                  L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_14,
                  L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_13,
                  L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_12,
                  L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_11,
                  L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_10,
                  L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_9,
                  L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_8,
                  L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_7,
                  L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_6,
                  L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_5,
                  L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_4,
                  L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_3,
                  L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_2,
                  L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_1,
                  L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_0}), .BoothXORCheck (
                  L1_3_L2_0_G2_MINI_ALU_BoothXORCheck), .BoothResult ({
                  \$dummy [544],\$dummy [545],\$dummy [546],\$dummy [547],
                  \$dummy [548],\$dummy [549],\$dummy [550],\$dummy [551]}), .BoothAddingOperand (
                  {L1_3_L2_0_G2_MINI_ALU_BoothOperand_16,
                  L1_3_L2_0_G2_MINI_ALU_BoothOperand_15,
                  L1_3_L2_0_G2_MINI_ALU_BoothOperand_14,
                  L1_3_L2_0_G2_MINI_ALU_BoothOperand_13,
                  L1_3_L2_0_G2_MINI_ALU_BoothOperand_12,
                  L1_3_L2_0_G2_MINI_ALU_BoothOperand_11,
                  L1_3_L2_0_G2_MINI_ALU_BoothOperand_10,
                  L1_3_L2_0_G2_MINI_ALU_BoothOperand_9,\$dummy [552],
                  \$dummy [553],\$dummy [554],\$dummy [555],\$dummy [556],
                  \$dummy [557],\$dummy [558],\$dummy [559],\$dummy [560]}), .BoothP (
                  {L1_3_L2_0_G2_MINI_ALU_BoothP_16,
                  L1_3_L2_0_G2_MINI_ALU_BoothP_15,
                  L1_3_L2_0_G2_MINI_ALU_BoothP_14,
                  L1_3_L2_0_G2_MINI_ALU_BoothP_13,
                  L1_3_L2_0_G2_MINI_ALU_BoothP_12,
                  L1_3_L2_0_G2_MINI_ALU_BoothP_11,
                  L1_3_L2_0_G2_MINI_ALU_BoothP_10,L1_3_L2_0_G2_MINI_ALU_BoothP_9
                  ,L1_3_L2_0_G2_MINI_ALU_BoothP_8,L1_3_L2_0_G2_MINI_ALU_BoothP_7
                  ,L1_3_L2_0_G2_MINI_ALU_BoothP_6,L1_3_L2_0_G2_MINI_ALU_BoothP_5
                  ,L1_3_L2_0_G2_MINI_ALU_BoothP_4,L1_3_L2_0_G2_MINI_ALU_BoothP_3
                  ,L1_3_L2_0_G2_MINI_ALU_BoothP_2,L1_3_L2_0_G2_MINI_ALU_BoothP_1
                  ,L1_3_L2_0_G2_MINI_ALU_BoothP_0}), .LargeWindowShifted ({
                  \$dummy [561],\$dummy [562],\$dummy [563],\$dummy [564],
                  \$dummy [565],\$dummy [566],\$dummy [567],\$dummy [568],
                  \$dummy [569],\$dummy [570],\$dummy [571],\$dummy [572],
                  \$dummy [573],\$dummy [574],\$dummy [575],\$dummy [576],
                  \$dummy [577]})) ;
    booth_adder_17_unfolded4 L1_3_L2_1_G2_MINI_ALU_BOOTH_ADDER (.AdderFirstOperand (
                             {L1ResultsLarge_6__16,L1ResultsLarge_6__15,
                             L1ResultsLarge_6__14,L1ResultsLarge_6__13,
                             L1ResultsLarge_6__12,L1ResultsLarge_6__11,
                             L1ResultsLarge_6__10,L1ResultsLarge_6__9,
                             L1ResultsLarge_6__8,L1ResultsLarge_6__7,
                             L1ResultsLarge_6__6,L1ResultsLarge_6__5,
                             L1ResultsLarge_6__4,L1ResultsLarge_6__3,
                             L1ResultsLarge_6__2,L1ResultsLarge_6__1,
                             L1ResultsLarge_6__0}), .AdderSecondOperand ({
                             L1ResultsLarge_7__16,L1ResultsLarge_7__15,
                             L1ResultsLarge_7__14,L1ResultsLarge_7__13,
                             L1ResultsLarge_7__12,L1ResultsLarge_7__11,
                             L1ResultsLarge_7__10,L1ResultsLarge_7__9,
                             L1ResultsLarge_7__8,L1ResultsLarge_7__7,
                             L1ResultsLarge_7__6,L1ResultsLarge_7__5,
                             L1ResultsLarge_7__4,L1ResultsLarge_7__3,
                             L1ResultsLarge_7__2,L1ResultsLarge_7__1,
                             L1ResultsLarge_7__0}), .BoothOperand ({
                             L1_3_L2_1_G2_MINI_ALU_BoothOperand_16,
                             L1_3_L2_1_G2_MINI_ALU_BoothOperand_15,
                             L1_3_L2_1_G2_MINI_ALU_BoothOperand_14,
                             L1_3_L2_1_G2_MINI_ALU_BoothOperand_13,
                             L1_3_L2_1_G2_MINI_ALU_BoothOperand_12,
                             L1_3_L2_1_G2_MINI_ALU_BoothOperand_11,
                             L1_3_L2_1_G2_MINI_ALU_BoothOperand_10,
                             L1_3_L2_1_G2_MINI_ALU_BoothOperand_9,
                             L1FirstOperands_12__16,L1FirstOperands_12__16,
                             L1FirstOperands_12__16,L1FirstOperands_12__16,
                             L1FirstOperands_12__16,L1FirstOperands_12__16,
                             L1FirstOperands_12__16,L1FirstOperands_12__16,
                             L1FirstOperands_12__16}), .BoothP ({
                             L1_3_L2_1_G2_MINI_ALU_BoothP_16,
                             L1_3_L2_1_G2_MINI_ALU_BoothP_15,
                             L1_3_L2_1_G2_MINI_ALU_BoothP_14,
                             L1_3_L2_1_G2_MINI_ALU_BoothP_13,
                             L1_3_L2_1_G2_MINI_ALU_BoothP_12,
                             L1_3_L2_1_G2_MINI_ALU_BoothP_11,
                             L1_3_L2_1_G2_MINI_ALU_BoothP_10,
                             L1_3_L2_1_G2_MINI_ALU_BoothP_9,
                             L1_3_L2_1_G2_MINI_ALU_BoothP_8,
                             L1_3_L2_1_G2_MINI_ALU_BoothP_7,
                             L1_3_L2_1_G2_MINI_ALU_BoothP_6,
                             L1_3_L2_1_G2_MINI_ALU_BoothP_5,
                             L1_3_L2_1_G2_MINI_ALU_BoothP_4,
                             L1_3_L2_1_G2_MINI_ALU_BoothP_3,
                             L1_3_L2_1_G2_MINI_ALU_BoothP_2,
                             L1_3_L2_1_G2_MINI_ALU_BoothP_1,
                             L1_3_L2_1_G2_MINI_ALU_BoothP_0}), .SelOperand (
                             nx3285), .Operation (
                             L1_3_L2_1_G2_MINI_ALU_BoothXORCheck), .AdderResult (
                             {L2ResultsLarge_3__16,L2ResultsLarge_3__15,
                             L2ResultsLarge_3__14,L2ResultsLarge_3__13,
                             L2ResultsLarge_3__12,L2ResultsLarge_3__11,
                             L2ResultsLarge_3__10,L2ResultsLarge_3__9,
                             L2ResultsLarge_3__8,L2ResultsLarge_3__7,
                             L2ResultsLarge_3__6,L2ResultsLarge_3__5,
                             L2ResultsLarge_3__4,L2ResultsLarge_3__3,
                             L2ResultsLarge_3__2,L2ResultsLarge_3__1,
                             L2ResultsLarge_3__0}), .AdderBoothResult ({
                             \$dummy [578],
                             L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_15,
                             L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_14,
                             L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_13,
                             L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_12,
                             L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_11,
                             L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_10,
                             L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_9,
                             L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_8,
                             L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_7,
                             L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_6,
                             L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_5,
                             L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_4,
                             L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_3,
                             L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_2,
                             L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_1,
                             L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_0})) ;
    booth_unit_17 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT (.CLK (CLK), .RST (RST), .Start (
                  Start), .Instr (Instr), .LoopingAndResultNotReady (nx3279), .Filter (
                  {FilterDin_3__1__7,FilterDin_3__1__6,FilterDin_3__1__5,
                  FilterDin_3__1__4,FilterDin_3__1__3,FilterDin_3__1__2,
                  FilterDin_3__1__1,FilterDin_3__1__0}), .Window ({
                  WindowDin_3__1__7,WindowDin_3__1__6,WindowDin_3__1__5,
                  WindowDin_3__1__4,WindowDin_3__1__3,WindowDin_3__1__2,
                  WindowDin_3__1__1,WindowDin_3__1__0}), .AdderBoothResult ({
                  L1FirstOperands_12__16,
                  L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_15,
                  L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_14,
                  L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_13,
                  L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_12,
                  L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_11,
                  L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_10,
                  L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_9,
                  L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_8,
                  L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_7,
                  L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_6,
                  L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_5,
                  L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_4,
                  L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_3,
                  L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_2,
                  L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_1,
                  L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_0}), .BoothXORCheck (
                  L1_3_L2_1_G2_MINI_ALU_BoothXORCheck), .BoothResult ({
                  \$dummy [579],\$dummy [580],\$dummy [581],\$dummy [582],
                  \$dummy [583],\$dummy [584],\$dummy [585],\$dummy [586]}), .BoothAddingOperand (
                  {L1_3_L2_1_G2_MINI_ALU_BoothOperand_16,
                  L1_3_L2_1_G2_MINI_ALU_BoothOperand_15,
                  L1_3_L2_1_G2_MINI_ALU_BoothOperand_14,
                  L1_3_L2_1_G2_MINI_ALU_BoothOperand_13,
                  L1_3_L2_1_G2_MINI_ALU_BoothOperand_12,
                  L1_3_L2_1_G2_MINI_ALU_BoothOperand_11,
                  L1_3_L2_1_G2_MINI_ALU_BoothOperand_10,
                  L1_3_L2_1_G2_MINI_ALU_BoothOperand_9,\$dummy [587],
                  \$dummy [588],\$dummy [589],\$dummy [590],\$dummy [591],
                  \$dummy [592],\$dummy [593],\$dummy [594],\$dummy [595]}), .BoothP (
                  {L1_3_L2_1_G2_MINI_ALU_BoothP_16,
                  L1_3_L2_1_G2_MINI_ALU_BoothP_15,
                  L1_3_L2_1_G2_MINI_ALU_BoothP_14,
                  L1_3_L2_1_G2_MINI_ALU_BoothP_13,
                  L1_3_L2_1_G2_MINI_ALU_BoothP_12,
                  L1_3_L2_1_G2_MINI_ALU_BoothP_11,
                  L1_3_L2_1_G2_MINI_ALU_BoothP_10,L1_3_L2_1_G2_MINI_ALU_BoothP_9
                  ,L1_3_L2_1_G2_MINI_ALU_BoothP_8,L1_3_L2_1_G2_MINI_ALU_BoothP_7
                  ,L1_3_L2_1_G2_MINI_ALU_BoothP_6,L1_3_L2_1_G2_MINI_ALU_BoothP_5
                  ,L1_3_L2_1_G2_MINI_ALU_BoothP_4,L1_3_L2_1_G2_MINI_ALU_BoothP_3
                  ,L1_3_L2_1_G2_MINI_ALU_BoothP_2,L1_3_L2_1_G2_MINI_ALU_BoothP_1
                  ,L1_3_L2_1_G2_MINI_ALU_BoothP_0}), .LargeWindowShifted ({
                  \$dummy [596],\$dummy [597],\$dummy [598],\$dummy [599],
                  \$dummy [600],\$dummy [601],\$dummy [602],\$dummy [603],
                  \$dummy [604],\$dummy [605],\$dummy [606],\$dummy [607],
                  \$dummy [608],\$dummy [609],\$dummy [610],\$dummy [611],
                  \$dummy [612]})) ;
    booth_adder_17_unfolded4 L1_3_L2_2_G2_MINI_ALU_BOOTH_ADDER (.AdderFirstOperand (
                             {L1ResultsLarge_8__16,L1ResultsLarge_8__15,
                             L1ResultsLarge_8__14,L1ResultsLarge_8__13,
                             L1ResultsLarge_8__12,L1ResultsLarge_8__11,
                             L1ResultsLarge_8__10,L1ResultsLarge_8__9,
                             L1ResultsLarge_8__8,L1ResultsLarge_8__7,
                             L1ResultsLarge_8__6,L1ResultsLarge_8__5,
                             L1ResultsLarge_8__4,L1ResultsLarge_8__3,
                             L1ResultsLarge_8__2,L1ResultsLarge_8__1,
                             L1ResultsLarge_8__0}), .AdderSecondOperand ({
                             L1ResultsLarge_9__16,L1ResultsLarge_9__15,
                             L1ResultsLarge_9__14,L1ResultsLarge_9__13,
                             L1ResultsLarge_9__12,L1ResultsLarge_9__11,
                             L1ResultsLarge_9__10,L1ResultsLarge_9__9,
                             L1ResultsLarge_9__8,L1ResultsLarge_9__7,
                             L1ResultsLarge_9__6,L1ResultsLarge_9__5,
                             L1ResultsLarge_9__4,L1ResultsLarge_9__3,
                             L1ResultsLarge_9__2,L1ResultsLarge_9__1,
                             L1ResultsLarge_9__0}), .BoothOperand ({
                             L1_3_L2_2_G2_MINI_ALU_BoothOperand_16,
                             L1_3_L2_2_G2_MINI_ALU_BoothOperand_15,
                             L1_3_L2_2_G2_MINI_ALU_BoothOperand_14,
                             L1_3_L2_2_G2_MINI_ALU_BoothOperand_13,
                             L1_3_L2_2_G2_MINI_ALU_BoothOperand_12,
                             L1_3_L2_2_G2_MINI_ALU_BoothOperand_11,
                             L1_3_L2_2_G2_MINI_ALU_BoothOperand_10,
                             L1_3_L2_2_G2_MINI_ALU_BoothOperand_9,
                             L1FirstOperands_12__16,L1FirstOperands_12__16,
                             L1FirstOperands_12__16,L1FirstOperands_12__16,
                             L1FirstOperands_12__16,L1FirstOperands_12__16,
                             L1FirstOperands_12__16,L1FirstOperands_12__16,
                             L1FirstOperands_12__16}), .BoothP ({
                             L1_3_L2_2_G2_MINI_ALU_BoothP_16,
                             L1_3_L2_2_G2_MINI_ALU_BoothP_15,
                             L1_3_L2_2_G2_MINI_ALU_BoothP_14,
                             L1_3_L2_2_G2_MINI_ALU_BoothP_13,
                             L1_3_L2_2_G2_MINI_ALU_BoothP_12,
                             L1_3_L2_2_G2_MINI_ALU_BoothP_11,
                             L1_3_L2_2_G2_MINI_ALU_BoothP_10,
                             L1_3_L2_2_G2_MINI_ALU_BoothP_9,
                             L1_3_L2_2_G2_MINI_ALU_BoothP_8,
                             L1_3_L2_2_G2_MINI_ALU_BoothP_7,
                             L1_3_L2_2_G2_MINI_ALU_BoothP_6,
                             L1_3_L2_2_G2_MINI_ALU_BoothP_5,
                             L1_3_L2_2_G2_MINI_ALU_BoothP_4,
                             L1_3_L2_2_G2_MINI_ALU_BoothP_3,
                             L1_3_L2_2_G2_MINI_ALU_BoothP_2,
                             L1_3_L2_2_G2_MINI_ALU_BoothP_1,
                             L1_3_L2_2_G2_MINI_ALU_BoothP_0}), .SelOperand (
                             nx3287), .Operation (
                             L1_3_L2_2_G2_MINI_ALU_BoothXORCheck), .AdderResult (
                             {L2ResultsLarge_4__16,L2ResultsLarge_4__15,
                             L2ResultsLarge_4__14,L2ResultsLarge_4__13,
                             L2ResultsLarge_4__12,L2ResultsLarge_4__11,
                             L2ResultsLarge_4__10,L2ResultsLarge_4__9,
                             L2ResultsLarge_4__8,L2ResultsLarge_4__7,
                             L2ResultsLarge_4__6,L2ResultsLarge_4__5,
                             L2ResultsLarge_4__4,L2ResultsLarge_4__3,
                             L2ResultsLarge_4__2,L2ResultsLarge_4__1,
                             L2ResultsLarge_4__0}), .AdderBoothResult ({
                             \$dummy [613],
                             L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_15,
                             L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_14,
                             L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_13,
                             L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_12,
                             L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_11,
                             L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_10,
                             L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_9,
                             L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_8,
                             L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_7,
                             L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_6,
                             L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_5,
                             L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_4,
                             L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_3,
                             L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_2,
                             L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_1,
                             L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_0})) ;
    booth_unit_17 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT (.CLK (CLK), .RST (RST), .Start (
                  Start), .Instr (Instr), .LoopingAndResultNotReady (nx3279), .Filter (
                  {FilterDin_3__2__7,FilterDin_3__2__6,FilterDin_3__2__5,
                  FilterDin_3__2__4,FilterDin_3__2__3,FilterDin_3__2__2,
                  FilterDin_3__2__1,FilterDin_3__2__0}), .Window ({
                  WindowDin_3__2__7,WindowDin_3__2__6,WindowDin_3__2__5,
                  WindowDin_3__2__4,WindowDin_3__2__3,WindowDin_3__2__2,
                  WindowDin_3__2__1,WindowDin_3__2__0}), .AdderBoothResult ({
                  L1FirstOperands_12__16,
                  L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_15,
                  L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_14,
                  L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_13,
                  L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_12,
                  L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_11,
                  L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_10,
                  L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_9,
                  L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_8,
                  L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_7,
                  L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_6,
                  L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_5,
                  L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_4,
                  L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_3,
                  L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_2,
                  L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_1,
                  L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_0}), .BoothXORCheck (
                  L1_3_L2_2_G2_MINI_ALU_BoothXORCheck), .BoothResult ({
                  \$dummy [614],\$dummy [615],\$dummy [616],\$dummy [617],
                  \$dummy [618],\$dummy [619],\$dummy [620],\$dummy [621]}), .BoothAddingOperand (
                  {L1_3_L2_2_G2_MINI_ALU_BoothOperand_16,
                  L1_3_L2_2_G2_MINI_ALU_BoothOperand_15,
                  L1_3_L2_2_G2_MINI_ALU_BoothOperand_14,
                  L1_3_L2_2_G2_MINI_ALU_BoothOperand_13,
                  L1_3_L2_2_G2_MINI_ALU_BoothOperand_12,
                  L1_3_L2_2_G2_MINI_ALU_BoothOperand_11,
                  L1_3_L2_2_G2_MINI_ALU_BoothOperand_10,
                  L1_3_L2_2_G2_MINI_ALU_BoothOperand_9,\$dummy [622],
                  \$dummy [623],\$dummy [624],\$dummy [625],\$dummy [626],
                  \$dummy [627],\$dummy [628],\$dummy [629],\$dummy [630]}), .BoothP (
                  {L1_3_L2_2_G2_MINI_ALU_BoothP_16,
                  L1_3_L2_2_G2_MINI_ALU_BoothP_15,
                  L1_3_L2_2_G2_MINI_ALU_BoothP_14,
                  L1_3_L2_2_G2_MINI_ALU_BoothP_13,
                  L1_3_L2_2_G2_MINI_ALU_BoothP_12,
                  L1_3_L2_2_G2_MINI_ALU_BoothP_11,
                  L1_3_L2_2_G2_MINI_ALU_BoothP_10,L1_3_L2_2_G2_MINI_ALU_BoothP_9
                  ,L1_3_L2_2_G2_MINI_ALU_BoothP_8,L1_3_L2_2_G2_MINI_ALU_BoothP_7
                  ,L1_3_L2_2_G2_MINI_ALU_BoothP_6,L1_3_L2_2_G2_MINI_ALU_BoothP_5
                  ,L1_3_L2_2_G2_MINI_ALU_BoothP_4,L1_3_L2_2_G2_MINI_ALU_BoothP_3
                  ,L1_3_L2_2_G2_MINI_ALU_BoothP_2,L1_3_L2_2_G2_MINI_ALU_BoothP_1
                  ,L1_3_L2_2_G2_MINI_ALU_BoothP_0}), .LargeWindowShifted ({
                  \$dummy [631],\$dummy [632],\$dummy [633],\$dummy [634],
                  \$dummy [635],\$dummy [636],\$dummy [637],\$dummy [638],
                  \$dummy [639],\$dummy [640],\$dummy [641],\$dummy [642],
                  \$dummy [643],\$dummy [644],\$dummy [645],\$dummy [646],
                  \$dummy [647]})) ;
    booth_adder_17_unfolded4 L1_3_L2_3_G2_MINI_ALU_BOOTH_ADDER (.AdderFirstOperand (
                             {L1ResultsLarge_10__16,L1ResultsLarge_10__15,
                             L1ResultsLarge_10__14,L1ResultsLarge_10__13,
                             L1ResultsLarge_10__12,L1ResultsLarge_10__11,
                             L1ResultsLarge_10__10,L1ResultsLarge_10__9,
                             L1ResultsLarge_10__8,L1ResultsLarge_10__7,
                             L1ResultsLarge_10__6,L1ResultsLarge_10__5,
                             L1ResultsLarge_10__4,L1ResultsLarge_10__3,
                             L1ResultsLarge_10__2,L1ResultsLarge_10__1,
                             L1ResultsLarge_10__0}), .AdderSecondOperand ({
                             L1ResultsLarge_11__16,L1ResultsLarge_11__15,
                             L1ResultsLarge_11__14,L1ResultsLarge_11__13,
                             L1ResultsLarge_11__12,L1ResultsLarge_11__11,
                             L1ResultsLarge_11__10,L1ResultsLarge_11__9,
                             L1ResultsLarge_11__8,L1ResultsLarge_11__7,
                             L1ResultsLarge_11__6,L1ResultsLarge_11__5,
                             L1ResultsLarge_11__4,L1ResultsLarge_11__3,
                             L1ResultsLarge_11__2,L1ResultsLarge_11__1,
                             L1ResultsLarge_11__0}), .BoothOperand ({
                             L1_3_L2_3_G2_MINI_ALU_BoothOperand_16,
                             L1_3_L2_3_G2_MINI_ALU_BoothOperand_15,
                             L1_3_L2_3_G2_MINI_ALU_BoothOperand_14,
                             L1_3_L2_3_G2_MINI_ALU_BoothOperand_13,
                             L1_3_L2_3_G2_MINI_ALU_BoothOperand_12,
                             L1_3_L2_3_G2_MINI_ALU_BoothOperand_11,
                             L1_3_L2_3_G2_MINI_ALU_BoothOperand_10,
                             L1_3_L2_3_G2_MINI_ALU_BoothOperand_9,
                             L1FirstOperands_12__16,L1FirstOperands_12__16,
                             L1FirstOperands_12__16,L1FirstOperands_12__16,
                             L1FirstOperands_12__16,L1FirstOperands_12__16,
                             L1FirstOperands_12__16,L1FirstOperands_12__16,
                             L1FirstOperands_12__16}), .BoothP ({
                             L1_3_L2_3_G2_MINI_ALU_BoothP_16,
                             L1_3_L2_3_G2_MINI_ALU_BoothP_15,
                             L1_3_L2_3_G2_MINI_ALU_BoothP_14,
                             L1_3_L2_3_G2_MINI_ALU_BoothP_13,
                             L1_3_L2_3_G2_MINI_ALU_BoothP_12,
                             L1_3_L2_3_G2_MINI_ALU_BoothP_11,
                             L1_3_L2_3_G2_MINI_ALU_BoothP_10,
                             L1_3_L2_3_G2_MINI_ALU_BoothP_9,
                             L1_3_L2_3_G2_MINI_ALU_BoothP_8,
                             L1_3_L2_3_G2_MINI_ALU_BoothP_7,
                             L1_3_L2_3_G2_MINI_ALU_BoothP_6,
                             L1_3_L2_3_G2_MINI_ALU_BoothP_5,
                             L1_3_L2_3_G2_MINI_ALU_BoothP_4,
                             L1_3_L2_3_G2_MINI_ALU_BoothP_3,
                             L1_3_L2_3_G2_MINI_ALU_BoothP_2,
                             L1_3_L2_3_G2_MINI_ALU_BoothP_1,
                             L1_3_L2_3_G2_MINI_ALU_BoothP_0}), .SelOperand (
                             nx3287), .Operation (
                             L1_3_L2_3_G2_MINI_ALU_BoothXORCheck), .AdderResult (
                             {L2ResultsLarge_5__16,L2ResultsLarge_5__15,
                             L2ResultsLarge_5__14,L2ResultsLarge_5__13,
                             L2ResultsLarge_5__12,L2ResultsLarge_5__11,
                             L2ResultsLarge_5__10,L2ResultsLarge_5__9,
                             L2ResultsLarge_5__8,L2ResultsLarge_5__7,
                             L2ResultsLarge_5__6,L2ResultsLarge_5__5,
                             L2ResultsLarge_5__4,L2ResultsLarge_5__3,
                             L2ResultsLarge_5__2,L2ResultsLarge_5__1,
                             L2ResultsLarge_5__0}), .AdderBoothResult ({
                             \$dummy [648],
                             L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_15,
                             L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_14,
                             L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_13,
                             L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_12,
                             L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_11,
                             L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_10,
                             L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_9,
                             L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_8,
                             L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_7,
                             L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_6,
                             L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_5,
                             L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_4,
                             L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_3,
                             L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_2,
                             L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_1,
                             L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_0})) ;
    booth_unit_17 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT (.CLK (CLK), .RST (RST), .Start (
                  Start), .Instr (Instr), .LoopingAndResultNotReady (nx3279), .Filter (
                  {FilterDin_3__3__7,FilterDin_3__3__6,FilterDin_3__3__5,
                  FilterDin_3__3__4,FilterDin_3__3__3,FilterDin_3__3__2,
                  FilterDin_3__3__1,FilterDin_3__3__0}), .Window ({
                  WindowDin_3__3__7,WindowDin_3__3__6,WindowDin_3__3__5,
                  WindowDin_3__3__4,WindowDin_3__3__3,WindowDin_3__3__2,
                  WindowDin_3__3__1,WindowDin_3__3__0}), .AdderBoothResult ({
                  L1FirstOperands_12__16,
                  L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_15,
                  L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_14,
                  L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_13,
                  L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_12,
                  L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_11,
                  L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_10,
                  L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_9,
                  L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_8,
                  L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_7,
                  L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_6,
                  L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_5,
                  L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_4,
                  L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_3,
                  L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_2,
                  L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_1,
                  L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_0}), .BoothXORCheck (
                  L1_3_L2_3_G2_MINI_ALU_BoothXORCheck), .BoothResult ({
                  \$dummy [649],\$dummy [650],\$dummy [651],\$dummy [652],
                  \$dummy [653],\$dummy [654],\$dummy [655],\$dummy [656]}), .BoothAddingOperand (
                  {L1_3_L2_3_G2_MINI_ALU_BoothOperand_16,
                  L1_3_L2_3_G2_MINI_ALU_BoothOperand_15,
                  L1_3_L2_3_G2_MINI_ALU_BoothOperand_14,
                  L1_3_L2_3_G2_MINI_ALU_BoothOperand_13,
                  L1_3_L2_3_G2_MINI_ALU_BoothOperand_12,
                  L1_3_L2_3_G2_MINI_ALU_BoothOperand_11,
                  L1_3_L2_3_G2_MINI_ALU_BoothOperand_10,
                  L1_3_L2_3_G2_MINI_ALU_BoothOperand_9,\$dummy [657],
                  \$dummy [658],\$dummy [659],\$dummy [660],\$dummy [661],
                  \$dummy [662],\$dummy [663],\$dummy [664],\$dummy [665]}), .BoothP (
                  {L1_3_L2_3_G2_MINI_ALU_BoothP_16,
                  L1_3_L2_3_G2_MINI_ALU_BoothP_15,
                  L1_3_L2_3_G2_MINI_ALU_BoothP_14,
                  L1_3_L2_3_G2_MINI_ALU_BoothP_13,
                  L1_3_L2_3_G2_MINI_ALU_BoothP_12,
                  L1_3_L2_3_G2_MINI_ALU_BoothP_11,
                  L1_3_L2_3_G2_MINI_ALU_BoothP_10,L1_3_L2_3_G2_MINI_ALU_BoothP_9
                  ,L1_3_L2_3_G2_MINI_ALU_BoothP_8,L1_3_L2_3_G2_MINI_ALU_BoothP_7
                  ,L1_3_L2_3_G2_MINI_ALU_BoothP_6,L1_3_L2_3_G2_MINI_ALU_BoothP_5
                  ,L1_3_L2_3_G2_MINI_ALU_BoothP_4,L1_3_L2_3_G2_MINI_ALU_BoothP_3
                  ,L1_3_L2_3_G2_MINI_ALU_BoothP_2,L1_3_L2_3_G2_MINI_ALU_BoothP_1
                  ,L1_3_L2_3_G2_MINI_ALU_BoothP_0}), .LargeWindowShifted ({
                  \$dummy [666],\$dummy [667],\$dummy [668],\$dummy [669],
                  \$dummy [670],\$dummy [671],\$dummy [672],\$dummy [673],
                  \$dummy [674],\$dummy [675],\$dummy [676],\$dummy [677],
                  \$dummy [678],\$dummy [679],\$dummy [680],\$dummy [681],
                  \$dummy [682]})) ;
    booth_adder_17_unfolded4 L1_3_L2_4_G3_MINI_ALU_BOOTH_ADDER (.AdderFirstOperand (
                             {L2ResultsLarge_0__16,L2ResultsLarge_0__15,
                             L2ResultsLarge_0__14,L2ResultsLarge_0__13,
                             L2ResultsLarge_0__12,L2ResultsLarge_0__11,
                             L2ResultsLarge_0__10,L2ResultsLarge_0__9,
                             L2ResultsLarge_0__8,L2ResultsLarge_0__7,
                             L2ResultsLarge_0__6,L2ResultsLarge_0__5,
                             L2ResultsLarge_0__4,L2ResultsLarge_0__3,
                             L2ResultsLarge_0__2,L2ResultsLarge_0__1,
                             L2ResultsLarge_0__0}), .AdderSecondOperand ({
                             L2ResultsLarge_1__16,L2ResultsLarge_1__15,
                             L2ResultsLarge_1__14,L2ResultsLarge_1__13,
                             L2ResultsLarge_1__12,L2ResultsLarge_1__11,
                             L2ResultsLarge_1__10,L2ResultsLarge_1__9,
                             L2ResultsLarge_1__8,L2ResultsLarge_1__7,
                             L2ResultsLarge_1__6,L2ResultsLarge_1__5,
                             L2ResultsLarge_1__4,L2ResultsLarge_1__3,
                             L2ResultsLarge_1__2,L2ResultsLarge_1__1,
                             L2ResultsLarge_1__0}), .BoothOperand ({
                             L1_3_L2_4_G3_MINI_ALU_BoothOperand_16,
                             L1_3_L2_4_G3_MINI_ALU_BoothOperand_15,
                             L1_3_L2_4_G3_MINI_ALU_BoothOperand_14,
                             L1_3_L2_4_G3_MINI_ALU_BoothOperand_13,
                             L1_3_L2_4_G3_MINI_ALU_BoothOperand_12,
                             L1_3_L2_4_G3_MINI_ALU_BoothOperand_11,
                             L1_3_L2_4_G3_MINI_ALU_BoothOperand_10,
                             L1_3_L2_4_G3_MINI_ALU_BoothOperand_9,
                             L1FirstOperands_12__16,L1FirstOperands_12__16,
                             L1FirstOperands_12__16,L1FirstOperands_12__16,
                             L1FirstOperands_12__16,L1FirstOperands_12__16,
                             L1FirstOperands_12__16,L1FirstOperands_12__16,
                             L1FirstOperands_12__16}), .BoothP ({
                             L1_3_L2_4_G3_MINI_ALU_BoothP_16,
                             L1_3_L2_4_G3_MINI_ALU_BoothP_15,
                             L1_3_L2_4_G3_MINI_ALU_BoothP_14,
                             L1_3_L2_4_G3_MINI_ALU_BoothP_13,
                             L1_3_L2_4_G3_MINI_ALU_BoothP_12,
                             L1_3_L2_4_G3_MINI_ALU_BoothP_11,
                             L1_3_L2_4_G3_MINI_ALU_BoothP_10,
                             L1_3_L2_4_G3_MINI_ALU_BoothP_9,
                             L1_3_L2_4_G3_MINI_ALU_BoothP_8,
                             L1_3_L2_4_G3_MINI_ALU_BoothP_7,
                             L1_3_L2_4_G3_MINI_ALU_BoothP_6,
                             L1_3_L2_4_G3_MINI_ALU_BoothP_5,
                             L1_3_L2_4_G3_MINI_ALU_BoothP_4,
                             L1_3_L2_4_G3_MINI_ALU_BoothP_3,
                             L1_3_L2_4_G3_MINI_ALU_BoothP_2,
                             L1_3_L2_4_G3_MINI_ALU_BoothP_1,
                             L1_3_L2_4_G3_MINI_ALU_BoothP_0}), .SelOperand (
                             nx3287), .Operation (
                             L1_3_L2_4_G3_MINI_ALU_BoothXORCheck), .AdderResult (
                             {L3ResultsLarge_0__16,L3ResultsLarge_0__15,
                             L3ResultsLarge_0__14,L3ResultsLarge_0__13,
                             L3ResultsLarge_0__12,L3ResultsLarge_0__11,
                             L3ResultsLarge_0__10,L3ResultsLarge_0__9,
                             L3ResultsLarge_0__8,L3ResultsLarge_0__7,
                             L3ResultsLarge_0__6,L3ResultsLarge_0__5,
                             L3ResultsLarge_0__4,L3ResultsLarge_0__3,
                             L3ResultsLarge_0__2,L3ResultsLarge_0__1,
                             L3ResultsLarge_0__0}), .AdderBoothResult ({
                             \$dummy [683],
                             L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_15,
                             L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_14,
                             L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_13,
                             L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_12,
                             L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_11,
                             L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_10,
                             L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_9,
                             L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_8,
                             L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_7,
                             L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_6,
                             L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_5,
                             L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_4,
                             L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_3,
                             L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_2,
                             L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_1,
                             L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_0})) ;
    booth_unit_17 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT (.CLK (CLK), .RST (RST), .Start (
                  Start), .Instr (Instr), .LoopingAndResultNotReady (nx3279), .Filter (
                  {FilterDin_3__4__7,FilterDin_3__4__6,FilterDin_3__4__5,
                  FilterDin_3__4__4,FilterDin_3__4__3,FilterDin_3__4__2,
                  FilterDin_3__4__1,FilterDin_3__4__0}), .Window ({
                  WindowDin_3__4__7,WindowDin_3__4__6,WindowDin_3__4__5,
                  WindowDin_3__4__4,WindowDin_3__4__3,WindowDin_3__4__2,
                  WindowDin_3__4__1,WindowDin_3__4__0}), .AdderBoothResult ({
                  L1FirstOperands_12__16,
                  L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_15,
                  L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_14,
                  L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_13,
                  L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_12,
                  L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_11,
                  L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_10,
                  L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_9,
                  L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_8,
                  L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_7,
                  L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_6,
                  L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_5,
                  L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_4,
                  L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_3,
                  L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_2,
                  L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_1,
                  L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_0}), .BoothXORCheck (
                  L1_3_L2_4_G3_MINI_ALU_BoothXORCheck), .BoothResult ({
                  \$dummy [684],\$dummy [685],\$dummy [686],\$dummy [687],
                  \$dummy [688],\$dummy [689],\$dummy [690],\$dummy [691]}), .BoothAddingOperand (
                  {L1_3_L2_4_G3_MINI_ALU_BoothOperand_16,
                  L1_3_L2_4_G3_MINI_ALU_BoothOperand_15,
                  L1_3_L2_4_G3_MINI_ALU_BoothOperand_14,
                  L1_3_L2_4_G3_MINI_ALU_BoothOperand_13,
                  L1_3_L2_4_G3_MINI_ALU_BoothOperand_12,
                  L1_3_L2_4_G3_MINI_ALU_BoothOperand_11,
                  L1_3_L2_4_G3_MINI_ALU_BoothOperand_10,
                  L1_3_L2_4_G3_MINI_ALU_BoothOperand_9,\$dummy [692],
                  \$dummy [693],\$dummy [694],\$dummy [695],\$dummy [696],
                  \$dummy [697],\$dummy [698],\$dummy [699],\$dummy [700]}), .BoothP (
                  {L1_3_L2_4_G3_MINI_ALU_BoothP_16,
                  L1_3_L2_4_G3_MINI_ALU_BoothP_15,
                  L1_3_L2_4_G3_MINI_ALU_BoothP_14,
                  L1_3_L2_4_G3_MINI_ALU_BoothP_13,
                  L1_3_L2_4_G3_MINI_ALU_BoothP_12,
                  L1_3_L2_4_G3_MINI_ALU_BoothP_11,
                  L1_3_L2_4_G3_MINI_ALU_BoothP_10,L1_3_L2_4_G3_MINI_ALU_BoothP_9
                  ,L1_3_L2_4_G3_MINI_ALU_BoothP_8,L1_3_L2_4_G3_MINI_ALU_BoothP_7
                  ,L1_3_L2_4_G3_MINI_ALU_BoothP_6,L1_3_L2_4_G3_MINI_ALU_BoothP_5
                  ,L1_3_L2_4_G3_MINI_ALU_BoothP_4,L1_3_L2_4_G3_MINI_ALU_BoothP_3
                  ,L1_3_L2_4_G3_MINI_ALU_BoothP_2,L1_3_L2_4_G3_MINI_ALU_BoothP_1
                  ,L1_3_L2_4_G3_MINI_ALU_BoothP_0}), .LargeWindowShifted ({
                  \$dummy [701],\$dummy [702],\$dummy [703],\$dummy [704],
                  \$dummy [705],\$dummy [706],\$dummy [707],\$dummy [708],
                  \$dummy [709],\$dummy [710],\$dummy [711],\$dummy [712],
                  \$dummy [713],\$dummy [714],\$dummy [715],\$dummy [716],
                  \$dummy [717]})) ;
    booth_adder_17_unfolded4 L1_4_L2_0_G3_MINI_ALU_BOOTH_ADDER (.AdderFirstOperand (
                             {L2ResultsLarge_2__16,L2ResultsLarge_2__15,
                             L2ResultsLarge_2__14,L2ResultsLarge_2__13,
                             L2ResultsLarge_2__12,L2ResultsLarge_2__11,
                             L2ResultsLarge_2__10,L2ResultsLarge_2__9,
                             L2ResultsLarge_2__8,L2ResultsLarge_2__7,
                             L2ResultsLarge_2__6,L2ResultsLarge_2__5,
                             L2ResultsLarge_2__4,L2ResultsLarge_2__3,
                             L2ResultsLarge_2__2,L2ResultsLarge_2__1,
                             L2ResultsLarge_2__0}), .AdderSecondOperand ({
                             L2ResultsLarge_3__16,L2ResultsLarge_3__15,
                             L2ResultsLarge_3__14,L2ResultsLarge_3__13,
                             L2ResultsLarge_3__12,L2ResultsLarge_3__11,
                             L2ResultsLarge_3__10,L2ResultsLarge_3__9,
                             L2ResultsLarge_3__8,L2ResultsLarge_3__7,
                             L2ResultsLarge_3__6,L2ResultsLarge_3__5,
                             L2ResultsLarge_3__4,L2ResultsLarge_3__3,
                             L2ResultsLarge_3__2,L2ResultsLarge_3__1,
                             L2ResultsLarge_3__0}), .BoothOperand ({
                             L1_4_L2_0_G3_MINI_ALU_BoothOperand_16,
                             L1_4_L2_0_G3_MINI_ALU_BoothOperand_15,
                             L1_4_L2_0_G3_MINI_ALU_BoothOperand_14,
                             L1_4_L2_0_G3_MINI_ALU_BoothOperand_13,
                             L1_4_L2_0_G3_MINI_ALU_BoothOperand_12,
                             L1_4_L2_0_G3_MINI_ALU_BoothOperand_11,
                             L1_4_L2_0_G3_MINI_ALU_BoothOperand_10,
                             L1_4_L2_0_G3_MINI_ALU_BoothOperand_9,
                             L1FirstOperands_12__16,L1FirstOperands_12__16,
                             L1FirstOperands_12__16,L1FirstOperands_12__16,
                             L1FirstOperands_12__16,L1FirstOperands_12__16,
                             L1FirstOperands_12__16,L1FirstOperands_12__16,
                             L1FirstOperands_12__16}), .BoothP ({
                             L1_4_L2_0_G3_MINI_ALU_BoothP_16,
                             L1_4_L2_0_G3_MINI_ALU_BoothP_15,
                             L1_4_L2_0_G3_MINI_ALU_BoothP_14,
                             L1_4_L2_0_G3_MINI_ALU_BoothP_13,
                             L1_4_L2_0_G3_MINI_ALU_BoothP_12,
                             L1_4_L2_0_G3_MINI_ALU_BoothP_11,
                             L1_4_L2_0_G3_MINI_ALU_BoothP_10,
                             L1_4_L2_0_G3_MINI_ALU_BoothP_9,
                             L1_4_L2_0_G3_MINI_ALU_BoothP_8,
                             L1_4_L2_0_G3_MINI_ALU_BoothP_7,
                             L1_4_L2_0_G3_MINI_ALU_BoothP_6,
                             L1_4_L2_0_G3_MINI_ALU_BoothP_5,
                             L1_4_L2_0_G3_MINI_ALU_BoothP_4,
                             L1_4_L2_0_G3_MINI_ALU_BoothP_3,
                             L1_4_L2_0_G3_MINI_ALU_BoothP_2,
                             L1_4_L2_0_G3_MINI_ALU_BoothP_1,
                             L1_4_L2_0_G3_MINI_ALU_BoothP_0}), .SelOperand (
                             nx3287), .Operation (
                             L1_4_L2_0_G3_MINI_ALU_BoothXORCheck), .AdderResult (
                             {L3ResultsLarge_1__16,L3ResultsLarge_1__15,
                             L3ResultsLarge_1__14,L3ResultsLarge_1__13,
                             L3ResultsLarge_1__12,L3ResultsLarge_1__11,
                             L3ResultsLarge_1__10,L3ResultsLarge_1__9,
                             L3ResultsLarge_1__8,L3ResultsLarge_1__7,
                             L3ResultsLarge_1__6,L3ResultsLarge_1__5,
                             L3ResultsLarge_1__4,L3ResultsLarge_1__3,
                             L3ResultsLarge_1__2,L3ResultsLarge_1__1,
                             L3ResultsLarge_1__0}), .AdderBoothResult ({
                             \$dummy [718],
                             L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_15,
                             L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_14,
                             L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_13,
                             L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_12,
                             L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_11,
                             L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_10,
                             L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_9,
                             L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_8,
                             L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_7,
                             L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_6,
                             L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_5,
                             L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_4,
                             L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_3,
                             L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_2,
                             L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_1,
                             L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_0})) ;
    booth_unit_17 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT (.CLK (CLK), .RST (RST), .Start (
                  Start), .Instr (Instr), .LoopingAndResultNotReady (nx3279), .Filter (
                  {FilterDin_4__0__7,FilterDin_4__0__6,FilterDin_4__0__5,
                  FilterDin_4__0__4,FilterDin_4__0__3,FilterDin_4__0__2,
                  FilterDin_4__0__1,FilterDin_4__0__0}), .Window ({
                  WindowDin_4__0__7,WindowDin_4__0__6,WindowDin_4__0__5,
                  WindowDin_4__0__4,WindowDin_4__0__3,WindowDin_4__0__2,
                  WindowDin_4__0__1,WindowDin_4__0__0}), .AdderBoothResult ({
                  L1FirstOperands_12__16,
                  L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_15,
                  L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_14,
                  L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_13,
                  L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_12,
                  L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_11,
                  L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_10,
                  L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_9,
                  L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_8,
                  L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_7,
                  L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_6,
                  L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_5,
                  L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_4,
                  L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_3,
                  L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_2,
                  L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_1,
                  L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_0}), .BoothXORCheck (
                  L1_4_L2_0_G3_MINI_ALU_BoothXORCheck), .BoothResult ({
                  \$dummy [719],\$dummy [720],\$dummy [721],\$dummy [722],
                  \$dummy [723],\$dummy [724],\$dummy [725],\$dummy [726]}), .BoothAddingOperand (
                  {L1_4_L2_0_G3_MINI_ALU_BoothOperand_16,
                  L1_4_L2_0_G3_MINI_ALU_BoothOperand_15,
                  L1_4_L2_0_G3_MINI_ALU_BoothOperand_14,
                  L1_4_L2_0_G3_MINI_ALU_BoothOperand_13,
                  L1_4_L2_0_G3_MINI_ALU_BoothOperand_12,
                  L1_4_L2_0_G3_MINI_ALU_BoothOperand_11,
                  L1_4_L2_0_G3_MINI_ALU_BoothOperand_10,
                  L1_4_L2_0_G3_MINI_ALU_BoothOperand_9,\$dummy [727],
                  \$dummy [728],\$dummy [729],\$dummy [730],\$dummy [731],
                  \$dummy [732],\$dummy [733],\$dummy [734],\$dummy [735]}), .BoothP (
                  {L1_4_L2_0_G3_MINI_ALU_BoothP_16,
                  L1_4_L2_0_G3_MINI_ALU_BoothP_15,
                  L1_4_L2_0_G3_MINI_ALU_BoothP_14,
                  L1_4_L2_0_G3_MINI_ALU_BoothP_13,
                  L1_4_L2_0_G3_MINI_ALU_BoothP_12,
                  L1_4_L2_0_G3_MINI_ALU_BoothP_11,
                  L1_4_L2_0_G3_MINI_ALU_BoothP_10,L1_4_L2_0_G3_MINI_ALU_BoothP_9
                  ,L1_4_L2_0_G3_MINI_ALU_BoothP_8,L1_4_L2_0_G3_MINI_ALU_BoothP_7
                  ,L1_4_L2_0_G3_MINI_ALU_BoothP_6,L1_4_L2_0_G3_MINI_ALU_BoothP_5
                  ,L1_4_L2_0_G3_MINI_ALU_BoothP_4,L1_4_L2_0_G3_MINI_ALU_BoothP_3
                  ,L1_4_L2_0_G3_MINI_ALU_BoothP_2,L1_4_L2_0_G3_MINI_ALU_BoothP_1
                  ,L1_4_L2_0_G3_MINI_ALU_BoothP_0}), .LargeWindowShifted ({
                  \$dummy [736],\$dummy [737],\$dummy [738],\$dummy [739],
                  \$dummy [740],\$dummy [741],\$dummy [742],\$dummy [743],
                  \$dummy [744],\$dummy [745],\$dummy [746],\$dummy [747],
                  \$dummy [748],\$dummy [749],\$dummy [750],\$dummy [751],
                  \$dummy [752]})) ;
    booth_adder_17_unfolded4 L1_4_L2_1_G3_MINI_ALU_BOOTH_ADDER (.AdderFirstOperand (
                             {L2ResultsLarge_4__16,L2ResultsLarge_4__15,
                             L2ResultsLarge_4__14,L2ResultsLarge_4__13,
                             L2ResultsLarge_4__12,L2ResultsLarge_4__11,
                             L2ResultsLarge_4__10,L2ResultsLarge_4__9,
                             L2ResultsLarge_4__8,L2ResultsLarge_4__7,
                             L2ResultsLarge_4__6,L2ResultsLarge_4__5,
                             L2ResultsLarge_4__4,L2ResultsLarge_4__3,
                             L2ResultsLarge_4__2,L2ResultsLarge_4__1,
                             L2ResultsLarge_4__0}), .AdderSecondOperand ({
                             L2ResultsLarge_5__16,L2ResultsLarge_5__15,
                             L2ResultsLarge_5__14,L2ResultsLarge_5__13,
                             L2ResultsLarge_5__12,L2ResultsLarge_5__11,
                             L2ResultsLarge_5__10,L2ResultsLarge_5__9,
                             L2ResultsLarge_5__8,L2ResultsLarge_5__7,
                             L2ResultsLarge_5__6,L2ResultsLarge_5__5,
                             L2ResultsLarge_5__4,L2ResultsLarge_5__3,
                             L2ResultsLarge_5__2,L2ResultsLarge_5__1,
                             L2ResultsLarge_5__0}), .BoothOperand ({
                             L1_4_L2_1_G3_MINI_ALU_BoothOperand_16,
                             L1_4_L2_1_G3_MINI_ALU_BoothOperand_15,
                             L1_4_L2_1_G3_MINI_ALU_BoothOperand_14,
                             L1_4_L2_1_G3_MINI_ALU_BoothOperand_13,
                             L1_4_L2_1_G3_MINI_ALU_BoothOperand_12,
                             L1_4_L2_1_G3_MINI_ALU_BoothOperand_11,
                             L1_4_L2_1_G3_MINI_ALU_BoothOperand_10,
                             L1_4_L2_1_G3_MINI_ALU_BoothOperand_9,
                             L1FirstOperands_12__16,L1FirstOperands_12__16,
                             L1FirstOperands_12__16,L1FirstOperands_12__16,
                             L1FirstOperands_12__16,L1FirstOperands_12__16,
                             L1FirstOperands_12__16,L1FirstOperands_12__16,
                             L1FirstOperands_12__16}), .BoothP ({
                             L1_4_L2_1_G3_MINI_ALU_BoothP_16,
                             L1_4_L2_1_G3_MINI_ALU_BoothP_15,
                             L1_4_L2_1_G3_MINI_ALU_BoothP_14,
                             L1_4_L2_1_G3_MINI_ALU_BoothP_13,
                             L1_4_L2_1_G3_MINI_ALU_BoothP_12,
                             L1_4_L2_1_G3_MINI_ALU_BoothP_11,
                             L1_4_L2_1_G3_MINI_ALU_BoothP_10,
                             L1_4_L2_1_G3_MINI_ALU_BoothP_9,
                             L1_4_L2_1_G3_MINI_ALU_BoothP_8,
                             L1_4_L2_1_G3_MINI_ALU_BoothP_7,
                             L1_4_L2_1_G3_MINI_ALU_BoothP_6,
                             L1_4_L2_1_G3_MINI_ALU_BoothP_5,
                             L1_4_L2_1_G3_MINI_ALU_BoothP_4,
                             L1_4_L2_1_G3_MINI_ALU_BoothP_3,
                             L1_4_L2_1_G3_MINI_ALU_BoothP_2,
                             L1_4_L2_1_G3_MINI_ALU_BoothP_1,
                             L1_4_L2_1_G3_MINI_ALU_BoothP_0}), .SelOperand (
                             nx3289), .Operation (
                             L1_4_L2_1_G3_MINI_ALU_BoothXORCheck), .AdderResult (
                             {L3ResultsLarge_2__16,L3ResultsLarge_2__15,
                             L3ResultsLarge_2__14,L3ResultsLarge_2__13,
                             L3ResultsLarge_2__12,L3ResultsLarge_2__11,
                             L3ResultsLarge_2__10,L3ResultsLarge_2__9,
                             L3ResultsLarge_2__8,L3ResultsLarge_2__7,
                             L3ResultsLarge_2__6,L3ResultsLarge_2__5,
                             L3ResultsLarge_2__4,L3ResultsLarge_2__3,
                             L3ResultsLarge_2__2,L3ResultsLarge_2__1,
                             L3ResultsLarge_2__0}), .AdderBoothResult ({
                             \$dummy [753],
                             L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_15,
                             L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_14,
                             L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_13,
                             L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_12,
                             L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_11,
                             L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_10,
                             L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_9,
                             L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_8,
                             L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_7,
                             L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_6,
                             L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_5,
                             L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_4,
                             L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_3,
                             L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_2,
                             L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_1,
                             L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_0})) ;
    booth_unit_17 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT (.CLK (CLK), .RST (RST), .Start (
                  Start), .Instr (Instr), .LoopingAndResultNotReady (nx3281), .Filter (
                  {FilterDin_4__1__7,FilterDin_4__1__6,FilterDin_4__1__5,
                  FilterDin_4__1__4,FilterDin_4__1__3,FilterDin_4__1__2,
                  FilterDin_4__1__1,FilterDin_4__1__0}), .Window ({
                  WindowDin_4__1__7,WindowDin_4__1__6,WindowDin_4__1__5,
                  WindowDin_4__1__4,WindowDin_4__1__3,WindowDin_4__1__2,
                  WindowDin_4__1__1,WindowDin_4__1__0}), .AdderBoothResult ({
                  L1FirstOperands_12__16,
                  L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_15,
                  L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_14,
                  L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_13,
                  L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_12,
                  L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_11,
                  L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_10,
                  L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_9,
                  L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_8,
                  L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_7,
                  L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_6,
                  L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_5,
                  L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_4,
                  L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_3,
                  L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_2,
                  L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_1,
                  L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_0}), .BoothXORCheck (
                  L1_4_L2_1_G3_MINI_ALU_BoothXORCheck), .BoothResult ({
                  \$dummy [754],\$dummy [755],\$dummy [756],\$dummy [757],
                  \$dummy [758],\$dummy [759],\$dummy [760],\$dummy [761]}), .BoothAddingOperand (
                  {L1_4_L2_1_G3_MINI_ALU_BoothOperand_16,
                  L1_4_L2_1_G3_MINI_ALU_BoothOperand_15,
                  L1_4_L2_1_G3_MINI_ALU_BoothOperand_14,
                  L1_4_L2_1_G3_MINI_ALU_BoothOperand_13,
                  L1_4_L2_1_G3_MINI_ALU_BoothOperand_12,
                  L1_4_L2_1_G3_MINI_ALU_BoothOperand_11,
                  L1_4_L2_1_G3_MINI_ALU_BoothOperand_10,
                  L1_4_L2_1_G3_MINI_ALU_BoothOperand_9,\$dummy [762],
                  \$dummy [763],\$dummy [764],\$dummy [765],\$dummy [766],
                  \$dummy [767],\$dummy [768],\$dummy [769],\$dummy [770]}), .BoothP (
                  {L1_4_L2_1_G3_MINI_ALU_BoothP_16,
                  L1_4_L2_1_G3_MINI_ALU_BoothP_15,
                  L1_4_L2_1_G3_MINI_ALU_BoothP_14,
                  L1_4_L2_1_G3_MINI_ALU_BoothP_13,
                  L1_4_L2_1_G3_MINI_ALU_BoothP_12,
                  L1_4_L2_1_G3_MINI_ALU_BoothP_11,
                  L1_4_L2_1_G3_MINI_ALU_BoothP_10,L1_4_L2_1_G3_MINI_ALU_BoothP_9
                  ,L1_4_L2_1_G3_MINI_ALU_BoothP_8,L1_4_L2_1_G3_MINI_ALU_BoothP_7
                  ,L1_4_L2_1_G3_MINI_ALU_BoothP_6,L1_4_L2_1_G3_MINI_ALU_BoothP_5
                  ,L1_4_L2_1_G3_MINI_ALU_BoothP_4,L1_4_L2_1_G3_MINI_ALU_BoothP_3
                  ,L1_4_L2_1_G3_MINI_ALU_BoothP_2,L1_4_L2_1_G3_MINI_ALU_BoothP_1
                  ,L1_4_L2_1_G3_MINI_ALU_BoothP_0}), .LargeWindowShifted ({
                  \$dummy [771],\$dummy [772],\$dummy [773],\$dummy [774],
                  \$dummy [775],\$dummy [776],\$dummy [777],\$dummy [778],
                  \$dummy [779],\$dummy [780],\$dummy [781],\$dummy [782],
                  \$dummy [783],\$dummy [784],\$dummy [785],\$dummy [786],
                  \$dummy [787]})) ;
    booth_adder_17_unfolded4 L1_4_L2_2_G4_MINI_ALU_BOOTH_ADDER (.AdderFirstOperand (
                             {L3ResultsLarge_0__16,L3ResultsLarge_0__15,
                             L3ResultsLarge_0__14,L3ResultsLarge_0__13,
                             L3ResultsLarge_0__12,L3ResultsLarge_0__11,
                             L3ResultsLarge_0__10,L3ResultsLarge_0__9,
                             L3ResultsLarge_0__8,L3ResultsLarge_0__7,
                             L3ResultsLarge_0__6,L3ResultsLarge_0__5,
                             L3ResultsLarge_0__4,L3ResultsLarge_0__3,
                             L3ResultsLarge_0__2,L3ResultsLarge_0__1,
                             L3ResultsLarge_0__0}), .AdderSecondOperand ({
                             L3ResultsLarge_1__16,L3ResultsLarge_1__15,
                             L3ResultsLarge_1__14,L3ResultsLarge_1__13,
                             L3ResultsLarge_1__12,L3ResultsLarge_1__11,
                             L3ResultsLarge_1__10,L3ResultsLarge_1__9,
                             L3ResultsLarge_1__8,L3ResultsLarge_1__7,
                             L3ResultsLarge_1__6,L3ResultsLarge_1__5,
                             L3ResultsLarge_1__4,L3ResultsLarge_1__3,
                             L3ResultsLarge_1__2,L3ResultsLarge_1__1,
                             L3ResultsLarge_1__0}), .BoothOperand ({
                             L1_4_L2_2_G4_MINI_ALU_BoothOperand_16,
                             L1_4_L2_2_G4_MINI_ALU_BoothOperand_15,
                             L1_4_L2_2_G4_MINI_ALU_BoothOperand_14,
                             L1_4_L2_2_G4_MINI_ALU_BoothOperand_13,
                             L1_4_L2_2_G4_MINI_ALU_BoothOperand_12,
                             L1_4_L2_2_G4_MINI_ALU_BoothOperand_11,
                             L1_4_L2_2_G4_MINI_ALU_BoothOperand_10,
                             L1_4_L2_2_G4_MINI_ALU_BoothOperand_9,
                             L1FirstOperands_12__16,L1FirstOperands_12__16,
                             L1FirstOperands_12__16,L1FirstOperands_12__16,
                             L1FirstOperands_12__16,L1FirstOperands_12__16,
                             L1FirstOperands_12__16,L1FirstOperands_12__16,
                             L1FirstOperands_12__16}), .BoothP ({
                             L1_4_L2_2_G4_MINI_ALU_BoothP_16,
                             L1_4_L2_2_G4_MINI_ALU_BoothP_15,
                             L1_4_L2_2_G4_MINI_ALU_BoothP_14,
                             L1_4_L2_2_G4_MINI_ALU_BoothP_13,
                             L1_4_L2_2_G4_MINI_ALU_BoothP_12,
                             L1_4_L2_2_G4_MINI_ALU_BoothP_11,
                             L1_4_L2_2_G4_MINI_ALU_BoothP_10,
                             L1_4_L2_2_G4_MINI_ALU_BoothP_9,
                             L1_4_L2_2_G4_MINI_ALU_BoothP_8,
                             L1_4_L2_2_G4_MINI_ALU_BoothP_7,
                             L1_4_L2_2_G4_MINI_ALU_BoothP_6,
                             L1_4_L2_2_G4_MINI_ALU_BoothP_5,
                             L1_4_L2_2_G4_MINI_ALU_BoothP_4,
                             L1_4_L2_2_G4_MINI_ALU_BoothP_3,
                             L1_4_L2_2_G4_MINI_ALU_BoothP_2,
                             L1_4_L2_2_G4_MINI_ALU_BoothP_1,
                             L1_4_L2_2_G4_MINI_ALU_BoothP_0}), .SelOperand (
                             nx3289), .Operation (
                             L1_4_L2_2_G4_MINI_ALU_BoothXORCheck), .AdderResult (
                             {L4ResultsLarge_0__16,L4ResultsLarge_0__15,
                             L4ResultsLarge_0__14,L4ResultsLarge_0__13,
                             L4ResultsLarge_0__12,L4ResultsLarge_0__11,
                             L4ResultsLarge_0__10,L4ResultsLarge_0__9,
                             L4ResultsLarge_0__8,L4ResultsLarge_0__7,
                             L4ResultsLarge_0__6,L4ResultsLarge_0__5,
                             L4ResultsLarge_0__4,L4ResultsLarge_0__3,
                             L4ResultsLarge_0__2,L4ResultsLarge_0__1,
                             L4ResultsLarge_0__0}), .AdderBoothResult ({
                             \$dummy [788],
                             L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_15,
                             L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_14,
                             L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_13,
                             L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_12,
                             L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_11,
                             L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_10,
                             L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_9,
                             L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_8,
                             L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_7,
                             L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_6,
                             L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_5,
                             L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_4,
                             L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_3,
                             L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_2,
                             L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_1,
                             L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_0})) ;
    booth_unit_17 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT (.CLK (CLK), .RST (RST), .Start (
                  Start), .Instr (Instr), .LoopingAndResultNotReady (nx3281), .Filter (
                  {FilterDin_4__2__7,FilterDin_4__2__6,FilterDin_4__2__5,
                  FilterDin_4__2__4,FilterDin_4__2__3,FilterDin_4__2__2,
                  FilterDin_4__2__1,FilterDin_4__2__0}), .Window ({
                  WindowDin_4__2__7,WindowDin_4__2__6,WindowDin_4__2__5,
                  WindowDin_4__2__4,WindowDin_4__2__3,WindowDin_4__2__2,
                  WindowDin_4__2__1,WindowDin_4__2__0}), .AdderBoothResult ({
                  L1FirstOperands_12__16,
                  L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_15,
                  L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_14,
                  L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_13,
                  L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_12,
                  L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_11,
                  L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_10,
                  L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_9,
                  L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_8,
                  L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_7,
                  L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_6,
                  L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_5,
                  L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_4,
                  L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_3,
                  L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_2,
                  L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_1,
                  L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_0}), .BoothXORCheck (
                  L1_4_L2_2_G4_MINI_ALU_BoothXORCheck), .BoothResult ({
                  \$dummy [789],\$dummy [790],\$dummy [791],\$dummy [792],
                  \$dummy [793],\$dummy [794],\$dummy [795],\$dummy [796]}), .BoothAddingOperand (
                  {L1_4_L2_2_G4_MINI_ALU_BoothOperand_16,
                  L1_4_L2_2_G4_MINI_ALU_BoothOperand_15,
                  L1_4_L2_2_G4_MINI_ALU_BoothOperand_14,
                  L1_4_L2_2_G4_MINI_ALU_BoothOperand_13,
                  L1_4_L2_2_G4_MINI_ALU_BoothOperand_12,
                  L1_4_L2_2_G4_MINI_ALU_BoothOperand_11,
                  L1_4_L2_2_G4_MINI_ALU_BoothOperand_10,
                  L1_4_L2_2_G4_MINI_ALU_BoothOperand_9,\$dummy [797],
                  \$dummy [798],\$dummy [799],\$dummy [800],\$dummy [801],
                  \$dummy [802],\$dummy [803],\$dummy [804],\$dummy [805]}), .BoothP (
                  {L1_4_L2_2_G4_MINI_ALU_BoothP_16,
                  L1_4_L2_2_G4_MINI_ALU_BoothP_15,
                  L1_4_L2_2_G4_MINI_ALU_BoothP_14,
                  L1_4_L2_2_G4_MINI_ALU_BoothP_13,
                  L1_4_L2_2_G4_MINI_ALU_BoothP_12,
                  L1_4_L2_2_G4_MINI_ALU_BoothP_11,
                  L1_4_L2_2_G4_MINI_ALU_BoothP_10,L1_4_L2_2_G4_MINI_ALU_BoothP_9
                  ,L1_4_L2_2_G4_MINI_ALU_BoothP_8,L1_4_L2_2_G4_MINI_ALU_BoothP_7
                  ,L1_4_L2_2_G4_MINI_ALU_BoothP_6,L1_4_L2_2_G4_MINI_ALU_BoothP_5
                  ,L1_4_L2_2_G4_MINI_ALU_BoothP_4,L1_4_L2_2_G4_MINI_ALU_BoothP_3
                  ,L1_4_L2_2_G4_MINI_ALU_BoothP_2,L1_4_L2_2_G4_MINI_ALU_BoothP_1
                  ,L1_4_L2_2_G4_MINI_ALU_BoothP_0}), .LargeWindowShifted ({
                  \$dummy [806],\$dummy [807],\$dummy [808],\$dummy [809],
                  \$dummy [810],\$dummy [811],\$dummy [812],\$dummy [813],
                  \$dummy [814],\$dummy [815],\$dummy [816],\$dummy [817],
                  \$dummy [818],\$dummy [819],\$dummy [820],\$dummy [821],
                  \$dummy [822]})) ;
    booth_adder_17_unfolded4 L1_4_L2_3_G5_MINI_ALU_BOOTH_ADDER (.AdderFirstOperand (
                             {L4ResultsLarge_0__16,L4ResultsLarge_0__15,
                             L4ResultsLarge_0__14,L4ResultsLarge_0__13,
                             L4ResultsLarge_0__12,L4ResultsLarge_0__11,
                             L4ResultsLarge_0__10,L4ResultsLarge_0__9,
                             L4ResultsLarge_0__8,L4ResultsLarge_0__7,
                             L4ResultsLarge_0__6,L4ResultsLarge_0__5,
                             L4ResultsLarge_0__4,L4ResultsLarge_0__3,
                             L4ResultsLarge_0__2,L4ResultsLarge_0__1,
                             L4ResultsLarge_0__0}), .AdderSecondOperand ({
                             L3ResultsLarge_2__16,L3ResultsLarge_2__15,
                             L3ResultsLarge_2__14,L3ResultsLarge_2__13,
                             L3ResultsLarge_2__12,L3ResultsLarge_2__11,
                             L3ResultsLarge_2__10,L3ResultsLarge_2__9,
                             L3ResultsLarge_2__8,L3ResultsLarge_2__7,
                             L3ResultsLarge_2__6,L3ResultsLarge_2__5,
                             L3ResultsLarge_2__4,L3ResultsLarge_2__3,
                             L3ResultsLarge_2__2,L3ResultsLarge_2__1,
                             L3ResultsLarge_2__0}), .BoothOperand ({
                             L1_4_L2_3_G5_MINI_ALU_BoothOperand_16,
                             L1_4_L2_3_G5_MINI_ALU_BoothOperand_15,
                             L1_4_L2_3_G5_MINI_ALU_BoothOperand_14,
                             L1_4_L2_3_G5_MINI_ALU_BoothOperand_13,
                             L1_4_L2_3_G5_MINI_ALU_BoothOperand_12,
                             L1_4_L2_3_G5_MINI_ALU_BoothOperand_11,
                             L1_4_L2_3_G5_MINI_ALU_BoothOperand_10,
                             L1_4_L2_3_G5_MINI_ALU_BoothOperand_9,
                             L1FirstOperands_12__16,L1FirstOperands_12__16,
                             L1FirstOperands_12__16,L1FirstOperands_12__16,
                             L1FirstOperands_12__16,L1FirstOperands_12__16,
                             L1FirstOperands_12__16,L1FirstOperands_12__16,
                             L1FirstOperands_12__16}), .BoothP ({
                             L1_4_L2_3_G5_MINI_ALU_BoothP_16,
                             L1_4_L2_3_G5_MINI_ALU_BoothP_15,
                             L1_4_L2_3_G5_MINI_ALU_BoothP_14,
                             L1_4_L2_3_G5_MINI_ALU_BoothP_13,
                             L1_4_L2_3_G5_MINI_ALU_BoothP_12,
                             L1_4_L2_3_G5_MINI_ALU_BoothP_11,
                             L1_4_L2_3_G5_MINI_ALU_BoothP_10,
                             L1_4_L2_3_G5_MINI_ALU_BoothP_9,
                             L1_4_L2_3_G5_MINI_ALU_BoothP_8,
                             L1_4_L2_3_G5_MINI_ALU_BoothP_7,
                             L1_4_L2_3_G5_MINI_ALU_BoothP_6,
                             L1_4_L2_3_G5_MINI_ALU_BoothP_5,
                             L1_4_L2_3_G5_MINI_ALU_BoothP_4,
                             L1_4_L2_3_G5_MINI_ALU_BoothP_3,
                             L1_4_L2_3_G5_MINI_ALU_BoothP_2,
                             L1_4_L2_3_G5_MINI_ALU_BoothP_1,
                             L1_4_L2_3_G5_MINI_ALU_BoothP_0}), .SelOperand (
                             nx3289), .Operation (
                             L1_4_L2_3_G5_MINI_ALU_BoothXORCheck), .AdderResult (
                             {L5FirstOperands_1__16,L5FirstOperands_1__15,
                             L5FirstOperands_1__14,L5FirstOperands_1__13,
                             L5FirstOperands_1__12,L5FirstOperands_1__11,
                             L5FirstOperands_1__10,L5FirstOperands_1__9,
                             L5FirstOperands_1__8,L5FirstOperands_1__7,
                             L5FirstOperands_1__6,L5FirstOperands_1__5,
                             L5FirstOperands_1__4,L5FirstOperands_1__3,
                             L5FirstOperands_1__2,L5FirstOperands_1__1,
                             L5FirstOperands_1__0}), .AdderBoothResult ({
                             \$dummy [823],
                             L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_15,
                             L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_14,
                             L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_13,
                             L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_12,
                             L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_11,
                             L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_10,
                             L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_9,
                             L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_8,
                             L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_7,
                             L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_6,
                             L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_5,
                             L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_4,
                             L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_3,
                             L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_2,
                             L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_1,
                             L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_0})) ;
    booth_unit_17 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT (.CLK (CLK), .RST (RST), .Start (
                  Start), .Instr (Instr), .LoopingAndResultNotReady (nx3281), .Filter (
                  {FilterDin_4__3__7,FilterDin_4__3__6,FilterDin_4__3__5,
                  FilterDin_4__3__4,FilterDin_4__3__3,FilterDin_4__3__2,
                  FilterDin_4__3__1,FilterDin_4__3__0}), .Window ({
                  WindowDin_4__3__7,WindowDin_4__3__6,WindowDin_4__3__5,
                  WindowDin_4__3__4,WindowDin_4__3__3,WindowDin_4__3__2,
                  WindowDin_4__3__1,WindowDin_4__3__0}), .AdderBoothResult ({
                  L1FirstOperands_12__16,
                  L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_15,
                  L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_14,
                  L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_13,
                  L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_12,
                  L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_11,
                  L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_10,
                  L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_9,
                  L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_8,
                  L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_7,
                  L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_6,
                  L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_5,
                  L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_4,
                  L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_3,
                  L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_2,
                  L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_1,
                  L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_0}), .BoothXORCheck (
                  L1_4_L2_3_G5_MINI_ALU_BoothXORCheck), .BoothResult ({
                  \$dummy [824],\$dummy [825],\$dummy [826],\$dummy [827],
                  \$dummy [828],\$dummy [829],\$dummy [830],\$dummy [831]}), .BoothAddingOperand (
                  {L1_4_L2_3_G5_MINI_ALU_BoothOperand_16,
                  L1_4_L2_3_G5_MINI_ALU_BoothOperand_15,
                  L1_4_L2_3_G5_MINI_ALU_BoothOperand_14,
                  L1_4_L2_3_G5_MINI_ALU_BoothOperand_13,
                  L1_4_L2_3_G5_MINI_ALU_BoothOperand_12,
                  L1_4_L2_3_G5_MINI_ALU_BoothOperand_11,
                  L1_4_L2_3_G5_MINI_ALU_BoothOperand_10,
                  L1_4_L2_3_G5_MINI_ALU_BoothOperand_9,\$dummy [832],
                  \$dummy [833],\$dummy [834],\$dummy [835],\$dummy [836],
                  \$dummy [837],\$dummy [838],\$dummy [839],\$dummy [840]}), .BoothP (
                  {L1_4_L2_3_G5_MINI_ALU_BoothP_16,
                  L1_4_L2_3_G5_MINI_ALU_BoothP_15,
                  L1_4_L2_3_G5_MINI_ALU_BoothP_14,
                  L1_4_L2_3_G5_MINI_ALU_BoothP_13,
                  L1_4_L2_3_G5_MINI_ALU_BoothP_12,
                  L1_4_L2_3_G5_MINI_ALU_BoothP_11,
                  L1_4_L2_3_G5_MINI_ALU_BoothP_10,L1_4_L2_3_G5_MINI_ALU_BoothP_9
                  ,L1_4_L2_3_G5_MINI_ALU_BoothP_8,L1_4_L2_3_G5_MINI_ALU_BoothP_7
                  ,L1_4_L2_3_G5_MINI_ALU_BoothP_6,L1_4_L2_3_G5_MINI_ALU_BoothP_5
                  ,L1_4_L2_3_G5_MINI_ALU_BoothP_4,L1_4_L2_3_G5_MINI_ALU_BoothP_3
                  ,L1_4_L2_3_G5_MINI_ALU_BoothP_2,L1_4_L2_3_G5_MINI_ALU_BoothP_1
                  ,L1_4_L2_3_G5_MINI_ALU_BoothP_0}), .LargeWindowShifted ({
                  \$dummy [841],\$dummy [842],\$dummy [843],\$dummy [844],
                  \$dummy [845],\$dummy [846],\$dummy [847],\$dummy [848],
                  \$dummy [849],\$dummy [850],\$dummy [851],\$dummy [852],
                  \$dummy [853],\$dummy [854],\$dummy [855],\$dummy [856],
                  \$dummy [857]})) ;
    booth_adder_17_unfolded5 L1_4_L2_4_G5_MINI_ALU_BOOTH_ADDER (.AdderFirstOperand (
                             {L5FirstOperands_1__16,L5FirstOperands_1__15,
                             L5FirstOperands_1__14,L5FirstOperands_1__13,
                             L5FirstOperands_1__12,L5FirstOperands_1__11,
                             L5FirstOperands_1__10,L5FirstOperands_1__9,
                             L5FirstOperands_1__8,L5FirstOperands_1__7,
                             L5FirstOperands_1__6,L5FirstOperands_1__5,
                             L5FirstOperands_1__4,L5FirstOperands_1__3,
                             L5FirstOperands_1__2,L5FirstOperands_1__1,
                             L5FirstOperands_1__0}), .AdderSecondOperand ({
                             L1FirstOperands_12__16,
                             L1_4_L2_4_G5_MINI_ALU_OperationResult_15,
                             L1_4_L2_4_G5_MINI_ALU_OperationResult_14,
                             L1_4_L2_4_G5_MINI_ALU_OperationResult_13,
                             L1_4_L2_4_G5_MINI_ALU_OperationResult_12,
                             L1_4_L2_4_G5_MINI_ALU_OperationResult_11,
                             L1_4_L2_4_G5_MINI_ALU_OperationResult_10,
                             L1_4_L2_4_G5_MINI_ALU_OperationResult_9,
                             L1_4_L2_4_G5_MINI_ALU_OperationResult_8,
                             L1_4_L2_4_G5_MINI_ALU_OperationResult_7,
                             L1_4_L2_4_G5_MINI_ALU_OperationResult_6,
                             L1_4_L2_4_G5_MINI_ALU_OperationResult_5,
                             L1_4_L2_4_G5_MINI_ALU_OperationResult_4,
                             L1_4_L2_4_G5_MINI_ALU_OperationResult_3,
                             L1_4_L2_4_G5_MINI_ALU_OperationResult_2,
                             L1_4_L2_4_G5_MINI_ALU_OperationResult_1,
                             L1_4_L2_4_G5_MINI_ALU_OperationResult_0}), .BoothOperand (
                             {L1_4_L2_4_G5_MINI_ALU_BoothOperand_16,
                             L1_4_L2_4_G5_MINI_ALU_BoothOperand_15,
                             L1_4_L2_4_G5_MINI_ALU_BoothOperand_14,
                             L1_4_L2_4_G5_MINI_ALU_BoothOperand_13,
                             L1_4_L2_4_G5_MINI_ALU_BoothOperand_12,
                             L1_4_L2_4_G5_MINI_ALU_BoothOperand_11,
                             L1_4_L2_4_G5_MINI_ALU_BoothOperand_10,
                             L1_4_L2_4_G5_MINI_ALU_BoothOperand_9,
                             L1FirstOperands_12__16,L1FirstOperands_12__16,
                             L1FirstOperands_12__16,L1FirstOperands_12__16,
                             L1FirstOperands_12__16,L1FirstOperands_12__16,
                             L1FirstOperands_12__16,L1FirstOperands_12__16,
                             L1FirstOperands_12__16}), .BoothP ({
                             L1_4_L2_4_G5_MINI_ALU_BoothP_16,
                             L1_4_L2_4_G5_MINI_ALU_BoothP_15,
                             L1_4_L2_4_G5_MINI_ALU_BoothP_14,
                             L1_4_L2_4_G5_MINI_ALU_BoothP_13,
                             L1_4_L2_4_G5_MINI_ALU_BoothP_12,
                             L1_4_L2_4_G5_MINI_ALU_BoothP_11,
                             L1_4_L2_4_G5_MINI_ALU_BoothP_10,
                             L1_4_L2_4_G5_MINI_ALU_BoothP_9,
                             L1_4_L2_4_G5_MINI_ALU_BoothP_8,
                             L1_4_L2_4_G5_MINI_ALU_BoothP_7,
                             L1_4_L2_4_G5_MINI_ALU_BoothP_6,
                             L1_4_L2_4_G5_MINI_ALU_BoothP_5,
                             L1_4_L2_4_G5_MINI_ALU_BoothP_4,
                             L1_4_L2_4_G5_MINI_ALU_BoothP_3,
                             L1_4_L2_4_G5_MINI_ALU_BoothP_2,
                             L1_4_L2_4_G5_MINI_ALU_BoothP_1,
                             L1_4_L2_4_G5_MINI_ALU_BoothP_0}), .SelOperand (
                             nx3289), .Operation (
                             L1_4_L2_4_G5_MINI_ALU_BoothXORCheck), .AdderResult (
                             {\$dummy [858],\$dummy [859],\$dummy [860],
                             \$dummy [861],\$dummy [862],\$dummy [863],
                             \$dummy [864],\$dummy [865],\$dummy [866],
                             L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_7,
                             L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_6,
                             L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_5,
                             L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_4,
                             L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_3,
                             L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_2,
                             L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_1,
                             L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_0}), .AdderBoothResult (
                             {\$dummy [867],
                             L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_15,
                             L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_14,
                             L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_13,
                             L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_12,
                             L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_11,
                             L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_10,
                             L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_9,
                             L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_8,
                             L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_7,
                             L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_6,
                             L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_5,
                             L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_4,
                             L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_3,
                             L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_2,
                             L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_1,
                             L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_0})) ;
    booth_unit_17 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT (.CLK (CLK), .RST (RST), .Start (
                  Start), .Instr (Instr), .LoopingAndResultNotReady (nx3281), .Filter (
                  {FilterDin_4__4__7,FilterDin_4__4__6,FilterDin_4__4__5,
                  FilterDin_4__4__4,FilterDin_4__4__3,FilterDin_4__4__2,
                  FilterDin_4__4__1,FilterDin_4__4__0}), .Window ({
                  WindowDin_4__4__7,WindowDin_4__4__6,WindowDin_4__4__5,
                  WindowDin_4__4__4,WindowDin_4__4__3,WindowDin_4__4__2,
                  WindowDin_4__4__1,WindowDin_4__4__0}), .AdderBoothResult ({
                  L1FirstOperands_12__16,
                  L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_15,
                  L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_14,
                  L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_13,
                  L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_12,
                  L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_11,
                  L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_10,
                  L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_9,
                  L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_8,
                  L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_7,
                  L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_6,
                  L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_5,
                  L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_4,
                  L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_3,
                  L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_2,
                  L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_1,
                  L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_0}), .BoothXORCheck (
                  L1_4_L2_4_G5_MINI_ALU_BoothXORCheck), .BoothResult ({
                  \$dummy [868],\$dummy [869],\$dummy [870],\$dummy [871],
                  \$dummy [872],\$dummy [873],\$dummy [874],\$dummy [875]}), .BoothAddingOperand (
                  {L1_4_L2_4_G5_MINI_ALU_BoothOperand_16,
                  L1_4_L2_4_G5_MINI_ALU_BoothOperand_15,
                  L1_4_L2_4_G5_MINI_ALU_BoothOperand_14,
                  L1_4_L2_4_G5_MINI_ALU_BoothOperand_13,
                  L1_4_L2_4_G5_MINI_ALU_BoothOperand_12,
                  L1_4_L2_4_G5_MINI_ALU_BoothOperand_11,
                  L1_4_L2_4_G5_MINI_ALU_BoothOperand_10,
                  L1_4_L2_4_G5_MINI_ALU_BoothOperand_9,\$dummy [876],
                  \$dummy [877],\$dummy [878],\$dummy [879],\$dummy [880],
                  \$dummy [881],\$dummy [882],\$dummy [883],\$dummy [884]}), .BoothP (
                  {L1_4_L2_4_G5_MINI_ALU_BoothP_16,
                  L1_4_L2_4_G5_MINI_ALU_BoothP_15,
                  L1_4_L2_4_G5_MINI_ALU_BoothP_14,
                  L1_4_L2_4_G5_MINI_ALU_BoothP_13,
                  L1_4_L2_4_G5_MINI_ALU_BoothP_12,
                  L1_4_L2_4_G5_MINI_ALU_BoothP_11,
                  L1_4_L2_4_G5_MINI_ALU_BoothP_10,L1_4_L2_4_G5_MINI_ALU_BoothP_9
                  ,L1_4_L2_4_G5_MINI_ALU_BoothP_8,L1_4_L2_4_G5_MINI_ALU_BoothP_7
                  ,L1_4_L2_4_G5_MINI_ALU_BoothP_6,L1_4_L2_4_G5_MINI_ALU_BoothP_5
                  ,L1_4_L2_4_G5_MINI_ALU_BoothP_4,L1_4_L2_4_G5_MINI_ALU_BoothP_3
                  ,L1_4_L2_4_G5_MINI_ALU_BoothP_2,L1_4_L2_4_G5_MINI_ALU_BoothP_1
                  ,L1_4_L2_4_G5_MINI_ALU_BoothP_0}), .LargeWindowShifted ({
                  \$dummy [885],\$dummy [886],\$dummy [887],\$dummy [888],
                  \$dummy [889],\$dummy [890],\$dummy [891],\$dummy [892],
                  \$dummy [893],\$dummy [894],\$dummy [895],\$dummy [896],
                  \$dummy [897],\$dummy [898],\$dummy [899],\$dummy [900],
                  \$dummy [901]})) ;
    nor02ii ix2855 (.Y (NOT__13497), .A0 (Instr), .A1 (nx2856)) ;
    nand03 ix2857 (.Y (nx2856), .A0 (CounterOut_0), .A1 (CounterOut_3), .A2 (
           nx2876)) ;
    or02 ix1037 (.Y (nx1036), .A0 (Start), .A1 (RST)) ;
    xnor2 ix1067 (.Y (nx1066), .A0 (CounterOut_3), .A1 (nx2868)) ;
    nand03 ix2869 (.Y (nx2868), .A0 (CounterOut_2), .A1 (CounterOut_1), .A2 (
           CounterOut_0)) ;
    xnor2 ix1059 (.Y (nx1058), .A0 (CounterOut_2), .A1 (nx2872)) ;
    fake_gnd ix2305 (.Y (L1FirstOperands_12__16)) ;
    mux21_ni ix109 (.Y (L1_4_L2_4_G5_MINI_ALU_OperationResult_0), .A0 (
             L1_4_L2_4_G5_MINI_ALU_BoothP_1), .A1 (WindowDin_4__4__0), .S0 (
             Instr)) ;
    mux21_ni ix117 (.Y (L1_4_L2_4_G5_MINI_ALU_OperationResult_1), .A0 (
             L1_4_L2_4_G5_MINI_ALU_BoothP_2), .A1 (WindowDin_4__4__1), .S0 (
             Instr)) ;
    mux21_ni ix125 (.Y (L1_4_L2_4_G5_MINI_ALU_OperationResult_2), .A0 (
             L1_4_L2_4_G5_MINI_ALU_BoothP_3), .A1 (WindowDin_4__4__2), .S0 (
             Instr)) ;
    mux21_ni ix133 (.Y (L1_4_L2_4_G5_MINI_ALU_OperationResult_3), .A0 (
             L1_4_L2_4_G5_MINI_ALU_BoothP_4), .A1 (WindowDin_4__4__3), .S0 (
             Instr)) ;
    mux21_ni ix141 (.Y (L1_4_L2_4_G5_MINI_ALU_OperationResult_4), .A0 (
             L1_4_L2_4_G5_MINI_ALU_BoothP_5), .A1 (WindowDin_4__4__4), .S0 (
             Instr)) ;
    mux21_ni ix149 (.Y (L1_4_L2_4_G5_MINI_ALU_OperationResult_5), .A0 (
             L1_4_L2_4_G5_MINI_ALU_BoothP_6), .A1 (WindowDin_4__4__5), .S0 (
             Instr)) ;
    mux21_ni ix157 (.Y (L1_4_L2_4_G5_MINI_ALU_OperationResult_6), .A0 (
             L1_4_L2_4_G5_MINI_ALU_BoothP_7), .A1 (WindowDin_4__4__6), .S0 (
             Instr)) ;
    mux21_ni ix165 (.Y (L1_4_L2_4_G5_MINI_ALU_OperationResult_7), .A0 (
             L1_4_L2_4_G5_MINI_ALU_BoothP_8), .A1 (WindowDin_4__4__7), .S0 (
             Instr)) ;
    nor02ii ix73 (.Y (L1_4_L2_4_G5_MINI_ALU_OperationResult_8), .A0 (Instr), .A1 (
            L1_4_L2_4_G5_MINI_ALU_BoothP_9)) ;
    nor02ii ix77 (.Y (L1_4_L2_4_G5_MINI_ALU_OperationResult_9), .A0 (Instr), .A1 (
            L1_4_L2_4_G5_MINI_ALU_BoothP_10)) ;
    nor02ii ix81 (.Y (L1_4_L2_4_G5_MINI_ALU_OperationResult_10), .A0 (Instr), .A1 (
            L1_4_L2_4_G5_MINI_ALU_BoothP_11)) ;
    nor02ii ix85 (.Y (L1_4_L2_4_G5_MINI_ALU_OperationResult_11), .A0 (Instr), .A1 (
            L1_4_L2_4_G5_MINI_ALU_BoothP_12)) ;
    nor02ii ix89 (.Y (L1_4_L2_4_G5_MINI_ALU_OperationResult_12), .A0 (Instr), .A1 (
            L1_4_L2_4_G5_MINI_ALU_BoothP_13)) ;
    nor02ii ix93 (.Y (L1_4_L2_4_G5_MINI_ALU_OperationResult_13), .A0 (Instr), .A1 (
            L1_4_L2_4_G5_MINI_ALU_BoothP_14)) ;
    nor02ii ix97 (.Y (L1_4_L2_4_G5_MINI_ALU_OperationResult_14), .A0 (Instr), .A1 (
            L1_4_L2_4_G5_MINI_ALU_BoothP_15)) ;
    nor02ii ix101 (.Y (L1_4_L2_4_G5_MINI_ALU_OperationResult_15), .A0 (Instr), .A1 (
            L1_4_L2_4_G5_MINI_ALU_BoothP_16)) ;
    mux21_ni ix1121 (.Y (L1_2_L2_1_G1_MINI_ALU_OperationResult_0), .A0 (
             L1_2_L2_1_G1_MINI_ALU_BoothP_1), .A1 (WindowDin_2__1__0), .S0 (
             Instr)) ;
    mux21_ni ix1129 (.Y (L1_2_L2_1_G1_MINI_ALU_OperationResult_1), .A0 (
             L1_2_L2_1_G1_MINI_ALU_BoothP_2), .A1 (WindowDin_2__1__1), .S0 (
             Instr)) ;
    mux21_ni ix1137 (.Y (L1_2_L2_1_G1_MINI_ALU_OperationResult_2), .A0 (
             L1_2_L2_1_G1_MINI_ALU_BoothP_3), .A1 (WindowDin_2__1__2), .S0 (
             Instr)) ;
    mux21_ni ix1145 (.Y (L1_2_L2_1_G1_MINI_ALU_OperationResult_3), .A0 (
             L1_2_L2_1_G1_MINI_ALU_BoothP_4), .A1 (WindowDin_2__1__3), .S0 (
             Instr)) ;
    mux21_ni ix1153 (.Y (L1_2_L2_1_G1_MINI_ALU_OperationResult_4), .A0 (
             L1_2_L2_1_G1_MINI_ALU_BoothP_5), .A1 (WindowDin_2__1__4), .S0 (
             Instr)) ;
    mux21_ni ix1161 (.Y (L1_2_L2_1_G1_MINI_ALU_OperationResult_5), .A0 (
             L1_2_L2_1_G1_MINI_ALU_BoothP_6), .A1 (WindowDin_2__1__5), .S0 (
             Instr)) ;
    mux21_ni ix1169 (.Y (L1_2_L2_1_G1_MINI_ALU_OperationResult_6), .A0 (
             L1_2_L2_1_G1_MINI_ALU_BoothP_7), .A1 (WindowDin_2__1__6), .S0 (
             Instr)) ;
    mux21_ni ix1177 (.Y (L1_2_L2_1_G1_MINI_ALU_OperationResult_7), .A0 (
             L1_2_L2_1_G1_MINI_ALU_BoothP_8), .A1 (WindowDin_2__1__7), .S0 (
             Instr)) ;
    nor02ii ix1085 (.Y (L1_2_L2_1_G1_MINI_ALU_OperationResult_8), .A0 (Instr), .A1 (
            L1_2_L2_1_G1_MINI_ALU_BoothP_9)) ;
    nor02ii ix1089 (.Y (L1_2_L2_1_G1_MINI_ALU_OperationResult_9), .A0 (Instr), .A1 (
            L1_2_L2_1_G1_MINI_ALU_BoothP_10)) ;
    nor02ii ix1093 (.Y (L1_2_L2_1_G1_MINI_ALU_OperationResult_10), .A0 (Instr), 
            .A1 (L1_2_L2_1_G1_MINI_ALU_BoothP_11)) ;
    nor02ii ix1097 (.Y (L1_2_L2_1_G1_MINI_ALU_OperationResult_11), .A0 (Instr), 
            .A1 (L1_2_L2_1_G1_MINI_ALU_BoothP_12)) ;
    nor02ii ix1101 (.Y (L1_2_L2_1_G1_MINI_ALU_OperationResult_12), .A0 (Instr), 
            .A1 (L1_2_L2_1_G1_MINI_ALU_BoothP_13)) ;
    nor02ii ix1105 (.Y (L1_2_L2_1_G1_MINI_ALU_OperationResult_13), .A0 (Instr), 
            .A1 (L1_2_L2_1_G1_MINI_ALU_BoothP_14)) ;
    nor02ii ix1109 (.Y (L1_2_L2_1_G1_MINI_ALU_OperationResult_14), .A0 (Instr), 
            .A1 (L1_2_L2_1_G1_MINI_ALU_BoothP_15)) ;
    nor02ii ix1113 (.Y (L1_2_L2_1_G1_MINI_ALU_OperationResult_15), .A0 (Instr), 
            .A1 (L1_2_L2_1_G1_MINI_ALU_BoothP_16)) ;
    mux21_ni ix1217 (.Y (L1_2_L2_0_G1_MINI_ALU_OperationResult_0), .A0 (
             L1_2_L2_0_G1_MINI_ALU_BoothP_1), .A1 (WindowDin_2__0__0), .S0 (
             Instr)) ;
    mux21_ni ix1225 (.Y (L1_2_L2_0_G1_MINI_ALU_OperationResult_1), .A0 (
             L1_2_L2_0_G1_MINI_ALU_BoothP_2), .A1 (WindowDin_2__0__1), .S0 (
             Instr)) ;
    mux21_ni ix1233 (.Y (L1_2_L2_0_G1_MINI_ALU_OperationResult_2), .A0 (
             L1_2_L2_0_G1_MINI_ALU_BoothP_3), .A1 (WindowDin_2__0__2), .S0 (
             Instr)) ;
    mux21_ni ix1241 (.Y (L1_2_L2_0_G1_MINI_ALU_OperationResult_3), .A0 (
             L1_2_L2_0_G1_MINI_ALU_BoothP_4), .A1 (WindowDin_2__0__3), .S0 (
             Instr)) ;
    mux21_ni ix1249 (.Y (L1_2_L2_0_G1_MINI_ALU_OperationResult_4), .A0 (
             L1_2_L2_0_G1_MINI_ALU_BoothP_5), .A1 (WindowDin_2__0__4), .S0 (
             Instr)) ;
    mux21_ni ix1257 (.Y (L1_2_L2_0_G1_MINI_ALU_OperationResult_5), .A0 (
             L1_2_L2_0_G1_MINI_ALU_BoothP_6), .A1 (WindowDin_2__0__5), .S0 (
             Instr)) ;
    mux21_ni ix1265 (.Y (L1_2_L2_0_G1_MINI_ALU_OperationResult_6), .A0 (
             L1_2_L2_0_G1_MINI_ALU_BoothP_7), .A1 (WindowDin_2__0__6), .S0 (
             Instr)) ;
    mux21_ni ix1273 (.Y (L1_2_L2_0_G1_MINI_ALU_OperationResult_7), .A0 (
             L1_2_L2_0_G1_MINI_ALU_BoothP_8), .A1 (WindowDin_2__0__7), .S0 (
             Instr)) ;
    nor02ii ix1181 (.Y (L1_2_L2_0_G1_MINI_ALU_OperationResult_8), .A0 (Instr), .A1 (
            L1_2_L2_0_G1_MINI_ALU_BoothP_9)) ;
    nor02ii ix1185 (.Y (L1_2_L2_0_G1_MINI_ALU_OperationResult_9), .A0 (Instr), .A1 (
            L1_2_L2_0_G1_MINI_ALU_BoothP_10)) ;
    nor02ii ix1189 (.Y (L1_2_L2_0_G1_MINI_ALU_OperationResult_10), .A0 (Instr), 
            .A1 (L1_2_L2_0_G1_MINI_ALU_BoothP_11)) ;
    nor02ii ix1193 (.Y (L1_2_L2_0_G1_MINI_ALU_OperationResult_11), .A0 (Instr), 
            .A1 (L1_2_L2_0_G1_MINI_ALU_BoothP_12)) ;
    nor02ii ix1197 (.Y (L1_2_L2_0_G1_MINI_ALU_OperationResult_12), .A0 (Instr), 
            .A1 (L1_2_L2_0_G1_MINI_ALU_BoothP_13)) ;
    nor02ii ix1201 (.Y (L1_2_L2_0_G1_MINI_ALU_OperationResult_13), .A0 (Instr), 
            .A1 (L1_2_L2_0_G1_MINI_ALU_BoothP_14)) ;
    nor02ii ix1205 (.Y (L1_2_L2_0_G1_MINI_ALU_OperationResult_14), .A0 (Instr), 
            .A1 (L1_2_L2_0_G1_MINI_ALU_BoothP_15)) ;
    nor02ii ix1209 (.Y (L1_2_L2_0_G1_MINI_ALU_OperationResult_15), .A0 (Instr), 
            .A1 (L1_2_L2_0_G1_MINI_ALU_BoothP_16)) ;
    mux21_ni ix1313 (.Y (L1_1_L2_4_G1_MINI_ALU_OperationResult_0), .A0 (
             L1_1_L2_4_G1_MINI_ALU_BoothP_1), .A1 (WindowDin_1__4__0), .S0 (
             Instr)) ;
    mux21_ni ix1321 (.Y (L1_1_L2_4_G1_MINI_ALU_OperationResult_1), .A0 (
             L1_1_L2_4_G1_MINI_ALU_BoothP_2), .A1 (WindowDin_1__4__1), .S0 (
             Instr)) ;
    mux21_ni ix1329 (.Y (L1_1_L2_4_G1_MINI_ALU_OperationResult_2), .A0 (
             L1_1_L2_4_G1_MINI_ALU_BoothP_3), .A1 (WindowDin_1__4__2), .S0 (
             Instr)) ;
    mux21_ni ix1337 (.Y (L1_1_L2_4_G1_MINI_ALU_OperationResult_3), .A0 (
             L1_1_L2_4_G1_MINI_ALU_BoothP_4), .A1 (WindowDin_1__4__3), .S0 (
             Instr)) ;
    mux21_ni ix1345 (.Y (L1_1_L2_4_G1_MINI_ALU_OperationResult_4), .A0 (
             L1_1_L2_4_G1_MINI_ALU_BoothP_5), .A1 (WindowDin_1__4__4), .S0 (
             Instr)) ;
    mux21_ni ix1353 (.Y (L1_1_L2_4_G1_MINI_ALU_OperationResult_5), .A0 (
             L1_1_L2_4_G1_MINI_ALU_BoothP_6), .A1 (WindowDin_1__4__5), .S0 (
             Instr)) ;
    mux21_ni ix1361 (.Y (L1_1_L2_4_G1_MINI_ALU_OperationResult_6), .A0 (
             L1_1_L2_4_G1_MINI_ALU_BoothP_7), .A1 (WindowDin_1__4__6), .S0 (
             Instr)) ;
    mux21_ni ix1369 (.Y (L1_1_L2_4_G1_MINI_ALU_OperationResult_7), .A0 (
             L1_1_L2_4_G1_MINI_ALU_BoothP_8), .A1 (WindowDin_1__4__7), .S0 (
             Instr)) ;
    nor02ii ix1277 (.Y (L1_1_L2_4_G1_MINI_ALU_OperationResult_8), .A0 (Instr), .A1 (
            L1_1_L2_4_G1_MINI_ALU_BoothP_9)) ;
    nor02ii ix1281 (.Y (L1_1_L2_4_G1_MINI_ALU_OperationResult_9), .A0 (Instr), .A1 (
            L1_1_L2_4_G1_MINI_ALU_BoothP_10)) ;
    nor02ii ix1285 (.Y (L1_1_L2_4_G1_MINI_ALU_OperationResult_10), .A0 (Instr), 
            .A1 (L1_1_L2_4_G1_MINI_ALU_BoothP_11)) ;
    nor02ii ix1289 (.Y (L1_1_L2_4_G1_MINI_ALU_OperationResult_11), .A0 (Instr), 
            .A1 (L1_1_L2_4_G1_MINI_ALU_BoothP_12)) ;
    nor02ii ix1293 (.Y (L1_1_L2_4_G1_MINI_ALU_OperationResult_12), .A0 (Instr), 
            .A1 (L1_1_L2_4_G1_MINI_ALU_BoothP_13)) ;
    nor02ii ix1297 (.Y (L1_1_L2_4_G1_MINI_ALU_OperationResult_13), .A0 (Instr), 
            .A1 (L1_1_L2_4_G1_MINI_ALU_BoothP_14)) ;
    nor02ii ix1301 (.Y (L1_1_L2_4_G1_MINI_ALU_OperationResult_14), .A0 (Instr), 
            .A1 (L1_1_L2_4_G1_MINI_ALU_BoothP_15)) ;
    nor02ii ix1305 (.Y (L1_1_L2_4_G1_MINI_ALU_OperationResult_15), .A0 (Instr), 
            .A1 (L1_1_L2_4_G1_MINI_ALU_BoothP_16)) ;
    mux21_ni ix1409 (.Y (L1_1_L2_3_G1_MINI_ALU_OperationResult_0), .A0 (
             L1_1_L2_3_G1_MINI_ALU_BoothP_1), .A1 (WindowDin_1__3__0), .S0 (
             Instr)) ;
    mux21_ni ix1417 (.Y (L1_1_L2_3_G1_MINI_ALU_OperationResult_1), .A0 (
             L1_1_L2_3_G1_MINI_ALU_BoothP_2), .A1 (WindowDin_1__3__1), .S0 (
             Instr)) ;
    mux21_ni ix1425 (.Y (L1_1_L2_3_G1_MINI_ALU_OperationResult_2), .A0 (
             L1_1_L2_3_G1_MINI_ALU_BoothP_3), .A1 (WindowDin_1__3__2), .S0 (
             Instr)) ;
    mux21_ni ix1433 (.Y (L1_1_L2_3_G1_MINI_ALU_OperationResult_3), .A0 (
             L1_1_L2_3_G1_MINI_ALU_BoothP_4), .A1 (WindowDin_1__3__3), .S0 (
             Instr)) ;
    mux21_ni ix1441 (.Y (L1_1_L2_3_G1_MINI_ALU_OperationResult_4), .A0 (
             L1_1_L2_3_G1_MINI_ALU_BoothP_5), .A1 (WindowDin_1__3__4), .S0 (
             Instr)) ;
    mux21_ni ix1449 (.Y (L1_1_L2_3_G1_MINI_ALU_OperationResult_5), .A0 (
             L1_1_L2_3_G1_MINI_ALU_BoothP_6), .A1 (WindowDin_1__3__5), .S0 (
             Instr)) ;
    mux21_ni ix1457 (.Y (L1_1_L2_3_G1_MINI_ALU_OperationResult_6), .A0 (
             L1_1_L2_3_G1_MINI_ALU_BoothP_7), .A1 (WindowDin_1__3__6), .S0 (
             Instr)) ;
    mux21_ni ix1465 (.Y (L1_1_L2_3_G1_MINI_ALU_OperationResult_7), .A0 (
             L1_1_L2_3_G1_MINI_ALU_BoothP_8), .A1 (WindowDin_1__3__7), .S0 (
             Instr)) ;
    nor02ii ix1373 (.Y (L1_1_L2_3_G1_MINI_ALU_OperationResult_8), .A0 (Instr), .A1 (
            L1_1_L2_3_G1_MINI_ALU_BoothP_9)) ;
    nor02ii ix1377 (.Y (L1_1_L2_3_G1_MINI_ALU_OperationResult_9), .A0 (Instr), .A1 (
            L1_1_L2_3_G1_MINI_ALU_BoothP_10)) ;
    nor02ii ix1381 (.Y (L1_1_L2_3_G1_MINI_ALU_OperationResult_10), .A0 (Instr), 
            .A1 (L1_1_L2_3_G1_MINI_ALU_BoothP_11)) ;
    nor02ii ix1385 (.Y (L1_1_L2_3_G1_MINI_ALU_OperationResult_11), .A0 (Instr), 
            .A1 (L1_1_L2_3_G1_MINI_ALU_BoothP_12)) ;
    nor02ii ix1389 (.Y (L1_1_L2_3_G1_MINI_ALU_OperationResult_12), .A0 (Instr), 
            .A1 (L1_1_L2_3_G1_MINI_ALU_BoothP_13)) ;
    nor02ii ix1393 (.Y (L1_1_L2_3_G1_MINI_ALU_OperationResult_13), .A0 (Instr), 
            .A1 (L1_1_L2_3_G1_MINI_ALU_BoothP_14)) ;
    nor02ii ix1397 (.Y (L1_1_L2_3_G1_MINI_ALU_OperationResult_14), .A0 (Instr), 
            .A1 (L1_1_L2_3_G1_MINI_ALU_BoothP_15)) ;
    nor02ii ix1401 (.Y (L1_1_L2_3_G1_MINI_ALU_OperationResult_15), .A0 (Instr), 
            .A1 (L1_1_L2_3_G1_MINI_ALU_BoothP_16)) ;
    mux21_ni ix1505 (.Y (L1_1_L2_2_G1_MINI_ALU_OperationResult_0), .A0 (
             L1_1_L2_2_G1_MINI_ALU_BoothP_1), .A1 (WindowDin_1__2__0), .S0 (
             Instr)) ;
    mux21_ni ix1513 (.Y (L1_1_L2_2_G1_MINI_ALU_OperationResult_1), .A0 (
             L1_1_L2_2_G1_MINI_ALU_BoothP_2), .A1 (WindowDin_1__2__1), .S0 (
             Instr)) ;
    mux21_ni ix1521 (.Y (L1_1_L2_2_G1_MINI_ALU_OperationResult_2), .A0 (
             L1_1_L2_2_G1_MINI_ALU_BoothP_3), .A1 (WindowDin_1__2__2), .S0 (
             Instr)) ;
    mux21_ni ix1529 (.Y (L1_1_L2_2_G1_MINI_ALU_OperationResult_3), .A0 (
             L1_1_L2_2_G1_MINI_ALU_BoothP_4), .A1 (WindowDin_1__2__3), .S0 (
             Instr)) ;
    mux21_ni ix1537 (.Y (L1_1_L2_2_G1_MINI_ALU_OperationResult_4), .A0 (
             L1_1_L2_2_G1_MINI_ALU_BoothP_5), .A1 (WindowDin_1__2__4), .S0 (
             Instr)) ;
    mux21_ni ix1545 (.Y (L1_1_L2_2_G1_MINI_ALU_OperationResult_5), .A0 (
             L1_1_L2_2_G1_MINI_ALU_BoothP_6), .A1 (WindowDin_1__2__5), .S0 (
             Instr)) ;
    mux21_ni ix1553 (.Y (L1_1_L2_2_G1_MINI_ALU_OperationResult_6), .A0 (
             L1_1_L2_2_G1_MINI_ALU_BoothP_7), .A1 (WindowDin_1__2__6), .S0 (
             Instr)) ;
    mux21_ni ix1561 (.Y (L1_1_L2_2_G1_MINI_ALU_OperationResult_7), .A0 (
             L1_1_L2_2_G1_MINI_ALU_BoothP_8), .A1 (WindowDin_1__2__7), .S0 (
             Instr)) ;
    nor02ii ix1469 (.Y (L1_1_L2_2_G1_MINI_ALU_OperationResult_8), .A0 (Instr), .A1 (
            L1_1_L2_2_G1_MINI_ALU_BoothP_9)) ;
    nor02ii ix1473 (.Y (L1_1_L2_2_G1_MINI_ALU_OperationResult_9), .A0 (Instr), .A1 (
            L1_1_L2_2_G1_MINI_ALU_BoothP_10)) ;
    nor02ii ix1477 (.Y (L1_1_L2_2_G1_MINI_ALU_OperationResult_10), .A0 (Instr), 
            .A1 (L1_1_L2_2_G1_MINI_ALU_BoothP_11)) ;
    nor02ii ix1481 (.Y (L1_1_L2_2_G1_MINI_ALU_OperationResult_11), .A0 (Instr), 
            .A1 (L1_1_L2_2_G1_MINI_ALU_BoothP_12)) ;
    nor02ii ix1485 (.Y (L1_1_L2_2_G1_MINI_ALU_OperationResult_12), .A0 (Instr), 
            .A1 (L1_1_L2_2_G1_MINI_ALU_BoothP_13)) ;
    nor02ii ix1489 (.Y (L1_1_L2_2_G1_MINI_ALU_OperationResult_13), .A0 (Instr), 
            .A1 (L1_1_L2_2_G1_MINI_ALU_BoothP_14)) ;
    nor02ii ix1493 (.Y (L1_1_L2_2_G1_MINI_ALU_OperationResult_14), .A0 (Instr), 
            .A1 (L1_1_L2_2_G1_MINI_ALU_BoothP_15)) ;
    nor02ii ix1497 (.Y (L1_1_L2_2_G1_MINI_ALU_OperationResult_15), .A0 (Instr), 
            .A1 (L1_1_L2_2_G1_MINI_ALU_BoothP_16)) ;
    mux21_ni ix1601 (.Y (L1_1_L2_1_G1_MINI_ALU_OperationResult_0), .A0 (
             L1_1_L2_1_G1_MINI_ALU_BoothP_1), .A1 (WindowDin_1__1__0), .S0 (
             Instr)) ;
    mux21_ni ix1609 (.Y (L1_1_L2_1_G1_MINI_ALU_OperationResult_1), .A0 (
             L1_1_L2_1_G1_MINI_ALU_BoothP_2), .A1 (WindowDin_1__1__1), .S0 (
             Instr)) ;
    mux21_ni ix1617 (.Y (L1_1_L2_1_G1_MINI_ALU_OperationResult_2), .A0 (
             L1_1_L2_1_G1_MINI_ALU_BoothP_3), .A1 (WindowDin_1__1__2), .S0 (
             Instr)) ;
    mux21_ni ix1625 (.Y (L1_1_L2_1_G1_MINI_ALU_OperationResult_3), .A0 (
             L1_1_L2_1_G1_MINI_ALU_BoothP_4), .A1 (WindowDin_1__1__3), .S0 (
             Instr)) ;
    mux21_ni ix1633 (.Y (L1_1_L2_1_G1_MINI_ALU_OperationResult_4), .A0 (
             L1_1_L2_1_G1_MINI_ALU_BoothP_5), .A1 (WindowDin_1__1__4), .S0 (
             Instr)) ;
    mux21_ni ix1641 (.Y (L1_1_L2_1_G1_MINI_ALU_OperationResult_5), .A0 (
             L1_1_L2_1_G1_MINI_ALU_BoothP_6), .A1 (WindowDin_1__1__5), .S0 (
             Instr)) ;
    mux21_ni ix1649 (.Y (L1_1_L2_1_G1_MINI_ALU_OperationResult_6), .A0 (
             L1_1_L2_1_G1_MINI_ALU_BoothP_7), .A1 (WindowDin_1__1__6), .S0 (
             Instr)) ;
    mux21_ni ix1657 (.Y (L1_1_L2_1_G1_MINI_ALU_OperationResult_7), .A0 (
             L1_1_L2_1_G1_MINI_ALU_BoothP_8), .A1 (WindowDin_1__1__7), .S0 (
             Instr)) ;
    nor02ii ix1565 (.Y (L1_1_L2_1_G1_MINI_ALU_OperationResult_8), .A0 (Instr), .A1 (
            L1_1_L2_1_G1_MINI_ALU_BoothP_9)) ;
    nor02ii ix1569 (.Y (L1_1_L2_1_G1_MINI_ALU_OperationResult_9), .A0 (Instr), .A1 (
            L1_1_L2_1_G1_MINI_ALU_BoothP_10)) ;
    nor02ii ix1573 (.Y (L1_1_L2_1_G1_MINI_ALU_OperationResult_10), .A0 (Instr), 
            .A1 (L1_1_L2_1_G1_MINI_ALU_BoothP_11)) ;
    nor02ii ix1577 (.Y (L1_1_L2_1_G1_MINI_ALU_OperationResult_11), .A0 (Instr), 
            .A1 (L1_1_L2_1_G1_MINI_ALU_BoothP_12)) ;
    nor02ii ix1581 (.Y (L1_1_L2_1_G1_MINI_ALU_OperationResult_12), .A0 (Instr), 
            .A1 (L1_1_L2_1_G1_MINI_ALU_BoothP_13)) ;
    nor02ii ix1585 (.Y (L1_1_L2_1_G1_MINI_ALU_OperationResult_13), .A0 (Instr), 
            .A1 (L1_1_L2_1_G1_MINI_ALU_BoothP_14)) ;
    nor02ii ix1589 (.Y (L1_1_L2_1_G1_MINI_ALU_OperationResult_14), .A0 (Instr), 
            .A1 (L1_1_L2_1_G1_MINI_ALU_BoothP_15)) ;
    nor02ii ix1593 (.Y (L1_1_L2_1_G1_MINI_ALU_OperationResult_15), .A0 (Instr), 
            .A1 (L1_1_L2_1_G1_MINI_ALU_BoothP_16)) ;
    mux21_ni ix1697 (.Y (L1_1_L2_0_G1_MINI_ALU_OperationResult_0), .A0 (
             L1_1_L2_0_G1_MINI_ALU_BoothP_1), .A1 (WindowDin_1__0__0), .S0 (
             Instr)) ;
    mux21_ni ix1705 (.Y (L1_1_L2_0_G1_MINI_ALU_OperationResult_1), .A0 (
             L1_1_L2_0_G1_MINI_ALU_BoothP_2), .A1 (WindowDin_1__0__1), .S0 (
             Instr)) ;
    mux21_ni ix1713 (.Y (L1_1_L2_0_G1_MINI_ALU_OperationResult_2), .A0 (
             L1_1_L2_0_G1_MINI_ALU_BoothP_3), .A1 (WindowDin_1__0__2), .S0 (
             Instr)) ;
    mux21_ni ix1721 (.Y (L1_1_L2_0_G1_MINI_ALU_OperationResult_3), .A0 (
             L1_1_L2_0_G1_MINI_ALU_BoothP_4), .A1 (WindowDin_1__0__3), .S0 (
             Instr)) ;
    mux21_ni ix1729 (.Y (L1_1_L2_0_G1_MINI_ALU_OperationResult_4), .A0 (
             L1_1_L2_0_G1_MINI_ALU_BoothP_5), .A1 (WindowDin_1__0__4), .S0 (
             Instr)) ;
    mux21_ni ix1737 (.Y (L1_1_L2_0_G1_MINI_ALU_OperationResult_5), .A0 (
             L1_1_L2_0_G1_MINI_ALU_BoothP_6), .A1 (WindowDin_1__0__5), .S0 (
             Instr)) ;
    mux21_ni ix1745 (.Y (L1_1_L2_0_G1_MINI_ALU_OperationResult_6), .A0 (
             L1_1_L2_0_G1_MINI_ALU_BoothP_7), .A1 (WindowDin_1__0__6), .S0 (
             Instr)) ;
    mux21_ni ix1753 (.Y (L1_1_L2_0_G1_MINI_ALU_OperationResult_7), .A0 (
             L1_1_L2_0_G1_MINI_ALU_BoothP_8), .A1 (WindowDin_1__0__7), .S0 (
             Instr)) ;
    nor02ii ix1661 (.Y (L1_1_L2_0_G1_MINI_ALU_OperationResult_8), .A0 (Instr), .A1 (
            L1_1_L2_0_G1_MINI_ALU_BoothP_9)) ;
    nor02ii ix1665 (.Y (L1_1_L2_0_G1_MINI_ALU_OperationResult_9), .A0 (Instr), .A1 (
            L1_1_L2_0_G1_MINI_ALU_BoothP_10)) ;
    nor02ii ix1669 (.Y (L1_1_L2_0_G1_MINI_ALU_OperationResult_10), .A0 (Instr), 
            .A1 (L1_1_L2_0_G1_MINI_ALU_BoothP_11)) ;
    nor02ii ix1673 (.Y (L1_1_L2_0_G1_MINI_ALU_OperationResult_11), .A0 (Instr), 
            .A1 (L1_1_L2_0_G1_MINI_ALU_BoothP_12)) ;
    nor02ii ix1677 (.Y (L1_1_L2_0_G1_MINI_ALU_OperationResult_12), .A0 (Instr), 
            .A1 (L1_1_L2_0_G1_MINI_ALU_BoothP_13)) ;
    nor02ii ix1681 (.Y (L1_1_L2_0_G1_MINI_ALU_OperationResult_13), .A0 (Instr), 
            .A1 (L1_1_L2_0_G1_MINI_ALU_BoothP_14)) ;
    nor02ii ix1685 (.Y (L1_1_L2_0_G1_MINI_ALU_OperationResult_14), .A0 (Instr), 
            .A1 (L1_1_L2_0_G1_MINI_ALU_BoothP_15)) ;
    nor02ii ix1689 (.Y (L1_1_L2_0_G1_MINI_ALU_OperationResult_15), .A0 (Instr), 
            .A1 (L1_1_L2_0_G1_MINI_ALU_BoothP_16)) ;
    mux21_ni ix1793 (.Y (L1_0_L2_4_G1_MINI_ALU_OperationResult_0), .A0 (
             L1_0_L2_4_G1_MINI_ALU_BoothP_1), .A1 (WindowDin_0__4__0), .S0 (
             Instr)) ;
    mux21_ni ix1801 (.Y (L1_0_L2_4_G1_MINI_ALU_OperationResult_1), .A0 (
             L1_0_L2_4_G1_MINI_ALU_BoothP_2), .A1 (WindowDin_0__4__1), .S0 (
             Instr)) ;
    mux21_ni ix1809 (.Y (L1_0_L2_4_G1_MINI_ALU_OperationResult_2), .A0 (
             L1_0_L2_4_G1_MINI_ALU_BoothP_3), .A1 (WindowDin_0__4__2), .S0 (
             Instr)) ;
    mux21_ni ix1817 (.Y (L1_0_L2_4_G1_MINI_ALU_OperationResult_3), .A0 (
             L1_0_L2_4_G1_MINI_ALU_BoothP_4), .A1 (WindowDin_0__4__3), .S0 (
             Instr)) ;
    mux21_ni ix1825 (.Y (L1_0_L2_4_G1_MINI_ALU_OperationResult_4), .A0 (
             L1_0_L2_4_G1_MINI_ALU_BoothP_5), .A1 (WindowDin_0__4__4), .S0 (
             Instr)) ;
    mux21_ni ix1833 (.Y (L1_0_L2_4_G1_MINI_ALU_OperationResult_5), .A0 (
             L1_0_L2_4_G1_MINI_ALU_BoothP_6), .A1 (WindowDin_0__4__5), .S0 (
             Instr)) ;
    mux21_ni ix1841 (.Y (L1_0_L2_4_G1_MINI_ALU_OperationResult_6), .A0 (
             L1_0_L2_4_G1_MINI_ALU_BoothP_7), .A1 (WindowDin_0__4__6), .S0 (
             Instr)) ;
    mux21_ni ix1849 (.Y (L1_0_L2_4_G1_MINI_ALU_OperationResult_7), .A0 (
             L1_0_L2_4_G1_MINI_ALU_BoothP_8), .A1 (WindowDin_0__4__7), .S0 (
             Instr)) ;
    nor02ii ix1757 (.Y (L1_0_L2_4_G1_MINI_ALU_OperationResult_8), .A0 (Instr), .A1 (
            L1_0_L2_4_G1_MINI_ALU_BoothP_9)) ;
    nor02ii ix1761 (.Y (L1_0_L2_4_G1_MINI_ALU_OperationResult_9), .A0 (Instr), .A1 (
            L1_0_L2_4_G1_MINI_ALU_BoothP_10)) ;
    nor02ii ix1765 (.Y (L1_0_L2_4_G1_MINI_ALU_OperationResult_10), .A0 (Instr), 
            .A1 (L1_0_L2_4_G1_MINI_ALU_BoothP_11)) ;
    nor02ii ix1769 (.Y (L1_0_L2_4_G1_MINI_ALU_OperationResult_11), .A0 (Instr), 
            .A1 (L1_0_L2_4_G1_MINI_ALU_BoothP_12)) ;
    nor02ii ix1773 (.Y (L1_0_L2_4_G1_MINI_ALU_OperationResult_12), .A0 (Instr), 
            .A1 (L1_0_L2_4_G1_MINI_ALU_BoothP_13)) ;
    nor02ii ix1777 (.Y (L1_0_L2_4_G1_MINI_ALU_OperationResult_13), .A0 (Instr), 
            .A1 (L1_0_L2_4_G1_MINI_ALU_BoothP_14)) ;
    nor02ii ix1781 (.Y (L1_0_L2_4_G1_MINI_ALU_OperationResult_14), .A0 (Instr), 
            .A1 (L1_0_L2_4_G1_MINI_ALU_BoothP_15)) ;
    nor02ii ix1785 (.Y (L1_0_L2_4_G1_MINI_ALU_OperationResult_15), .A0 (Instr), 
            .A1 (L1_0_L2_4_G1_MINI_ALU_BoothP_16)) ;
    mux21_ni ix1889 (.Y (L1_0_L2_3_G1_MINI_ALU_OperationResult_0), .A0 (
             L1_0_L2_3_G1_MINI_ALU_BoothP_1), .A1 (WindowDin_0__3__0), .S0 (
             Instr)) ;
    mux21_ni ix1897 (.Y (L1_0_L2_3_G1_MINI_ALU_OperationResult_1), .A0 (
             L1_0_L2_3_G1_MINI_ALU_BoothP_2), .A1 (WindowDin_0__3__1), .S0 (
             Instr)) ;
    mux21_ni ix1905 (.Y (L1_0_L2_3_G1_MINI_ALU_OperationResult_2), .A0 (
             L1_0_L2_3_G1_MINI_ALU_BoothP_3), .A1 (WindowDin_0__3__2), .S0 (
             Instr)) ;
    mux21_ni ix1913 (.Y (L1_0_L2_3_G1_MINI_ALU_OperationResult_3), .A0 (
             L1_0_L2_3_G1_MINI_ALU_BoothP_4), .A1 (WindowDin_0__3__3), .S0 (
             Instr)) ;
    mux21_ni ix1921 (.Y (L1_0_L2_3_G1_MINI_ALU_OperationResult_4), .A0 (
             L1_0_L2_3_G1_MINI_ALU_BoothP_5), .A1 (WindowDin_0__3__4), .S0 (
             Instr)) ;
    mux21_ni ix1929 (.Y (L1_0_L2_3_G1_MINI_ALU_OperationResult_5), .A0 (
             L1_0_L2_3_G1_MINI_ALU_BoothP_6), .A1 (WindowDin_0__3__5), .S0 (
             Instr)) ;
    mux21_ni ix1937 (.Y (L1_0_L2_3_G1_MINI_ALU_OperationResult_6), .A0 (
             L1_0_L2_3_G1_MINI_ALU_BoothP_7), .A1 (WindowDin_0__3__6), .S0 (
             Instr)) ;
    mux21_ni ix1945 (.Y (L1_0_L2_3_G1_MINI_ALU_OperationResult_7), .A0 (
             L1_0_L2_3_G1_MINI_ALU_BoothP_8), .A1 (WindowDin_0__3__7), .S0 (
             Instr)) ;
    nor02ii ix1853 (.Y (L1_0_L2_3_G1_MINI_ALU_OperationResult_8), .A0 (Instr), .A1 (
            L1_0_L2_3_G1_MINI_ALU_BoothP_9)) ;
    nor02ii ix1857 (.Y (L1_0_L2_3_G1_MINI_ALU_OperationResult_9), .A0 (Instr), .A1 (
            L1_0_L2_3_G1_MINI_ALU_BoothP_10)) ;
    nor02ii ix1861 (.Y (L1_0_L2_3_G1_MINI_ALU_OperationResult_10), .A0 (Instr), 
            .A1 (L1_0_L2_3_G1_MINI_ALU_BoothP_11)) ;
    nor02ii ix1865 (.Y (L1_0_L2_3_G1_MINI_ALU_OperationResult_11), .A0 (Instr), 
            .A1 (L1_0_L2_3_G1_MINI_ALU_BoothP_12)) ;
    nor02ii ix1869 (.Y (L1_0_L2_3_G1_MINI_ALU_OperationResult_12), .A0 (Instr), 
            .A1 (L1_0_L2_3_G1_MINI_ALU_BoothP_13)) ;
    nor02ii ix1873 (.Y (L1_0_L2_3_G1_MINI_ALU_OperationResult_13), .A0 (Instr), 
            .A1 (L1_0_L2_3_G1_MINI_ALU_BoothP_14)) ;
    nor02ii ix1877 (.Y (L1_0_L2_3_G1_MINI_ALU_OperationResult_14), .A0 (Instr), 
            .A1 (L1_0_L2_3_G1_MINI_ALU_BoothP_15)) ;
    nor02ii ix1881 (.Y (L1_0_L2_3_G1_MINI_ALU_OperationResult_15), .A0 (Instr), 
            .A1 (L1_0_L2_3_G1_MINI_ALU_BoothP_16)) ;
    mux21_ni ix1985 (.Y (L1_0_L2_2_G1_MINI_ALU_OperationResult_0), .A0 (
             L1_0_L2_2_G1_MINI_ALU_BoothP_1), .A1 (WindowDin_0__2__0), .S0 (
             Instr)) ;
    mux21_ni ix1993 (.Y (L1_0_L2_2_G1_MINI_ALU_OperationResult_1), .A0 (
             L1_0_L2_2_G1_MINI_ALU_BoothP_2), .A1 (WindowDin_0__2__1), .S0 (
             Instr)) ;
    mux21_ni ix2001 (.Y (L1_0_L2_2_G1_MINI_ALU_OperationResult_2), .A0 (
             L1_0_L2_2_G1_MINI_ALU_BoothP_3), .A1 (WindowDin_0__2__2), .S0 (
             Instr)) ;
    mux21_ni ix2009 (.Y (L1_0_L2_2_G1_MINI_ALU_OperationResult_3), .A0 (
             L1_0_L2_2_G1_MINI_ALU_BoothP_4), .A1 (WindowDin_0__2__3), .S0 (
             Instr)) ;
    mux21_ni ix2017 (.Y (L1_0_L2_2_G1_MINI_ALU_OperationResult_4), .A0 (
             L1_0_L2_2_G1_MINI_ALU_BoothP_5), .A1 (WindowDin_0__2__4), .S0 (
             Instr)) ;
    mux21_ni ix2025 (.Y (L1_0_L2_2_G1_MINI_ALU_OperationResult_5), .A0 (
             L1_0_L2_2_G1_MINI_ALU_BoothP_6), .A1 (WindowDin_0__2__5), .S0 (
             Instr)) ;
    mux21_ni ix2033 (.Y (L1_0_L2_2_G1_MINI_ALU_OperationResult_6), .A0 (
             L1_0_L2_2_G1_MINI_ALU_BoothP_7), .A1 (WindowDin_0__2__6), .S0 (
             Instr)) ;
    mux21_ni ix2041 (.Y (L1_0_L2_2_G1_MINI_ALU_OperationResult_7), .A0 (
             L1_0_L2_2_G1_MINI_ALU_BoothP_8), .A1 (WindowDin_0__2__7), .S0 (
             Instr)) ;
    nor02ii ix1949 (.Y (L1_0_L2_2_G1_MINI_ALU_OperationResult_8), .A0 (Instr), .A1 (
            L1_0_L2_2_G1_MINI_ALU_BoothP_9)) ;
    nor02ii ix1953 (.Y (L1_0_L2_2_G1_MINI_ALU_OperationResult_9), .A0 (Instr), .A1 (
            L1_0_L2_2_G1_MINI_ALU_BoothP_10)) ;
    nor02ii ix1957 (.Y (L1_0_L2_2_G1_MINI_ALU_OperationResult_10), .A0 (Instr), 
            .A1 (L1_0_L2_2_G1_MINI_ALU_BoothP_11)) ;
    nor02ii ix1961 (.Y (L1_0_L2_2_G1_MINI_ALU_OperationResult_11), .A0 (Instr), 
            .A1 (L1_0_L2_2_G1_MINI_ALU_BoothP_12)) ;
    nor02ii ix1965 (.Y (L1_0_L2_2_G1_MINI_ALU_OperationResult_12), .A0 (Instr), 
            .A1 (L1_0_L2_2_G1_MINI_ALU_BoothP_13)) ;
    nor02ii ix1969 (.Y (L1_0_L2_2_G1_MINI_ALU_OperationResult_13), .A0 (Instr), 
            .A1 (L1_0_L2_2_G1_MINI_ALU_BoothP_14)) ;
    nor02ii ix1973 (.Y (L1_0_L2_2_G1_MINI_ALU_OperationResult_14), .A0 (Instr), 
            .A1 (L1_0_L2_2_G1_MINI_ALU_BoothP_15)) ;
    nor02ii ix1977 (.Y (L1_0_L2_2_G1_MINI_ALU_OperationResult_15), .A0 (Instr), 
            .A1 (L1_0_L2_2_G1_MINI_ALU_BoothP_16)) ;
    mux21_ni ix2081 (.Y (L1_0_L2_1_G1_MINI_ALU_OperationResult_0), .A0 (
             L1_0_L2_1_G1_MINI_ALU_BoothP_1), .A1 (WindowDin_0__1__0), .S0 (
             Instr)) ;
    mux21_ni ix2089 (.Y (L1_0_L2_1_G1_MINI_ALU_OperationResult_1), .A0 (
             L1_0_L2_1_G1_MINI_ALU_BoothP_2), .A1 (WindowDin_0__1__1), .S0 (
             Instr)) ;
    mux21_ni ix2097 (.Y (L1_0_L2_1_G1_MINI_ALU_OperationResult_2), .A0 (
             L1_0_L2_1_G1_MINI_ALU_BoothP_3), .A1 (WindowDin_0__1__2), .S0 (
             Instr)) ;
    mux21_ni ix2105 (.Y (L1_0_L2_1_G1_MINI_ALU_OperationResult_3), .A0 (
             L1_0_L2_1_G1_MINI_ALU_BoothP_4), .A1 (WindowDin_0__1__3), .S0 (
             Instr)) ;
    mux21_ni ix2113 (.Y (L1_0_L2_1_G1_MINI_ALU_OperationResult_4), .A0 (
             L1_0_L2_1_G1_MINI_ALU_BoothP_5), .A1 (WindowDin_0__1__4), .S0 (
             Instr)) ;
    mux21_ni ix2121 (.Y (L1_0_L2_1_G1_MINI_ALU_OperationResult_5), .A0 (
             L1_0_L2_1_G1_MINI_ALU_BoothP_6), .A1 (WindowDin_0__1__5), .S0 (
             Instr)) ;
    mux21_ni ix2129 (.Y (L1_0_L2_1_G1_MINI_ALU_OperationResult_6), .A0 (
             L1_0_L2_1_G1_MINI_ALU_BoothP_7), .A1 (WindowDin_0__1__6), .S0 (
             Instr)) ;
    mux21_ni ix2137 (.Y (L1_0_L2_1_G1_MINI_ALU_OperationResult_7), .A0 (
             L1_0_L2_1_G1_MINI_ALU_BoothP_8), .A1 (WindowDin_0__1__7), .S0 (
             Instr)) ;
    nor02ii ix2045 (.Y (L1_0_L2_1_G1_MINI_ALU_OperationResult_8), .A0 (Instr), .A1 (
            L1_0_L2_1_G1_MINI_ALU_BoothP_9)) ;
    nor02ii ix2049 (.Y (L1_0_L2_1_G1_MINI_ALU_OperationResult_9), .A0 (Instr), .A1 (
            L1_0_L2_1_G1_MINI_ALU_BoothP_10)) ;
    nor02ii ix2053 (.Y (L1_0_L2_1_G1_MINI_ALU_OperationResult_10), .A0 (Instr), 
            .A1 (L1_0_L2_1_G1_MINI_ALU_BoothP_11)) ;
    nor02ii ix2057 (.Y (L1_0_L2_1_G1_MINI_ALU_OperationResult_11), .A0 (Instr), 
            .A1 (L1_0_L2_1_G1_MINI_ALU_BoothP_12)) ;
    nor02ii ix2061 (.Y (L1_0_L2_1_G1_MINI_ALU_OperationResult_12), .A0 (Instr), 
            .A1 (L1_0_L2_1_G1_MINI_ALU_BoothP_13)) ;
    nor02ii ix2065 (.Y (L1_0_L2_1_G1_MINI_ALU_OperationResult_13), .A0 (Instr), 
            .A1 (L1_0_L2_1_G1_MINI_ALU_BoothP_14)) ;
    nor02ii ix2069 (.Y (L1_0_L2_1_G1_MINI_ALU_OperationResult_14), .A0 (Instr), 
            .A1 (L1_0_L2_1_G1_MINI_ALU_BoothP_15)) ;
    nor02ii ix2073 (.Y (L1_0_L2_1_G1_MINI_ALU_OperationResult_15), .A0 (Instr), 
            .A1 (L1_0_L2_1_G1_MINI_ALU_BoothP_16)) ;
    mux21_ni ix2177 (.Y (L1_0_L2_0_G1_MINI_ALU_OperationResult_0), .A0 (
             L1_0_L2_0_G1_MINI_ALU_BoothP_1), .A1 (WindowDin_0__0__0), .S0 (
             Instr)) ;
    mux21_ni ix2185 (.Y (L1_0_L2_0_G1_MINI_ALU_OperationResult_1), .A0 (
             L1_0_L2_0_G1_MINI_ALU_BoothP_2), .A1 (WindowDin_0__0__1), .S0 (
             Instr)) ;
    mux21_ni ix2193 (.Y (L1_0_L2_0_G1_MINI_ALU_OperationResult_2), .A0 (
             L1_0_L2_0_G1_MINI_ALU_BoothP_3), .A1 (WindowDin_0__0__2), .S0 (
             Instr)) ;
    mux21_ni ix2201 (.Y (L1_0_L2_0_G1_MINI_ALU_OperationResult_3), .A0 (
             L1_0_L2_0_G1_MINI_ALU_BoothP_4), .A1 (WindowDin_0__0__3), .S0 (
             Instr)) ;
    mux21_ni ix2209 (.Y (L1_0_L2_0_G1_MINI_ALU_OperationResult_4), .A0 (
             L1_0_L2_0_G1_MINI_ALU_BoothP_5), .A1 (WindowDin_0__0__4), .S0 (
             Instr)) ;
    mux21_ni ix2217 (.Y (L1_0_L2_0_G1_MINI_ALU_OperationResult_5), .A0 (
             L1_0_L2_0_G1_MINI_ALU_BoothP_6), .A1 (WindowDin_0__0__5), .S0 (
             Instr)) ;
    mux21_ni ix2225 (.Y (L1_0_L2_0_G1_MINI_ALU_OperationResult_6), .A0 (
             L1_0_L2_0_G1_MINI_ALU_BoothP_7), .A1 (WindowDin_0__0__6), .S0 (
             Instr)) ;
    mux21_ni ix2233 (.Y (L1_0_L2_0_G1_MINI_ALU_OperationResult_7), .A0 (
             L1_0_L2_0_G1_MINI_ALU_BoothP_8), .A1 (WindowDin_0__0__7), .S0 (
             Instr)) ;
    nor02ii ix2141 (.Y (L1_0_L2_0_G1_MINI_ALU_OperationResult_8), .A0 (Instr), .A1 (
            L1_0_L2_0_G1_MINI_ALU_BoothP_9)) ;
    nor02ii ix2145 (.Y (L1_0_L2_0_G1_MINI_ALU_OperationResult_9), .A0 (Instr), .A1 (
            L1_0_L2_0_G1_MINI_ALU_BoothP_10)) ;
    nor02ii ix2149 (.Y (L1_0_L2_0_G1_MINI_ALU_OperationResult_10), .A0 (Instr), 
            .A1 (L1_0_L2_0_G1_MINI_ALU_BoothP_11)) ;
    nor02ii ix2153 (.Y (L1_0_L2_0_G1_MINI_ALU_OperationResult_11), .A0 (Instr), 
            .A1 (L1_0_L2_0_G1_MINI_ALU_BoothP_12)) ;
    nor02ii ix2157 (.Y (L1_0_L2_0_G1_MINI_ALU_OperationResult_12), .A0 (Instr), 
            .A1 (L1_0_L2_0_G1_MINI_ALU_BoothP_13)) ;
    nor02ii ix2161 (.Y (L1_0_L2_0_G1_MINI_ALU_OperationResult_13), .A0 (Instr), 
            .A1 (L1_0_L2_0_G1_MINI_ALU_BoothP_14)) ;
    nor02ii ix2165 (.Y (L1_0_L2_0_G1_MINI_ALU_OperationResult_14), .A0 (Instr), 
            .A1 (L1_0_L2_0_G1_MINI_ALU_BoothP_15)) ;
    nor02ii ix2169 (.Y (L1_0_L2_0_G1_MINI_ALU_OperationResult_15), .A0 (Instr), 
            .A1 (L1_0_L2_0_G1_MINI_ALU_BoothP_16)) ;
    mux21_ni ix973 (.Y (L1FirstOperands_11__0), .A0 (
             L1_2_L2_2_G1_MINI_ALU_BoothP_1), .A1 (WindowDin_2__2__0), .S0 (
             Instr)) ;
    mux21_ni ix981 (.Y (L1FirstOperands_11__1), .A0 (
             L1_2_L2_2_G1_MINI_ALU_BoothP_2), .A1 (WindowDin_2__2__1), .S0 (
             Instr)) ;
    mux21_ni ix989 (.Y (L1FirstOperands_11__2), .A0 (
             L1_2_L2_2_G1_MINI_ALU_BoothP_3), .A1 (WindowDin_2__2__2), .S0 (
             Instr)) ;
    mux21_ni ix997 (.Y (L1FirstOperands_11__3), .A0 (
             L1_2_L2_2_G1_MINI_ALU_BoothP_4), .A1 (WindowDin_2__2__3), .S0 (
             Instr)) ;
    mux21_ni ix1005 (.Y (L1FirstOperands_11__4), .A0 (
             L1_2_L2_2_G1_MINI_ALU_BoothP_5), .A1 (WindowDin_2__2__4), .S0 (
             Instr)) ;
    mux21_ni ix1013 (.Y (L1FirstOperands_11__5), .A0 (
             L1_2_L2_2_G1_MINI_ALU_BoothP_6), .A1 (WindowDin_2__2__5), .S0 (
             Instr)) ;
    mux21_ni ix1021 (.Y (L1FirstOperands_11__6), .A0 (
             L1_2_L2_2_G1_MINI_ALU_BoothP_7), .A1 (WindowDin_2__2__6), .S0 (
             Instr)) ;
    mux21_ni ix1029 (.Y (L1FirstOperands_11__7), .A0 (
             L1_2_L2_2_G1_MINI_ALU_BoothP_8), .A1 (WindowDin_2__2__7), .S0 (
             Instr)) ;
    nor02ii ix937 (.Y (L1FirstOperands_11__8), .A0 (Instr), .A1 (
            L1_2_L2_2_G1_MINI_ALU_BoothP_9)) ;
    nor02ii ix941 (.Y (L1FirstOperands_11__9), .A0 (Instr), .A1 (
            L1_2_L2_2_G1_MINI_ALU_BoothP_10)) ;
    nor02ii ix945 (.Y (L1FirstOperands_11__10), .A0 (Instr), .A1 (
            L1_2_L2_2_G1_MINI_ALU_BoothP_11)) ;
    nor02ii ix949 (.Y (L1FirstOperands_11__11), .A0 (Instr), .A1 (
            L1_2_L2_2_G1_MINI_ALU_BoothP_12)) ;
    nor02ii ix953 (.Y (L1FirstOperands_11__12), .A0 (Instr), .A1 (
            L1_2_L2_2_G1_MINI_ALU_BoothP_13)) ;
    nor02ii ix957 (.Y (L1FirstOperands_11__13), .A0 (Instr), .A1 (
            L1_2_L2_2_G1_MINI_ALU_BoothP_14)) ;
    nor02ii ix961 (.Y (L1FirstOperands_11__14), .A0 (Instr), .A1 (
            L1_2_L2_2_G1_MINI_ALU_BoothP_15)) ;
    nor02ii ix965 (.Y (L1FirstOperands_11__15), .A0 (Instr), .A1 (
            L1_2_L2_2_G1_MINI_ALU_BoothP_16)) ;
    mux21_ni ix397 (.Y (L1FirstOperands_10__0), .A0 (
             L1_3_L2_3_G2_MINI_ALU_BoothP_1), .A1 (WindowDin_3__3__0), .S0 (
             Instr)) ;
    mux21_ni ix405 (.Y (L1FirstOperands_10__1), .A0 (
             L1_3_L2_3_G2_MINI_ALU_BoothP_2), .A1 (WindowDin_3__3__1), .S0 (
             Instr)) ;
    mux21_ni ix413 (.Y (L1FirstOperands_10__2), .A0 (
             L1_3_L2_3_G2_MINI_ALU_BoothP_3), .A1 (WindowDin_3__3__2), .S0 (
             Instr)) ;
    mux21_ni ix421 (.Y (L1FirstOperands_10__3), .A0 (
             L1_3_L2_3_G2_MINI_ALU_BoothP_4), .A1 (WindowDin_3__3__3), .S0 (
             Instr)) ;
    mux21_ni ix429 (.Y (L1FirstOperands_10__4), .A0 (
             L1_3_L2_3_G2_MINI_ALU_BoothP_5), .A1 (WindowDin_3__3__4), .S0 (
             Instr)) ;
    mux21_ni ix437 (.Y (L1FirstOperands_10__5), .A0 (
             L1_3_L2_3_G2_MINI_ALU_BoothP_6), .A1 (WindowDin_3__3__5), .S0 (
             Instr)) ;
    mux21_ni ix445 (.Y (L1FirstOperands_10__6), .A0 (
             L1_3_L2_3_G2_MINI_ALU_BoothP_7), .A1 (WindowDin_3__3__6), .S0 (
             Instr)) ;
    mux21_ni ix453 (.Y (L1FirstOperands_10__7), .A0 (
             L1_3_L2_3_G2_MINI_ALU_BoothP_8), .A1 (WindowDin_3__3__7), .S0 (
             Instr)) ;
    nor02ii ix361 (.Y (L1FirstOperands_10__8), .A0 (Instr), .A1 (
            L1_3_L2_3_G2_MINI_ALU_BoothP_9)) ;
    nor02ii ix365 (.Y (L1FirstOperands_10__9), .A0 (Instr), .A1 (
            L1_3_L2_3_G2_MINI_ALU_BoothP_10)) ;
    nor02ii ix369 (.Y (L1FirstOperands_10__10), .A0 (Instr), .A1 (
            L1_3_L2_3_G2_MINI_ALU_BoothP_11)) ;
    nor02ii ix373 (.Y (L1FirstOperands_10__11), .A0 (Instr), .A1 (
            L1_3_L2_3_G2_MINI_ALU_BoothP_12)) ;
    nor02ii ix377 (.Y (L1FirstOperands_10__12), .A0 (Instr), .A1 (
            L1_3_L2_3_G2_MINI_ALU_BoothP_13)) ;
    nor02ii ix381 (.Y (L1FirstOperands_10__13), .A0 (Instr), .A1 (
            L1_3_L2_3_G2_MINI_ALU_BoothP_14)) ;
    nor02ii ix385 (.Y (L1FirstOperands_10__14), .A0 (Instr), .A1 (
            L1_3_L2_3_G2_MINI_ALU_BoothP_15)) ;
    nor02ii ix389 (.Y (L1FirstOperands_10__15), .A0 (Instr), .A1 (
            L1_3_L2_3_G2_MINI_ALU_BoothP_16)) ;
    mux21_ni ix493 (.Y (L1FirstOperands_8__0), .A0 (
             L1_3_L2_2_G2_MINI_ALU_BoothP_1), .A1 (WindowDin_3__2__0), .S0 (
             Instr)) ;
    mux21_ni ix501 (.Y (L1FirstOperands_8__1), .A0 (
             L1_3_L2_2_G2_MINI_ALU_BoothP_2), .A1 (WindowDin_3__2__1), .S0 (
             Instr)) ;
    mux21_ni ix509 (.Y (L1FirstOperands_8__2), .A0 (
             L1_3_L2_2_G2_MINI_ALU_BoothP_3), .A1 (WindowDin_3__2__2), .S0 (
             Instr)) ;
    mux21_ni ix517 (.Y (L1FirstOperands_8__3), .A0 (
             L1_3_L2_2_G2_MINI_ALU_BoothP_4), .A1 (WindowDin_3__2__3), .S0 (
             Instr)) ;
    mux21_ni ix525 (.Y (L1FirstOperands_8__4), .A0 (
             L1_3_L2_2_G2_MINI_ALU_BoothP_5), .A1 (WindowDin_3__2__4), .S0 (
             Instr)) ;
    mux21_ni ix533 (.Y (L1FirstOperands_8__5), .A0 (
             L1_3_L2_2_G2_MINI_ALU_BoothP_6), .A1 (WindowDin_3__2__5), .S0 (
             Instr)) ;
    mux21_ni ix541 (.Y (L1FirstOperands_8__6), .A0 (
             L1_3_L2_2_G2_MINI_ALU_BoothP_7), .A1 (WindowDin_3__2__6), .S0 (
             Instr)) ;
    mux21_ni ix549 (.Y (L1FirstOperands_8__7), .A0 (
             L1_3_L2_2_G2_MINI_ALU_BoothP_8), .A1 (WindowDin_3__2__7), .S0 (
             Instr)) ;
    nor02ii ix457 (.Y (L1FirstOperands_8__8), .A0 (Instr), .A1 (
            L1_3_L2_2_G2_MINI_ALU_BoothP_9)) ;
    nor02ii ix461 (.Y (L1FirstOperands_8__9), .A0 (Instr), .A1 (
            L1_3_L2_2_G2_MINI_ALU_BoothP_10)) ;
    nor02ii ix465 (.Y (L1FirstOperands_8__10), .A0 (Instr), .A1 (
            L1_3_L2_2_G2_MINI_ALU_BoothP_11)) ;
    nor02ii ix469 (.Y (L1FirstOperands_8__11), .A0 (Instr), .A1 (
            L1_3_L2_2_G2_MINI_ALU_BoothP_12)) ;
    nor02ii ix473 (.Y (L1FirstOperands_8__12), .A0 (Instr), .A1 (
            L1_3_L2_2_G2_MINI_ALU_BoothP_13)) ;
    nor02ii ix477 (.Y (L1FirstOperands_8__13), .A0 (Instr), .A1 (
            L1_3_L2_2_G2_MINI_ALU_BoothP_14)) ;
    nor02ii ix481 (.Y (L1FirstOperands_8__14), .A0 (Instr), .A1 (
            L1_3_L2_2_G2_MINI_ALU_BoothP_15)) ;
    nor02ii ix485 (.Y (L1FirstOperands_8__15), .A0 (Instr), .A1 (
            L1_3_L2_2_G2_MINI_ALU_BoothP_16)) ;
    mux21_ni ix205 (.Y (L1FirstOperands_7__0), .A0 (
             L1_4_L2_3_G5_MINI_ALU_BoothP_1), .A1 (WindowDin_4__3__0), .S0 (
             Instr)) ;
    mux21_ni ix213 (.Y (L1FirstOperands_7__1), .A0 (
             L1_4_L2_3_G5_MINI_ALU_BoothP_2), .A1 (WindowDin_4__3__1), .S0 (
             Instr)) ;
    mux21_ni ix221 (.Y (L1FirstOperands_7__2), .A0 (
             L1_4_L2_3_G5_MINI_ALU_BoothP_3), .A1 (WindowDin_4__3__2), .S0 (
             Instr)) ;
    mux21_ni ix229 (.Y (L1FirstOperands_7__3), .A0 (
             L1_4_L2_3_G5_MINI_ALU_BoothP_4), .A1 (WindowDin_4__3__3), .S0 (
             Instr)) ;
    mux21_ni ix237 (.Y (L1FirstOperands_7__4), .A0 (
             L1_4_L2_3_G5_MINI_ALU_BoothP_5), .A1 (WindowDin_4__3__4), .S0 (
             Instr)) ;
    mux21_ni ix245 (.Y (L1FirstOperands_7__5), .A0 (
             L1_4_L2_3_G5_MINI_ALU_BoothP_6), .A1 (WindowDin_4__3__5), .S0 (
             Instr)) ;
    mux21_ni ix253 (.Y (L1FirstOperands_7__6), .A0 (
             L1_4_L2_3_G5_MINI_ALU_BoothP_7), .A1 (WindowDin_4__3__6), .S0 (
             Instr)) ;
    mux21_ni ix261 (.Y (L1FirstOperands_7__7), .A0 (
             L1_4_L2_3_G5_MINI_ALU_BoothP_8), .A1 (WindowDin_4__3__7), .S0 (
             Instr)) ;
    nor02ii ix169 (.Y (L1FirstOperands_7__8), .A0 (Instr), .A1 (
            L1_4_L2_3_G5_MINI_ALU_BoothP_9)) ;
    nor02ii ix173 (.Y (L1FirstOperands_7__9), .A0 (Instr), .A1 (
            L1_4_L2_3_G5_MINI_ALU_BoothP_10)) ;
    nor02ii ix177 (.Y (L1FirstOperands_7__10), .A0 (Instr), .A1 (
            L1_4_L2_3_G5_MINI_ALU_BoothP_11)) ;
    nor02ii ix181 (.Y (L1FirstOperands_7__11), .A0 (Instr), .A1 (
            L1_4_L2_3_G5_MINI_ALU_BoothP_12)) ;
    nor02ii ix185 (.Y (L1FirstOperands_7__12), .A0 (Instr), .A1 (
            L1_4_L2_3_G5_MINI_ALU_BoothP_13)) ;
    nor02ii ix189 (.Y (L1FirstOperands_7__13), .A0 (Instr), .A1 (
            L1_4_L2_3_G5_MINI_ALU_BoothP_14)) ;
    nor02ii ix193 (.Y (L1FirstOperands_7__14), .A0 (Instr), .A1 (
            L1_4_L2_3_G5_MINI_ALU_BoothP_15)) ;
    nor02ii ix197 (.Y (L1FirstOperands_7__15), .A0 (Instr), .A1 (
            L1_4_L2_3_G5_MINI_ALU_BoothP_16)) ;
    mux21_ni ix589 (.Y (L1FirstOperands_6__0), .A0 (
             L1_3_L2_1_G2_MINI_ALU_BoothP_1), .A1 (WindowDin_3__1__0), .S0 (
             Instr)) ;
    mux21_ni ix597 (.Y (L1FirstOperands_6__1), .A0 (
             L1_3_L2_1_G2_MINI_ALU_BoothP_2), .A1 (WindowDin_3__1__1), .S0 (
             Instr)) ;
    mux21_ni ix605 (.Y (L1FirstOperands_6__2), .A0 (
             L1_3_L2_1_G2_MINI_ALU_BoothP_3), .A1 (WindowDin_3__1__2), .S0 (
             Instr)) ;
    mux21_ni ix613 (.Y (L1FirstOperands_6__3), .A0 (
             L1_3_L2_1_G2_MINI_ALU_BoothP_4), .A1 (WindowDin_3__1__3), .S0 (
             Instr)) ;
    mux21_ni ix621 (.Y (L1FirstOperands_6__4), .A0 (
             L1_3_L2_1_G2_MINI_ALU_BoothP_5), .A1 (WindowDin_3__1__4), .S0 (
             Instr)) ;
    mux21_ni ix629 (.Y (L1FirstOperands_6__5), .A0 (
             L1_3_L2_1_G2_MINI_ALU_BoothP_6), .A1 (WindowDin_3__1__5), .S0 (
             Instr)) ;
    mux21_ni ix637 (.Y (L1FirstOperands_6__6), .A0 (
             L1_3_L2_1_G2_MINI_ALU_BoothP_7), .A1 (WindowDin_3__1__6), .S0 (
             Instr)) ;
    mux21_ni ix645 (.Y (L1FirstOperands_6__7), .A0 (
             L1_3_L2_1_G2_MINI_ALU_BoothP_8), .A1 (WindowDin_3__1__7), .S0 (
             Instr)) ;
    nor02ii ix553 (.Y (L1FirstOperands_6__8), .A0 (Instr), .A1 (
            L1_3_L2_1_G2_MINI_ALU_BoothP_9)) ;
    nor02ii ix557 (.Y (L1FirstOperands_6__9), .A0 (Instr), .A1 (
            L1_3_L2_1_G2_MINI_ALU_BoothP_10)) ;
    nor02ii ix561 (.Y (L1FirstOperands_6__10), .A0 (Instr), .A1 (
            L1_3_L2_1_G2_MINI_ALU_BoothP_11)) ;
    nor02ii ix565 (.Y (L1FirstOperands_6__11), .A0 (Instr), .A1 (
            L1_3_L2_1_G2_MINI_ALU_BoothP_12)) ;
    nor02ii ix569 (.Y (L1FirstOperands_6__12), .A0 (Instr), .A1 (
            L1_3_L2_1_G2_MINI_ALU_BoothP_13)) ;
    nor02ii ix573 (.Y (L1FirstOperands_6__13), .A0 (Instr), .A1 (
            L1_3_L2_1_G2_MINI_ALU_BoothP_14)) ;
    nor02ii ix577 (.Y (L1FirstOperands_6__14), .A0 (Instr), .A1 (
            L1_3_L2_1_G2_MINI_ALU_BoothP_15)) ;
    nor02ii ix581 (.Y (L1FirstOperands_6__15), .A0 (Instr), .A1 (
            L1_3_L2_1_G2_MINI_ALU_BoothP_16)) ;
    mux21_ni ix685 (.Y (L1FirstOperands_4__0), .A0 (
             L1_3_L2_0_G2_MINI_ALU_BoothP_1), .A1 (WindowDin_3__0__0), .S0 (
             Instr)) ;
    mux21_ni ix693 (.Y (L1FirstOperands_4__1), .A0 (
             L1_3_L2_0_G2_MINI_ALU_BoothP_2), .A1 (WindowDin_3__0__1), .S0 (
             Instr)) ;
    mux21_ni ix701 (.Y (L1FirstOperands_4__2), .A0 (
             L1_3_L2_0_G2_MINI_ALU_BoothP_3), .A1 (WindowDin_3__0__2), .S0 (
             Instr)) ;
    mux21_ni ix709 (.Y (L1FirstOperands_4__3), .A0 (
             L1_3_L2_0_G2_MINI_ALU_BoothP_4), .A1 (WindowDin_3__0__3), .S0 (
             Instr)) ;
    mux21_ni ix717 (.Y (L1FirstOperands_4__4), .A0 (
             L1_3_L2_0_G2_MINI_ALU_BoothP_5), .A1 (WindowDin_3__0__4), .S0 (
             Instr)) ;
    mux21_ni ix725 (.Y (L1FirstOperands_4__5), .A0 (
             L1_3_L2_0_G2_MINI_ALU_BoothP_6), .A1 (WindowDin_3__0__5), .S0 (
             Instr)) ;
    mux21_ni ix733 (.Y (L1FirstOperands_4__6), .A0 (
             L1_3_L2_0_G2_MINI_ALU_BoothP_7), .A1 (WindowDin_3__0__6), .S0 (
             Instr)) ;
    mux21_ni ix741 (.Y (L1FirstOperands_4__7), .A0 (
             L1_3_L2_0_G2_MINI_ALU_BoothP_8), .A1 (WindowDin_3__0__7), .S0 (
             Instr)) ;
    nor02ii ix649 (.Y (L1FirstOperands_4__8), .A0 (Instr), .A1 (
            L1_3_L2_0_G2_MINI_ALU_BoothP_9)) ;
    nor02ii ix653 (.Y (L1FirstOperands_4__9), .A0 (Instr), .A1 (
            L1_3_L2_0_G2_MINI_ALU_BoothP_10)) ;
    nor02ii ix657 (.Y (L1FirstOperands_4__10), .A0 (Instr), .A1 (
            L1_3_L2_0_G2_MINI_ALU_BoothP_11)) ;
    nor02ii ix661 (.Y (L1FirstOperands_4__11), .A0 (Instr), .A1 (
            L1_3_L2_0_G2_MINI_ALU_BoothP_12)) ;
    nor02ii ix665 (.Y (L1FirstOperands_4__12), .A0 (Instr), .A1 (
            L1_3_L2_0_G2_MINI_ALU_BoothP_13)) ;
    nor02ii ix669 (.Y (L1FirstOperands_4__13), .A0 (Instr), .A1 (
            L1_3_L2_0_G2_MINI_ALU_BoothP_14)) ;
    nor02ii ix673 (.Y (L1FirstOperands_4__14), .A0 (Instr), .A1 (
            L1_3_L2_0_G2_MINI_ALU_BoothP_15)) ;
    nor02ii ix677 (.Y (L1FirstOperands_4__15), .A0 (Instr), .A1 (
            L1_3_L2_0_G2_MINI_ALU_BoothP_16)) ;
    mux21_ni ix301 (.Y (L1FirstOperands_3__0), .A0 (
             L1_4_L2_2_G4_MINI_ALU_BoothP_1), .A1 (WindowDin_4__2__0), .S0 (
             Instr)) ;
    mux21_ni ix309 (.Y (L1FirstOperands_3__1), .A0 (
             L1_4_L2_2_G4_MINI_ALU_BoothP_2), .A1 (WindowDin_4__2__1), .S0 (
             Instr)) ;
    mux21_ni ix317 (.Y (L1FirstOperands_3__2), .A0 (
             L1_4_L2_2_G4_MINI_ALU_BoothP_3), .A1 (WindowDin_4__2__2), .S0 (
             Instr)) ;
    mux21_ni ix325 (.Y (L1FirstOperands_3__3), .A0 (
             L1_4_L2_2_G4_MINI_ALU_BoothP_4), .A1 (WindowDin_4__2__3), .S0 (
             Instr)) ;
    mux21_ni ix333 (.Y (L1FirstOperands_3__4), .A0 (
             L1_4_L2_2_G4_MINI_ALU_BoothP_5), .A1 (WindowDin_4__2__4), .S0 (
             Instr)) ;
    mux21_ni ix341 (.Y (L1FirstOperands_3__5), .A0 (
             L1_4_L2_2_G4_MINI_ALU_BoothP_6), .A1 (WindowDin_4__2__5), .S0 (
             Instr)) ;
    mux21_ni ix349 (.Y (L1FirstOperands_3__6), .A0 (
             L1_4_L2_2_G4_MINI_ALU_BoothP_7), .A1 (WindowDin_4__2__6), .S0 (
             Instr)) ;
    mux21_ni ix357 (.Y (L1FirstOperands_3__7), .A0 (
             L1_4_L2_2_G4_MINI_ALU_BoothP_8), .A1 (WindowDin_4__2__7), .S0 (
             Instr)) ;
    nor02ii ix265 (.Y (L1FirstOperands_3__8), .A0 (Instr), .A1 (
            L1_4_L2_2_G4_MINI_ALU_BoothP_9)) ;
    nor02ii ix269 (.Y (L1FirstOperands_3__9), .A0 (Instr), .A1 (
            L1_4_L2_2_G4_MINI_ALU_BoothP_10)) ;
    nor02ii ix273 (.Y (L1FirstOperands_3__10), .A0 (Instr), .A1 (
            L1_4_L2_2_G4_MINI_ALU_BoothP_11)) ;
    nor02ii ix277 (.Y (L1FirstOperands_3__11), .A0 (Instr), .A1 (
            L1_4_L2_2_G4_MINI_ALU_BoothP_12)) ;
    nor02ii ix281 (.Y (L1FirstOperands_3__12), .A0 (Instr), .A1 (
            L1_4_L2_2_G4_MINI_ALU_BoothP_13)) ;
    nor02ii ix285 (.Y (L1FirstOperands_3__13), .A0 (Instr), .A1 (
            L1_4_L2_2_G4_MINI_ALU_BoothP_14)) ;
    nor02ii ix289 (.Y (L1FirstOperands_3__14), .A0 (Instr), .A1 (
            L1_4_L2_2_G4_MINI_ALU_BoothP_15)) ;
    nor02ii ix293 (.Y (L1FirstOperands_3__15), .A0 (Instr), .A1 (
            L1_4_L2_2_G4_MINI_ALU_BoothP_16)) ;
    mux21_ni ix781 (.Y (L1FirstOperands_2__0), .A0 (
             L1_2_L2_4_G2_MINI_ALU_BoothP_1), .A1 (WindowDin_2__4__0), .S0 (
             Instr)) ;
    mux21_ni ix789 (.Y (L1FirstOperands_2__1), .A0 (
             L1_2_L2_4_G2_MINI_ALU_BoothP_2), .A1 (WindowDin_2__4__1), .S0 (
             Instr)) ;
    mux21_ni ix797 (.Y (L1FirstOperands_2__2), .A0 (
             L1_2_L2_4_G2_MINI_ALU_BoothP_3), .A1 (WindowDin_2__4__2), .S0 (
             Instr)) ;
    mux21_ni ix805 (.Y (L1FirstOperands_2__3), .A0 (
             L1_2_L2_4_G2_MINI_ALU_BoothP_4), .A1 (WindowDin_2__4__3), .S0 (
             Instr)) ;
    mux21_ni ix813 (.Y (L1FirstOperands_2__4), .A0 (
             L1_2_L2_4_G2_MINI_ALU_BoothP_5), .A1 (WindowDin_2__4__4), .S0 (
             Instr)) ;
    mux21_ni ix821 (.Y (L1FirstOperands_2__5), .A0 (
             L1_2_L2_4_G2_MINI_ALU_BoothP_6), .A1 (WindowDin_2__4__5), .S0 (
             Instr)) ;
    mux21_ni ix829 (.Y (L1FirstOperands_2__6), .A0 (
             L1_2_L2_4_G2_MINI_ALU_BoothP_7), .A1 (WindowDin_2__4__6), .S0 (
             Instr)) ;
    mux21_ni ix837 (.Y (L1FirstOperands_2__7), .A0 (
             L1_2_L2_4_G2_MINI_ALU_BoothP_8), .A1 (WindowDin_2__4__7), .S0 (
             Instr)) ;
    nor02ii ix745 (.Y (L1FirstOperands_2__8), .A0 (Instr), .A1 (
            L1_2_L2_4_G2_MINI_ALU_BoothP_9)) ;
    nor02ii ix749 (.Y (L1FirstOperands_2__9), .A0 (Instr), .A1 (
            L1_2_L2_4_G2_MINI_ALU_BoothP_10)) ;
    nor02ii ix753 (.Y (L1FirstOperands_2__10), .A0 (Instr), .A1 (
            L1_2_L2_4_G2_MINI_ALU_BoothP_11)) ;
    nor02ii ix757 (.Y (L1FirstOperands_2__11), .A0 (Instr), .A1 (
            L1_2_L2_4_G2_MINI_ALU_BoothP_12)) ;
    nor02ii ix761 (.Y (L1FirstOperands_2__12), .A0 (Instr), .A1 (
            L1_2_L2_4_G2_MINI_ALU_BoothP_13)) ;
    nor02ii ix765 (.Y (L1FirstOperands_2__13), .A0 (Instr), .A1 (
            L1_2_L2_4_G2_MINI_ALU_BoothP_14)) ;
    nor02ii ix769 (.Y (L1FirstOperands_2__14), .A0 (Instr), .A1 (
            L1_2_L2_4_G2_MINI_ALU_BoothP_15)) ;
    nor02ii ix773 (.Y (L1FirstOperands_2__15), .A0 (Instr), .A1 (
            L1_2_L2_4_G2_MINI_ALU_BoothP_16)) ;
    mux21_ni ix877 (.Y (L1FirstOperands_0__0), .A0 (
             L1_2_L2_3_G2_MINI_ALU_BoothP_1), .A1 (WindowDin_2__3__0), .S0 (
             Instr)) ;
    mux21_ni ix885 (.Y (L1FirstOperands_0__1), .A0 (
             L1_2_L2_3_G2_MINI_ALU_BoothP_2), .A1 (WindowDin_2__3__1), .S0 (
             Instr)) ;
    mux21_ni ix893 (.Y (L1FirstOperands_0__2), .A0 (
             L1_2_L2_3_G2_MINI_ALU_BoothP_3), .A1 (WindowDin_2__3__2), .S0 (
             Instr)) ;
    mux21_ni ix901 (.Y (L1FirstOperands_0__3), .A0 (
             L1_2_L2_3_G2_MINI_ALU_BoothP_4), .A1 (WindowDin_2__3__3), .S0 (
             Instr)) ;
    mux21_ni ix909 (.Y (L1FirstOperands_0__4), .A0 (
             L1_2_L2_3_G2_MINI_ALU_BoothP_5), .A1 (WindowDin_2__3__4), .S0 (
             Instr)) ;
    mux21_ni ix917 (.Y (L1FirstOperands_0__5), .A0 (
             L1_2_L2_3_G2_MINI_ALU_BoothP_6), .A1 (WindowDin_2__3__5), .S0 (
             Instr)) ;
    mux21_ni ix925 (.Y (L1FirstOperands_0__6), .A0 (
             L1_2_L2_3_G2_MINI_ALU_BoothP_7), .A1 (WindowDin_2__3__6), .S0 (
             Instr)) ;
    mux21_ni ix933 (.Y (L1FirstOperands_0__7), .A0 (
             L1_2_L2_3_G2_MINI_ALU_BoothP_8), .A1 (WindowDin_2__3__7), .S0 (
             Instr)) ;
    nor02ii ix841 (.Y (L1FirstOperands_0__8), .A0 (Instr), .A1 (
            L1_2_L2_3_G2_MINI_ALU_BoothP_9)) ;
    nor02ii ix845 (.Y (L1FirstOperands_0__9), .A0 (Instr), .A1 (
            L1_2_L2_3_G2_MINI_ALU_BoothP_10)) ;
    nor02ii ix849 (.Y (L1FirstOperands_0__10), .A0 (Instr), .A1 (
            L1_2_L2_3_G2_MINI_ALU_BoothP_11)) ;
    nor02ii ix853 (.Y (L1FirstOperands_0__11), .A0 (Instr), .A1 (
            L1_2_L2_3_G2_MINI_ALU_BoothP_12)) ;
    nor02ii ix857 (.Y (L1FirstOperands_0__12), .A0 (Instr), .A1 (
            L1_2_L2_3_G2_MINI_ALU_BoothP_13)) ;
    nor02ii ix861 (.Y (L1FirstOperands_0__13), .A0 (Instr), .A1 (
            L1_2_L2_3_G2_MINI_ALU_BoothP_14)) ;
    nor02ii ix865 (.Y (L1FirstOperands_0__14), .A0 (Instr), .A1 (
            L1_2_L2_3_G2_MINI_ALU_BoothP_15)) ;
    nor02ii ix869 (.Y (L1FirstOperands_0__15), .A0 (Instr), .A1 (
            L1_2_L2_3_G2_MINI_ALU_BoothP_16)) ;
    nor02ii ix2243 (.Y (LoopingAndResultNotReady), .A0 (nx3233), .A1 (nx2856)) ;
    nor04 ix3234 (.Y (nx3233), .A0 (CounterOut_0), .A1 (CounterOut_1), .A2 (
          CounterOut_2), .A3 (CounterOut_3)) ;
    oai21 ix29 (.Y (Result[0]), .A0 (nx3236), .A1 (Instr), .B0 (nx3238)) ;
    inv01 ix3237 (.Y (nx3236), .A (L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_0)) ;
    aoi32 ix3239 (.Y (nx3238), .A0 (L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_5), .A1 (
          FilterSize), .A2 (Instr), .B0 (
          L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_3), .B1 (nx22)) ;
    nor02ii ix23 (.Y (nx22), .A0 (FilterSize), .A1 (Instr)) ;
    oai21 ix41 (.Y (Result[1]), .A0 (nx3242), .A1 (Instr), .B0 (nx3244)) ;
    inv01 ix3243 (.Y (nx3242), .A (L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_1)) ;
    aoi32 ix3245 (.Y (nx3244), .A0 (L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_6), .A1 (
          FilterSize), .A2 (Instr), .B0 (
          L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_4), .B1 (nx22)) ;
    oai21 ix53 (.Y (Result[2]), .A0 (nx3247), .A1 (Instr), .B0 (nx3249)) ;
    inv01 ix3248 (.Y (nx3247), .A (L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_2)) ;
    aoi32 ix3250 (.Y (nx3249), .A0 (L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_7), .A1 (
          FilterSize), .A2 (Instr), .B0 (
          L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_5), .B1 (nx22)) ;
    nor02ii ix3 (.Y (Result[5]), .A0 (Instr), .A1 (
            L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_5)) ;
    nor02ii ix7 (.Y (Result[6]), .A0 (Instr), .A1 (
            L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_6)) ;
    nor02ii ix11 (.Y (Result[7]), .A0 (Instr), .A1 (
            L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_7)) ;
    inv01 ix1079 (.Y (Done), .A (NOT__13497)) ;
    inv01 ix3272 (.Y (nx3273), .A (LoopingAndResultNotReady)) ;
    inv01 ix3274 (.Y (nx3275), .A (nx3273)) ;
    inv01 ix3276 (.Y (nx3277), .A (nx3273)) ;
    inv01 ix3278 (.Y (nx3279), .A (nx3273)) ;
    inv01 ix3280 (.Y (nx3281), .A (nx3273)) ;
    inv01 ix3282 (.Y (nx3283), .A (Done)) ;
    inv01 ix3284 (.Y (nx3285), .A (Done)) ;
    inv01 ix3286 (.Y (nx3287), .A (Done)) ;
    inv01 ix3288 (.Y (nx3289), .A (Done)) ;
    and02 ix1033 (.Y (nx1032), .A0 (NOT__13497), .A1 (CLK)) ;
    or02 ix2873 (.Y (nx2872), .A0 (nx2876), .A1 (NOT_CounterOut_0)) ;
    xnor2 ix1047 (.Y (nx1046), .A0 (nx2876), .A1 (CounterOut_0)) ;
    ao22 ix61 (.Y (Result[3]), .A0 (L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_6), .A1 (
         nx22), .B0 (L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_3), .B1 (nx3303)) ;
    inv01 ix3302 (.Y (nx3303), .A (Instr)) ;
    ao22 ix69 (.Y (Result[4]), .A0 (L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_7), .A1 (
         nx22), .B0 (L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_4), .B1 (nx3303)) ;
    latchr ACCELERATOR_COUNTER_lat_Dout_0__u1 (.QB (nx5), .D (NOT_CounterOut_0)
           , .CLK (nx1032), .R (nx1036)) ;
    inv01 ACCELERATOR_COUNTER_lat_Dout_0__u2 (.Y (CounterOut_0), .A (nx5)) ;
    buf02 ACCELERATOR_COUNTER_lat_Dout_0__u3 (.Y (NOT_CounterOut_0), .A (nx5)) ;
    latchr ACCELERATOR_COUNTER_lat_Dout_3__u1 (.QB (nx3304), .D (nx1066), .CLK (
           nx1032), .R (nx1036)) ;
    inv01 ACCELERATOR_COUNTER_lat_Dout_3__u2 (.Y (CounterOut_3), .A (nx3304)) ;
    buf02 ACCELERATOR_COUNTER_lat_Dout_3__u3 (.Y (nx1), .A (nx3304)) ;
    latchr ACCELERATOR_COUNTER_lat_Dout_2__u1 (.QB (nx3306), .D (nx1058), .CLK (
           nx1032), .R (nx1036)) ;
    inv01 ACCELERATOR_COUNTER_lat_Dout_2__u2 (.Y (CounterOut_2), .A (nx3306)) ;
    buf02 ACCELERATOR_COUNTER_lat_Dout_2__u3 (.Y (nx3305), .A (nx3306)) ;
    latchr ACCELERATOR_COUNTER_lat_Dout_1__u1 (.QB (nx3308), .D (nx1046), .CLK (
           nx1032), .R (nx1036)) ;
    inv01 ACCELERATOR_COUNTER_lat_Dout_1__u2 (.Y (CounterOut_1), .A (nx3308)) ;
    buf02 ACCELERATOR_COUNTER_lat_Dout_1__u3 (.Y (nx2876), .A (nx3308)) ;
endmodule


module booth_adder_17_unfolded5 ( AdderFirstOperand, AdderSecondOperand, 
                                  BoothOperand, BoothP, SelOperand, Operation, 
                                  AdderResult, AdderBoothResult ) ;

    input [16:0]AdderFirstOperand ;
    input [16:0]AdderSecondOperand ;
    input [16:0]BoothOperand ;
    input [16:0]BoothP ;
    input SelOperand ;
    input Operation ;
    output [16:0]AdderResult ;
    output [16:0]AdderBoothResult ;

    wire AdderResult_16_rename, AdderResult_15_rename, AdderResult_14_rename, 
         AdderResult_13_rename, AdderResult_12_rename, AdderResult_11_rename, 
         AdderResult_10_rename, AdderResult_9_rename, AdderResult_8_rename, 
         FirstOperand_16, FirstOperand_15, FirstOperand_14, FirstOperand_13, 
         FirstOperand_12, FirstOperand_11, FirstOperand_10, FirstOperand_9, 
         FirstOperand_8, FirstOperand_7, FirstOperand_6, FirstOperand_5, 
         FirstOperand_4, FirstOperand_3, FirstOperand_2, FirstOperand_1, 
         FirstOperand_0, SecondOperand_16, SecondOperand_15, SecondOperand_14, 
         SecondOperand_13, SecondOperand_12, SecondOperand_11, SecondOperand_10, 
         SecondOperand_9, SecondOperand_8, SecondOperand_7, SecondOperand_6, 
         SecondOperand_5, SecondOperand_4, SecondOperand_3, SecondOperand_2, 
         SecondOperand_1, SecondOperand_0, nx224, nx227, nx229, nx231, nx233, 
         nx235, nx237, nx239, nx241, nx243;
    wire [0:0] \$dummy ;




    assign AdderResult[16] = AdderBoothResult[16] ;
    assign AdderResult[15] = AdderBoothResult[16] ;
    assign AdderResult[14] = AdderBoothResult[16] ;
    assign AdderResult[13] = AdderBoothResult[16] ;
    assign AdderResult[12] = AdderBoothResult[16] ;
    assign AdderResult[11] = AdderBoothResult[16] ;
    assign AdderResult[10] = AdderBoothResult[16] ;
    assign AdderResult[9] = AdderBoothResult[16] ;
    assign AdderResult[8] = AdderBoothResult[16] ;
    adder_17 ADDER (.A ({FirstOperand_16,FirstOperand_15,FirstOperand_14,
             FirstOperand_13,FirstOperand_12,FirstOperand_11,FirstOperand_10,
             FirstOperand_9,FirstOperand_8,FirstOperand_7,FirstOperand_6,
             FirstOperand_5,FirstOperand_4,FirstOperand_3,FirstOperand_2,
             FirstOperand_1,FirstOperand_0}), .B ({SecondOperand_16,
             SecondOperand_15,SecondOperand_14,SecondOperand_13,SecondOperand_12
             ,SecondOperand_11,SecondOperand_10,SecondOperand_9,SecondOperand_8,
             SecondOperand_7,SecondOperand_6,SecondOperand_5,SecondOperand_4,
             SecondOperand_3,SecondOperand_2,SecondOperand_1,SecondOperand_0}), 
             .Cin (AdderBoothResult[16]), .Sum ({AdderResult_16_rename,
             AdderResult_15_rename,AdderResult_14_rename,AdderResult_13_rename,
             AdderResult_12_rename,AdderResult_11_rename,AdderResult_10_rename,
             AdderResult_9_rename,AdderResult_8_rename,AdderResult[7],
             AdderResult[6],AdderResult[5],AdderResult[4],AdderResult[3],
             AdderResult[2],AdderResult[1],AdderResult[0]}), .Cout (\$dummy [0])
             ) ;
    fake_gnd ix47 (.Y (AdderBoothResult[16])) ;
    mux21_ni ix137 (.Y (SecondOperand_0), .A0 (AdderSecondOperand[0]), .A1 (
             BoothP[0]), .S0 (nx235)) ;
    mux21_ni ix145 (.Y (SecondOperand_1), .A0 (AdderSecondOperand[1]), .A1 (
             BoothP[1]), .S0 (nx235)) ;
    mux21_ni ix153 (.Y (SecondOperand_2), .A0 (AdderSecondOperand[2]), .A1 (
             BoothP[2]), .S0 (nx235)) ;
    mux21_ni ix161 (.Y (SecondOperand_3), .A0 (AdderSecondOperand[3]), .A1 (
             BoothP[3]), .S0 (nx235)) ;
    mux21_ni ix169 (.Y (SecondOperand_4), .A0 (AdderSecondOperand[4]), .A1 (
             BoothP[4]), .S0 (nx235)) ;
    mux21_ni ix177 (.Y (SecondOperand_5), .A0 (AdderSecondOperand[5]), .A1 (
             BoothP[5]), .S0 (nx235)) ;
    mux21_ni ix185 (.Y (SecondOperand_6), .A0 (AdderSecondOperand[6]), .A1 (
             BoothP[6]), .S0 (nx235)) ;
    mux21_ni ix193 (.Y (SecondOperand_7), .A0 (AdderSecondOperand[7]), .A1 (
             BoothP[7]), .S0 (nx237)) ;
    mux21_ni ix201 (.Y (SecondOperand_8), .A0 (AdderSecondOperand[8]), .A1 (
             BoothP[8]), .S0 (nx237)) ;
    mux21_ni ix209 (.Y (SecondOperand_9), .A0 (AdderSecondOperand[9]), .A1 (
             BoothP[9]), .S0 (nx237)) ;
    mux21_ni ix217 (.Y (SecondOperand_10), .A0 (AdderSecondOperand[10]), .A1 (
             BoothP[10]), .S0 (nx237)) ;
    mux21_ni ix225 (.Y (SecondOperand_11), .A0 (AdderSecondOperand[11]), .A1 (
             BoothP[11]), .S0 (nx237)) ;
    mux21_ni ix233 (.Y (SecondOperand_12), .A0 (AdderSecondOperand[12]), .A1 (
             BoothP[12]), .S0 (nx237)) ;
    mux21_ni ix241 (.Y (SecondOperand_13), .A0 (AdderSecondOperand[13]), .A1 (
             BoothP[13]), .S0 (nx237)) ;
    mux21_ni ix249 (.Y (SecondOperand_14), .A0 (AdderSecondOperand[14]), .A1 (
             BoothP[14]), .S0 (nx239)) ;
    mux21_ni ix257 (.Y (SecondOperand_15), .A0 (AdderSecondOperand[15]), .A1 (
             BoothP[15]), .S0 (nx239)) ;
    nor02ii ix261 (.Y (FirstOperand_0), .A0 (nx239), .A1 (AdderFirstOperand[0])
            ) ;
    nor02ii ix265 (.Y (FirstOperand_1), .A0 (nx239), .A1 (AdderFirstOperand[1])
            ) ;
    nor02ii ix269 (.Y (FirstOperand_2), .A0 (nx239), .A1 (AdderFirstOperand[2])
            ) ;
    nor02ii ix273 (.Y (FirstOperand_3), .A0 (nx239), .A1 (AdderFirstOperand[3])
            ) ;
    nor02ii ix277 (.Y (FirstOperand_4), .A0 (nx239), .A1 (AdderFirstOperand[4])
            ) ;
    nor02ii ix281 (.Y (FirstOperand_5), .A0 (nx241), .A1 (AdderFirstOperand[5])
            ) ;
    nor02ii ix285 (.Y (FirstOperand_6), .A0 (nx241), .A1 (AdderFirstOperand[6])
            ) ;
    nor02ii ix289 (.Y (FirstOperand_7), .A0 (nx241), .A1 (AdderFirstOperand[7])
            ) ;
    nor02ii ix293 (.Y (FirstOperand_8), .A0 (nx241), .A1 (AdderFirstOperand[8])
            ) ;
    mux21_ni ix301 (.Y (FirstOperand_9), .A0 (AdderFirstOperand[9]), .A1 (
             BoothOperand[9]), .S0 (nx241)) ;
    mux21_ni ix309 (.Y (FirstOperand_10), .A0 (AdderFirstOperand[10]), .A1 (
             BoothOperand[10]), .S0 (nx241)) ;
    mux21_ni ix317 (.Y (FirstOperand_11), .A0 (AdderFirstOperand[11]), .A1 (
             BoothOperand[11]), .S0 (nx241)) ;
    mux21_ni ix325 (.Y (FirstOperand_12), .A0 (AdderFirstOperand[12]), .A1 (
             BoothOperand[12]), .S0 (nx243)) ;
    mux21_ni ix333 (.Y (FirstOperand_13), .A0 (AdderFirstOperand[13]), .A1 (
             BoothOperand[13]), .S0 (nx243)) ;
    mux21_ni ix341 (.Y (FirstOperand_14), .A0 (AdderFirstOperand[14]), .A1 (
             BoothOperand[14]), .S0 (nx243)) ;
    mux21_ni ix349 (.Y (FirstOperand_15), .A0 (AdderFirstOperand[15]), .A1 (
             BoothOperand[15]), .S0 (nx243)) ;
    mux21_ni ix357 (.Y (FirstOperand_16), .A0 (AdderFirstOperand[16]), .A1 (
             BoothOperand[16]), .S0 (nx243)) ;
    mux21_ni ix7 (.Y (AdderBoothResult[0]), .A0 (BoothP[1]), .A1 (AdderResult[1]
             ), .S0 (nx227)) ;
    mux21_ni ix15 (.Y (AdderBoothResult[1]), .A0 (BoothP[2]), .A1 (
             AdderResult[2]), .S0 (nx227)) ;
    mux21_ni ix23 (.Y (AdderBoothResult[2]), .A0 (BoothP[3]), .A1 (
             AdderResult[3]), .S0 (nx227)) ;
    mux21_ni ix31 (.Y (AdderBoothResult[3]), .A0 (BoothP[4]), .A1 (
             AdderResult[4]), .S0 (nx227)) ;
    mux21_ni ix39 (.Y (AdderBoothResult[4]), .A0 (BoothP[5]), .A1 (
             AdderResult[5]), .S0 (nx227)) ;
    mux21_ni ix49 (.Y (AdderBoothResult[5]), .A0 (BoothP[6]), .A1 (
             AdderResult[6]), .S0 (nx227)) ;
    mux21_ni ix55 (.Y (AdderBoothResult[6]), .A0 (BoothP[7]), .A1 (
             AdderResult[7]), .S0 (nx227)) ;
    mux21_ni ix63 (.Y (AdderBoothResult[7]), .A0 (BoothP[8]), .A1 (
             AdderResult_8_rename), .S0 (nx229)) ;
    mux21_ni ix71 (.Y (AdderBoothResult[8]), .A0 (BoothP[9]), .A1 (
             AdderResult_9_rename), .S0 (nx229)) ;
    mux21_ni ix79 (.Y (AdderBoothResult[9]), .A0 (BoothP[10]), .A1 (
             AdderResult_10_rename), .S0 (nx229)) ;
    mux21_ni ix87 (.Y (AdderBoothResult[10]), .A0 (BoothP[11]), .A1 (
             AdderResult_11_rename), .S0 (nx229)) ;
    mux21_ni ix95 (.Y (AdderBoothResult[11]), .A0 (BoothP[12]), .A1 (
             AdderResult_12_rename), .S0 (nx229)) ;
    mux21_ni ix103 (.Y (AdderBoothResult[12]), .A0 (BoothP[13]), .A1 (
             AdderResult_13_rename), .S0 (nx229)) ;
    mux21_ni ix111 (.Y (AdderBoothResult[13]), .A0 (BoothP[14]), .A1 (
             AdderResult_14_rename), .S0 (nx229)) ;
    mux21_ni ix119 (.Y (AdderBoothResult[14]), .A0 (BoothP[15]), .A1 (
             AdderResult_15_rename), .S0 (nx231)) ;
    mux21_ni ix127 (.Y (AdderBoothResult[15]), .A0 (BoothP[16]), .A1 (
             AdderResult_16_rename), .S0 (nx231)) ;
    and02 ix129 (.Y (SecondOperand_16), .A0 (nx243), .A1 (BoothP[16])) ;
    inv01 ix223 (.Y (nx224), .A (Operation)) ;
    inv02 ix226 (.Y (nx227), .A (nx224)) ;
    inv02 ix228 (.Y (nx229), .A (nx224)) ;
    inv02 ix230 (.Y (nx231), .A (nx224)) ;
    inv01 ix232 (.Y (nx233), .A (SelOperand)) ;
    inv02 ix234 (.Y (nx235), .A (nx233)) ;
    inv02 ix236 (.Y (nx237), .A (nx233)) ;
    inv02 ix238 (.Y (nx239), .A (nx233)) ;
    inv02 ix240 (.Y (nx241), .A (nx233)) ;
    inv02 ix242 (.Y (nx243), .A (nx233)) ;
endmodule


module booth_adder_17_unfolded4 ( AdderFirstOperand, AdderSecondOperand, 
                                  BoothOperand, BoothP, SelOperand, Operation, 
                                  AdderResult, AdderBoothResult ) ;

    input [16:0]AdderFirstOperand ;
    input [16:0]AdderSecondOperand ;
    input [16:0]BoothOperand ;
    input [16:0]BoothP ;
    input SelOperand ;
    input Operation ;
    output [16:0]AdderResult ;
    output [16:0]AdderBoothResult ;

    wire FirstOperand_16, FirstOperand_15, FirstOperand_14, FirstOperand_13, 
         FirstOperand_12, FirstOperand_11, FirstOperand_10, FirstOperand_9, 
         FirstOperand_8, FirstOperand_7, FirstOperand_6, FirstOperand_5, 
         FirstOperand_4, FirstOperand_3, FirstOperand_2, FirstOperand_1, 
         FirstOperand_0, SecondOperand_16, SecondOperand_15, SecondOperand_14, 
         SecondOperand_13, SecondOperand_12, SecondOperand_11, SecondOperand_10, 
         SecondOperand_9, SecondOperand_8, SecondOperand_7, SecondOperand_6, 
         SecondOperand_5, SecondOperand_4, SecondOperand_3, SecondOperand_2, 
         SecondOperand_1, SecondOperand_0, nx220, nx222, nx225, nx227, nx229, 
         nx231, nx233, nx235, nx237, nx239;
    wire [0:0] \$dummy ;




    adder_17 ADDER (.A ({FirstOperand_16,FirstOperand_15,FirstOperand_14,
             FirstOperand_13,FirstOperand_12,FirstOperand_11,FirstOperand_10,
             FirstOperand_9,FirstOperand_8,FirstOperand_7,FirstOperand_6,
             FirstOperand_5,FirstOperand_4,FirstOperand_3,FirstOperand_2,
             FirstOperand_1,FirstOperand_0}), .B ({SecondOperand_16,
             SecondOperand_15,SecondOperand_14,SecondOperand_13,SecondOperand_12
             ,SecondOperand_11,SecondOperand_10,SecondOperand_9,SecondOperand_8,
             SecondOperand_7,SecondOperand_6,SecondOperand_5,SecondOperand_4,
             SecondOperand_3,SecondOperand_2,SecondOperand_1,SecondOperand_0}), 
             .Cin (AdderBoothResult[16]), .Sum ({AdderResult[16],AdderResult[15]
             ,AdderResult[14],AdderResult[13],AdderResult[12],AdderResult[11],
             AdderResult[10],AdderResult[9],AdderResult[8],AdderResult[7],
             AdderResult[6],AdderResult[5],AdderResult[4],AdderResult[3],
             AdderResult[2],AdderResult[1],AdderResult[0]}), .Cout (\$dummy [0])
             ) ;
    fake_gnd ix45 (.Y (AdderBoothResult[16])) ;
    mux21_ni ix135 (.Y (SecondOperand_0), .A0 (AdderSecondOperand[0]), .A1 (
             BoothP[0]), .S0 (nx231)) ;
    mux21_ni ix143 (.Y (SecondOperand_1), .A0 (AdderSecondOperand[1]), .A1 (
             BoothP[1]), .S0 (nx231)) ;
    mux21_ni ix151 (.Y (SecondOperand_2), .A0 (AdderSecondOperand[2]), .A1 (
             BoothP[2]), .S0 (nx231)) ;
    mux21_ni ix159 (.Y (SecondOperand_3), .A0 (AdderSecondOperand[3]), .A1 (
             BoothP[3]), .S0 (nx231)) ;
    mux21_ni ix167 (.Y (SecondOperand_4), .A0 (AdderSecondOperand[4]), .A1 (
             BoothP[4]), .S0 (nx231)) ;
    mux21_ni ix175 (.Y (SecondOperand_5), .A0 (AdderSecondOperand[5]), .A1 (
             BoothP[5]), .S0 (nx231)) ;
    mux21_ni ix183 (.Y (SecondOperand_6), .A0 (AdderSecondOperand[6]), .A1 (
             BoothP[6]), .S0 (nx231)) ;
    mux21_ni ix191 (.Y (SecondOperand_7), .A0 (AdderSecondOperand[7]), .A1 (
             BoothP[7]), .S0 (nx233)) ;
    mux21_ni ix199 (.Y (SecondOperand_8), .A0 (AdderSecondOperand[8]), .A1 (
             BoothP[8]), .S0 (nx233)) ;
    mux21_ni ix207 (.Y (SecondOperand_9), .A0 (AdderSecondOperand[9]), .A1 (
             BoothP[9]), .S0 (nx233)) ;
    mux21_ni ix215 (.Y (SecondOperand_10), .A0 (AdderSecondOperand[10]), .A1 (
             BoothP[10]), .S0 (nx233)) ;
    mux21_ni ix223 (.Y (SecondOperand_11), .A0 (AdderSecondOperand[11]), .A1 (
             BoothP[11]), .S0 (nx233)) ;
    mux21_ni ix231 (.Y (SecondOperand_12), .A0 (AdderSecondOperand[12]), .A1 (
             BoothP[12]), .S0 (nx233)) ;
    mux21_ni ix239 (.Y (SecondOperand_13), .A0 (AdderSecondOperand[13]), .A1 (
             BoothP[13]), .S0 (nx233)) ;
    mux21_ni ix247 (.Y (SecondOperand_14), .A0 (AdderSecondOperand[14]), .A1 (
             BoothP[14]), .S0 (nx235)) ;
    mux21_ni ix255 (.Y (SecondOperand_15), .A0 (AdderSecondOperand[15]), .A1 (
             BoothP[15]), .S0 (nx235)) ;
    mux21_ni ix263 (.Y (SecondOperand_16), .A0 (AdderSecondOperand[16]), .A1 (
             BoothP[16]), .S0 (nx235)) ;
    nor02ii ix267 (.Y (FirstOperand_0), .A0 (nx235), .A1 (AdderFirstOperand[0])
            ) ;
    nor02ii ix271 (.Y (FirstOperand_1), .A0 (nx235), .A1 (AdderFirstOperand[1])
            ) ;
    nor02ii ix275 (.Y (FirstOperand_2), .A0 (nx235), .A1 (AdderFirstOperand[2])
            ) ;
    nor02ii ix279 (.Y (FirstOperand_3), .A0 (nx235), .A1 (AdderFirstOperand[3])
            ) ;
    nor02ii ix283 (.Y (FirstOperand_4), .A0 (nx237), .A1 (AdderFirstOperand[4])
            ) ;
    nor02ii ix287 (.Y (FirstOperand_5), .A0 (nx237), .A1 (AdderFirstOperand[5])
            ) ;
    nor02ii ix291 (.Y (FirstOperand_6), .A0 (nx237), .A1 (AdderFirstOperand[6])
            ) ;
    nor02ii ix295 (.Y (FirstOperand_7), .A0 (nx237), .A1 (AdderFirstOperand[7])
            ) ;
    nor02ii ix299 (.Y (FirstOperand_8), .A0 (nx237), .A1 (AdderFirstOperand[8])
            ) ;
    mux21_ni ix307 (.Y (FirstOperand_9), .A0 (AdderFirstOperand[9]), .A1 (
             BoothOperand[9]), .S0 (nx237)) ;
    mux21_ni ix315 (.Y (FirstOperand_10), .A0 (AdderFirstOperand[10]), .A1 (
             BoothOperand[10]), .S0 (nx237)) ;
    mux21_ni ix323 (.Y (FirstOperand_11), .A0 (AdderFirstOperand[11]), .A1 (
             BoothOperand[11]), .S0 (nx239)) ;
    mux21_ni ix331 (.Y (FirstOperand_12), .A0 (AdderFirstOperand[12]), .A1 (
             BoothOperand[12]), .S0 (nx239)) ;
    mux21_ni ix339 (.Y (FirstOperand_13), .A0 (AdderFirstOperand[13]), .A1 (
             BoothOperand[13]), .S0 (nx239)) ;
    mux21_ni ix347 (.Y (FirstOperand_14), .A0 (AdderFirstOperand[14]), .A1 (
             BoothOperand[14]), .S0 (nx239)) ;
    mux21_ni ix355 (.Y (FirstOperand_15), .A0 (AdderFirstOperand[15]), .A1 (
             BoothOperand[15]), .S0 (nx239)) ;
    mux21_ni ix363 (.Y (FirstOperand_16), .A0 (AdderFirstOperand[16]), .A1 (
             BoothOperand[16]), .S0 (nx239)) ;
    mux21_ni ix7 (.Y (AdderBoothResult[0]), .A0 (BoothP[1]), .A1 (AdderResult[1]
             ), .S0 (nx222)) ;
    mux21_ni ix15 (.Y (AdderBoothResult[1]), .A0 (BoothP[2]), .A1 (
             AdderResult[2]), .S0 (nx222)) ;
    mux21_ni ix23 (.Y (AdderBoothResult[2]), .A0 (BoothP[3]), .A1 (
             AdderResult[3]), .S0 (nx222)) ;
    mux21_ni ix31 (.Y (AdderBoothResult[3]), .A0 (BoothP[4]), .A1 (
             AdderResult[4]), .S0 (nx222)) ;
    mux21_ni ix39 (.Y (AdderBoothResult[4]), .A0 (BoothP[5]), .A1 (
             AdderResult[5]), .S0 (nx222)) ;
    mux21_ni ix48 (.Y (AdderBoothResult[5]), .A0 (BoothP[6]), .A1 (
             AdderResult[6]), .S0 (nx222)) ;
    mux21_ni ix55 (.Y (AdderBoothResult[6]), .A0 (BoothP[7]), .A1 (
             AdderResult[7]), .S0 (nx222)) ;
    mux21_ni ix63 (.Y (AdderBoothResult[7]), .A0 (BoothP[8]), .A1 (
             AdderResult[8]), .S0 (nx225)) ;
    mux21_ni ix71 (.Y (AdderBoothResult[8]), .A0 (BoothP[9]), .A1 (
             AdderResult[9]), .S0 (nx225)) ;
    mux21_ni ix79 (.Y (AdderBoothResult[9]), .A0 (BoothP[10]), .A1 (
             AdderResult[10]), .S0 (nx225)) ;
    mux21_ni ix87 (.Y (AdderBoothResult[10]), .A0 (BoothP[11]), .A1 (
             AdderResult[11]), .S0 (nx225)) ;
    mux21_ni ix95 (.Y (AdderBoothResult[11]), .A0 (BoothP[12]), .A1 (
             AdderResult[12]), .S0 (nx225)) ;
    mux21_ni ix103 (.Y (AdderBoothResult[12]), .A0 (BoothP[13]), .A1 (
             AdderResult[13]), .S0 (nx225)) ;
    mux21_ni ix111 (.Y (AdderBoothResult[13]), .A0 (BoothP[14]), .A1 (
             AdderResult[14]), .S0 (nx225)) ;
    mux21_ni ix119 (.Y (AdderBoothResult[14]), .A0 (BoothP[15]), .A1 (
             AdderResult[15]), .S0 (nx227)) ;
    mux21_ni ix127 (.Y (AdderBoothResult[15]), .A0 (BoothP[16]), .A1 (
             AdderResult[16]), .S0 (nx227)) ;
    inv01 ix219 (.Y (nx220), .A (Operation)) ;
    inv02 ix221 (.Y (nx222), .A (nx220)) ;
    inv02 ix224 (.Y (nx225), .A (nx220)) ;
    inv02 ix226 (.Y (nx227), .A (nx220)) ;
    inv01 ix228 (.Y (nx229), .A (SelOperand)) ;
    inv02 ix230 (.Y (nx231), .A (nx229)) ;
    inv02 ix232 (.Y (nx233), .A (nx229)) ;
    inv02 ix234 (.Y (nx235), .A (nx229)) ;
    inv02 ix236 (.Y (nx237), .A (nx229)) ;
    inv02 ix238 (.Y (nx239), .A (nx229)) ;
endmodule


module booth_unit_17_unfolded1 ( CLK, RST, Start, Instr, 
                                 LoopingAndResultNotReady, Filter, Window, 
                                 AdderBoothResult, BoothXORCheck, BoothResult, 
                                 BoothAddingOperand, BoothP, LargeWindowShifted
                                  ) ;

    input CLK ;
    input RST ;
    input Start ;
    input Instr ;
    input LoopingAndResultNotReady ;
    input [7:0]Filter ;
    input [7:0]Window ;
    input [16:0]AdderBoothResult ;
    output BoothXORCheck ;
    output [7:0]BoothResult ;
    output [16:0]BoothAddingOperand ;
    output [16:0]BoothP ;
    output [16:0]LargeWindowShifted ;

    wire BoothP_0_rename, RegisterPEN, RegisterPDin_16, RegisterPDin_15, 
         RegisterPDin_14, RegisterPDin_13, RegisterPDin_12, RegisterPDin_11, 
         RegisterPDin_10, RegisterPDin_9, RegisterPDin_8, RegisterPDin_7, 
         RegisterPDin_6, RegisterPDin_5, RegisterPDin_4, RegisterPDin_3, 
         RegisterPDin_2, RegisterPDin_1, RegisterPDin_0, RegisterSDout_10, nx12, 
         nx20, RegisterADout_10, RegisterSDout_11, nx52, nx60, RegisterADout_11, 
         RegisterSDout_12, nx92, nx100, RegisterADout_12, RegisterSDout_13, 
         nx132, nx140, RegisterADout_13, RegisterSDout_14, nx172, nx180, 
         RegisterADout_14, RegisterSDout_15, nx212, nx220, RegisterADout_15, 
         RegisterSDout_16, nx246, RegisterADout_16, nx69, nx79, nx89, nx99, 
         nx109, nx119, nx129, nx139, nx149, nx159, nx169, nx179, nx189, nx199, 
         nx209, nx224, nx226, nx235, nx249, nx261, nx273, nx286, nx299, nx315, 
         nx324, nx326, nx328;
    wire [14:0] \$dummy ;




    assign BoothResult[7] = LargeWindowShifted[16] ;
    assign BoothResult[6] = LargeWindowShifted[16] ;
    assign BoothResult[5] = LargeWindowShifted[16] ;
    assign BoothResult[4] = LargeWindowShifted[16] ;
    assign BoothResult[3] = LargeWindowShifted[16] ;
    assign BoothResult[2] = LargeWindowShifted[16] ;
    assign BoothResult[1] = LargeWindowShifted[16] ;
    assign BoothResult[0] = LargeWindowShifted[16] ;
    assign BoothAddingOperand[8] = LargeWindowShifted[16] ;
    assign BoothAddingOperand[7] = LargeWindowShifted[16] ;
    assign BoothAddingOperand[6] = LargeWindowShifted[16] ;
    assign BoothAddingOperand[5] = LargeWindowShifted[16] ;
    assign BoothAddingOperand[4] = LargeWindowShifted[16] ;
    assign BoothAddingOperand[3] = LargeWindowShifted[16] ;
    assign BoothAddingOperand[2] = LargeWindowShifted[16] ;
    assign BoothAddingOperand[1] = LargeWindowShifted[16] ;
    assign BoothAddingOperand[0] = LargeWindowShifted[16] ;
    assign BoothP[0] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[15] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[14] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[13] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[12] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[11] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[10] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[9] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[8] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[7] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[6] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[5] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[4] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[3] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[2] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[1] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[0] = LargeWindowShifted[16] ;
    register_edge_17 REGISTER_P (.CLK (CLK), .RST (RST), .EN (RegisterPEN), .Din (
                     {RegisterPDin_16,RegisterPDin_15,RegisterPDin_14,
                     RegisterPDin_13,RegisterPDin_12,RegisterPDin_11,
                     RegisterPDin_10,RegisterPDin_9,RegisterPDin_8,
                     RegisterPDin_7,RegisterPDin_6,RegisterPDin_5,RegisterPDin_4
                     ,RegisterPDin_3,RegisterPDin_2,RegisterPDin_1,
                     RegisterPDin_0}), .Dout ({BoothP[16],BoothP[15],BoothP[14],
                     BoothP[13],BoothP[12],BoothP[11],BoothP[10],BoothP[9],
                     BoothP[8],BoothP[7],BoothP[6],BoothP[5],BoothP[4],BoothP[3]
                     ,BoothP[2],BoothP[1],BoothP_0_rename})) ;
    mux_4x1_17 P_INPUT_DATA_MUX (.A ({LargeWindowShifted[16],
               AdderBoothResult[15],AdderBoothResult[14],AdderBoothResult[13],
               AdderBoothResult[12],AdderBoothResult[11],AdderBoothResult[10],
               AdderBoothResult[9],AdderBoothResult[8],AdderBoothResult[7],
               AdderBoothResult[6],AdderBoothResult[5],AdderBoothResult[4],
               AdderBoothResult[3],AdderBoothResult[2],AdderBoothResult[1],
               AdderBoothResult[0]}), .B ({LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16]}), .C ({
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],Window[7],Window[6]
               ,Window[5],Window[4],Window[3],Window[2],Window[1],Window[0],
               LargeWindowShifted[16]}), .D ({LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16]}), .S ({Start,Instr
               }), .Dout ({RegisterPDin_16,RegisterPDin_15,RegisterPDin_14,
               RegisterPDin_13,RegisterPDin_12,RegisterPDin_11,RegisterPDin_10,
               RegisterPDin_9,RegisterPDin_8,RegisterPDin_7,RegisterPDin_6,
               RegisterPDin_5,RegisterPDin_4,RegisterPDin_3,RegisterPDin_2,
               RegisterPDin_1,RegisterPDin_0})) ;
    fake_gnd ix43 (.Y (LargeWindowShifted[16])) ;
    dff REGISTER_A_reg_Dout_9 (.Q (BoothAddingOperand[9]), .QB (\$dummy [0]), .D (
        nx209), .CLK (CLK)) ;
    ao32 ix210 (.Y (nx209), .A0 (nx324), .A1 (Filter[0]), .A2 (Start), .B0 (
         BoothAddingOperand[9]), .B1 (nx326)) ;
    inv01 ix225 (.Y (nx224), .A (RST)) ;
    nor02_2x ix227 (.Y (nx226), .A0 (Start), .A1 (RST)) ;
    or02 ix287 (.Y (RegisterPEN), .A0 (Start), .A1 (LoopingAndResultNotReady)) ;
    dff REGISTER_S_reg_Dout_10 (.Q (RegisterSDout_10), .QB (\$dummy [1]), .D (
        nx69), .CLK (CLK)) ;
    mux21_ni ix70 (.Y (nx69), .A0 (nx20), .A1 (RegisterSDout_10), .S0 (nx326)) ;
    aoi21 ix21 (.Y (nx20), .A0 (Filter[1]), .A1 (Filter[0]), .B0 (nx235)) ;
    or02 ix236 (.Y (nx235), .A0 (RST), .A1 (nx12)) ;
    nor02_2x ix13 (.Y (nx12), .A0 (Filter[0]), .A1 (Filter[1])) ;
    dff REGISTER_A_reg_Dout_10 (.Q (RegisterADout_10), .QB (\$dummy [2]), .D (
        nx79), .CLK (CLK)) ;
    ao32 ix80 (.Y (nx79), .A0 (nx324), .A1 (Filter[1]), .A2 (Start), .B0 (
         RegisterADout_10), .B1 (nx326)) ;
    dff REGISTER_S_reg_Dout_11 (.Q (RegisterSDout_11), .QB (\$dummy [3]), .D (
        nx89), .CLK (CLK)) ;
    mux21_ni ix90 (.Y (nx89), .A0 (nx60), .A1 (RegisterSDout_11), .S0 (nx326)) ;
    nor03_2x ix61 (.Y (nx60), .A0 (nx249), .A1 (RST), .A2 (nx52)) ;
    nor02ii ix250 (.Y (nx249), .A0 (nx12), .A1 (Filter[2])) ;
    nor03_2x ix53 (.Y (nx52), .A0 (Filter[2]), .A1 (Filter[0]), .A2 (Filter[1])
             ) ;
    dff REGISTER_A_reg_Dout_11 (.Q (RegisterADout_11), .QB (\$dummy [4]), .D (
        nx99), .CLK (CLK)) ;
    ao32 ix100 (.Y (nx99), .A0 (nx324), .A1 (Filter[2]), .A2 (Start), .B0 (
         RegisterADout_11), .B1 (nx326)) ;
    dff REGISTER_S_reg_Dout_12 (.Q (RegisterSDout_12), .QB (\$dummy [5]), .D (
        nx109), .CLK (CLK)) ;
    mux21_ni ix110 (.Y (nx109), .A0 (nx100), .A1 (RegisterSDout_12), .S0 (nx326)
             ) ;
    nor03_2x ix101 (.Y (nx100), .A0 (nx261), .A1 (RST), .A2 (nx92)) ;
    nor02ii ix262 (.Y (nx261), .A0 (nx52), .A1 (Filter[3])) ;
    nor04 ix93 (.Y (nx92), .A0 (Filter[3]), .A1 (Filter[2]), .A2 (Filter[0]), .A3 (
          Filter[1])) ;
    dff REGISTER_A_reg_Dout_12 (.Q (RegisterADout_12), .QB (\$dummy [6]), .D (
        nx119), .CLK (CLK)) ;
    ao32 ix120 (.Y (nx119), .A0 (nx324), .A1 (Filter[3]), .A2 (Start), .B0 (
         RegisterADout_12), .B1 (nx326)) ;
    dff REGISTER_S_reg_Dout_13 (.Q (RegisterSDout_13), .QB (\$dummy [7]), .D (
        nx129), .CLK (CLK)) ;
    mux21_ni ix130 (.Y (nx129), .A0 (nx140), .A1 (RegisterSDout_13), .S0 (nx328)
             ) ;
    nor03_2x ix141 (.Y (nx140), .A0 (nx273), .A1 (RST), .A2 (nx132)) ;
    nor02ii ix274 (.Y (nx273), .A0 (nx92), .A1 (Filter[4])) ;
    nor02ii ix133 (.Y (nx132), .A0 (Filter[4]), .A1 (nx92)) ;
    dff REGISTER_A_reg_Dout_13 (.Q (RegisterADout_13), .QB (\$dummy [8]), .D (
        nx139), .CLK (CLK)) ;
    ao32 ix140 (.Y (nx139), .A0 (nx324), .A1 (Filter[4]), .A2 (Start), .B0 (
         RegisterADout_13), .B1 (nx328)) ;
    dff REGISTER_S_reg_Dout_14 (.Q (RegisterSDout_14), .QB (\$dummy [9]), .D (
        nx149), .CLK (CLK)) ;
    mux21_ni ix150 (.Y (nx149), .A0 (nx180), .A1 (RegisterSDout_14), .S0 (nx328)
             ) ;
    nor03_2x ix181 (.Y (nx180), .A0 (nx286), .A1 (RST), .A2 (nx172)) ;
    nor02ii ix288 (.Y (nx286), .A0 (nx132), .A1 (Filter[5])) ;
    nor02ii ix173 (.Y (nx172), .A0 (Filter[5]), .A1 (nx132)) ;
    dff REGISTER_A_reg_Dout_14 (.Q (RegisterADout_14), .QB (\$dummy [10]), .D (
        nx159), .CLK (CLK)) ;
    ao32 ix160 (.Y (nx159), .A0 (nx324), .A1 (Filter[5]), .A2 (Start), .B0 (
         RegisterADout_14), .B1 (nx328)) ;
    dff REGISTER_S_reg_Dout_15 (.Q (RegisterSDout_15), .QB (\$dummy [11]), .D (
        nx169), .CLK (CLK)) ;
    mux21_ni ix170 (.Y (nx169), .A0 (nx220), .A1 (RegisterSDout_15), .S0 (nx328)
             ) ;
    nor03_2x ix221 (.Y (nx220), .A0 (nx299), .A1 (RST), .A2 (nx212)) ;
    nor02ii ix300 (.Y (nx299), .A0 (nx172), .A1 (Filter[6])) ;
    nor02ii ix213 (.Y (nx212), .A0 (Filter[6]), .A1 (nx172)) ;
    dff REGISTER_A_reg_Dout_15 (.Q (RegisterADout_15), .QB (\$dummy [12]), .D (
        nx179), .CLK (CLK)) ;
    ao32 ix180 (.Y (nx179), .A0 (nx324), .A1 (Filter[6]), .A2 (Start), .B0 (
         RegisterADout_15), .B1 (nx328)) ;
    dff REGISTER_S_reg_Dout_16 (.Q (RegisterSDout_16), .QB (\$dummy [13]), .D (
        nx189), .CLK (CLK)) ;
    ao32 ix190 (.Y (nx189), .A0 (nx224), .A1 (nx246), .A2 (Start), .B0 (
         RegisterSDout_16), .B1 (nx328)) ;
    xnor2 ix247 (.Y (nx246), .A0 (Filter[7]), .A1 (nx212)) ;
    dff REGISTER_A_reg_Dout_16 (.Q (RegisterADout_16), .QB (\$dummy [14]), .D (
        nx199), .CLK (CLK)) ;
    ao32 ix200 (.Y (nx199), .A0 (nx224), .A1 (Filter[7]), .A2 (Start), .B0 (
         RegisterADout_16), .B1 (nx226)) ;
    inv02 ix316 (.Y (nx315), .A (BoothP_0_rename)) ;
    inv01 ix323 (.Y (nx324), .A (RST)) ;
    nor02_2x ix325 (.Y (nx326), .A0 (Start), .A1 (RST)) ;
    nor02_2x ix327 (.Y (nx328), .A0 (Start), .A1 (RST)) ;
    mux21_ni ix46 (.Y (BoothAddingOperand[10]), .A0 (RegisterADout_10), .A1 (
             RegisterSDout_10), .S0 (nx315)) ;
    mux21_ni ix85 (.Y (BoothAddingOperand[11]), .A0 (RegisterADout_11), .A1 (
             RegisterSDout_11), .S0 (nx315)) ;
    mux21_ni ix125 (.Y (BoothAddingOperand[12]), .A0 (RegisterADout_12), .A1 (
             RegisterSDout_12), .S0 (nx315)) ;
    mux21_ni ix165 (.Y (BoothAddingOperand[13]), .A0 (RegisterADout_13), .A1 (
             RegisterSDout_13), .S0 (nx315)) ;
    mux21_ni ix205 (.Y (BoothAddingOperand[14]), .A0 (RegisterADout_14), .A1 (
             RegisterSDout_14), .S0 (nx315)) ;
    mux21_ni ix245 (.Y (BoothAddingOperand[15]), .A0 (RegisterADout_15), .A1 (
             RegisterSDout_15), .S0 (nx315)) ;
    mux21_ni ix275 (.Y (BoothAddingOperand[16]), .A0 (RegisterADout_16), .A1 (
             RegisterSDout_16), .S0 (nx315)) ;
    xor2 ix289 (.Y (BoothXORCheck), .A0 (BoothP[1]), .A1 (BoothP_0_rename)) ;
endmodule


module booth_adder_17_unfolded3 ( AdderFirstOperand, AdderSecondOperand, 
                                  BoothOperand, BoothP, SelOperand, Operation, 
                                  AdderResult, AdderBoothResult ) ;

    input [16:0]AdderFirstOperand ;
    input [16:0]AdderSecondOperand ;
    input [16:0]BoothOperand ;
    input [16:0]BoothP ;
    input SelOperand ;
    input Operation ;
    output [16:0]AdderResult ;
    output [16:0]AdderBoothResult ;

    wire AdderResult_16_rename, AdderResult_15_rename, AdderResult_14_rename, 
         AdderResult_13_rename, AdderResult_12_rename, AdderResult_11_rename, 
         AdderResult_10_rename, AdderResult_9_rename, FirstOperand_16, 
         FirstOperand_15, FirstOperand_14, FirstOperand_13, FirstOperand_12, 
         FirstOperand_11, FirstOperand_10, FirstOperand_9, SecondOperand_16, 
         SecondOperand_15, SecondOperand_14, SecondOperand_13, SecondOperand_12, 
         SecondOperand_11, SecondOperand_10, SecondOperand_9, SecondOperand_8, 
         SecondOperand_7, SecondOperand_6, SecondOperand_5, SecondOperand_4, 
         nx143, nx153, nx155, nx158, nx161, nx164, nx167, nx182, nx184, nx186, 
         nx188, nx190, nx192, nx194;
    wire [9:0] \$dummy ;




    assign AdderResult[16] = AdderBoothResult[16] ;
    assign AdderResult[15] = AdderBoothResult[16] ;
    assign AdderResult[14] = AdderBoothResult[16] ;
    assign AdderResult[13] = AdderBoothResult[16] ;
    assign AdderResult[12] = AdderBoothResult[16] ;
    assign AdderResult[11] = AdderBoothResult[16] ;
    assign AdderResult[10] = AdderBoothResult[16] ;
    assign AdderResult[9] = AdderBoothResult[16] ;
    assign AdderResult[8] = AdderBoothResult[16] ;
    assign AdderResult[7] = AdderBoothResult[16] ;
    assign AdderResult[6] = AdderBoothResult[16] ;
    assign AdderResult[5] = AdderBoothResult[16] ;
    assign AdderResult[4] = AdderBoothResult[16] ;
    assign AdderResult[3] = AdderBoothResult[16] ;
    assign AdderResult[2] = AdderBoothResult[16] ;
    assign AdderResult[1] = AdderBoothResult[16] ;
    assign AdderResult[0] = AdderBoothResult[16] ;
    adder_17_unfolded1 ADDER (.A ({FirstOperand_16,FirstOperand_15,
                       FirstOperand_14,FirstOperand_13,FirstOperand_12,
                       FirstOperand_11,FirstOperand_10,FirstOperand_9,
                       AdderBoothResult[16],AdderBoothResult[16],
                       AdderBoothResult[16],AdderBoothResult[16],
                       AdderBoothResult[16],AdderBoothResult[16],
                       AdderBoothResult[16],AdderBoothResult[16],
                       AdderBoothResult[16]}), .B ({SecondOperand_16,
                       SecondOperand_15,SecondOperand_14,SecondOperand_13,
                       SecondOperand_12,SecondOperand_11,SecondOperand_10,
                       SecondOperand_9,SecondOperand_8,SecondOperand_7,
                       SecondOperand_6,SecondOperand_5,SecondOperand_4,
                       AdderBoothResult[16],AdderBoothResult[16],
                       AdderBoothResult[16],AdderBoothResult[16]}), .Cin (
                       AdderBoothResult[16]), .Sum ({AdderResult_16_rename,
                       AdderResult_15_rename,AdderResult_14_rename,
                       AdderResult_13_rename,AdderResult_12_rename,
                       AdderResult_11_rename,AdderResult_10_rename,
                       AdderResult_9_rename,\$dummy [0],\$dummy [1],\$dummy [2],
                       \$dummy [3],\$dummy [4],\$dummy [5],\$dummy [6],
                       \$dummy [7],\$dummy [8]}), .Cout (\$dummy [9])) ;
    fake_gnd ix59 (.Y (AdderBoothResult[16])) ;
    and02 ix15 (.Y (SecondOperand_4), .A0 (BoothP[4]), .A1 (nx186)) ;
    and02 ix25 (.Y (SecondOperand_5), .A0 (BoothP[5]), .A1 (nx186)) ;
    and02 ix35 (.Y (SecondOperand_6), .A0 (BoothP[6]), .A1 (nx186)) ;
    and02 ix45 (.Y (SecondOperand_7), .A0 (BoothP[7]), .A1 (nx186)) ;
    and02 ix55 (.Y (SecondOperand_8), .A0 (BoothP[8]), .A1 (nx186)) ;
    and02 ix125 (.Y (SecondOperand_9), .A0 (BoothP[9]), .A1 (nx186)) ;
    and02 ix127 (.Y (SecondOperand_10), .A0 (BoothP[10]), .A1 (nx186)) ;
    and02 ix129 (.Y (SecondOperand_11), .A0 (BoothP[11]), .A1 (nx188)) ;
    and02 ix131 (.Y (SecondOperand_12), .A0 (BoothP[12]), .A1 (nx188)) ;
    and02 ix133 (.Y (SecondOperand_13), .A0 (BoothP[13]), .A1 (nx188)) ;
    and02 ix135 (.Y (SecondOperand_14), .A0 (BoothP[14]), .A1 (nx188)) ;
    and02 ix137 (.Y (SecondOperand_15), .A0 (BoothP[15]), .A1 (nx188)) ;
    and02 ix139 (.Y (SecondOperand_16), .A0 (BoothP[16]), .A1 (nx188)) ;
    and02 ix141 (.Y (FirstOperand_9), .A0 (BoothOperand[9]), .A1 (nx188)) ;
    and02 ix143 (.Y (FirstOperand_10), .A0 (BoothOperand[10]), .A1 (nx190)) ;
    and02 ix145 (.Y (FirstOperand_11), .A0 (BoothOperand[11]), .A1 (nx190)) ;
    and02 ix147 (.Y (FirstOperand_12), .A0 (BoothOperand[12]), .A1 (nx190)) ;
    and02 ix149 (.Y (FirstOperand_13), .A0 (BoothOperand[13]), .A1 (nx190)) ;
    and02 ix151 (.Y (FirstOperand_14), .A0 (BoothOperand[14]), .A1 (nx190)) ;
    and02 ix153 (.Y (FirstOperand_15), .A0 (BoothOperand[15]), .A1 (nx190)) ;
    and02 ix155 (.Y (FirstOperand_16), .A0 (nx190), .A1 (BoothOperand[16])) ;
    nor02ii ix5 (.Y (AdderBoothResult[0]), .A0 (nx143), .A1 (BoothP[1])) ;
    nor02ii ix7 (.Y (AdderBoothResult[1]), .A0 (nx143), .A1 (BoothP[2])) ;
    nor02ii ix9 (.Y (AdderBoothResult[2]), .A0 (nx143), .A1 (BoothP[3])) ;
    aoi21 ix19 (.Y (AdderBoothResult[3]), .A0 (nx182), .A1 (nx194), .B0 (nx155)
          ) ;
    inv01 ix154 (.Y (nx153), .A (SelOperand)) ;
    inv01 ix156 (.Y (nx155), .A (BoothP[4])) ;
    aoi21 ix29 (.Y (AdderBoothResult[4]), .A0 (nx182), .A1 (nx194), .B0 (nx158)
          ) ;
    inv01 ix159 (.Y (nx158), .A (BoothP[5])) ;
    aoi21 ix39 (.Y (AdderBoothResult[5]), .A0 (nx182), .A1 (nx194), .B0 (nx161)
          ) ;
    inv01 ix162 (.Y (nx161), .A (BoothP[6])) ;
    aoi21 ix49 (.Y (AdderBoothResult[6]), .A0 (nx182), .A1 (nx194), .B0 (nx164)
          ) ;
    inv01 ix165 (.Y (nx164), .A (BoothP[7])) ;
    aoi21 ix61 (.Y (AdderBoothResult[7]), .A0 (nx182), .A1 (nx194), .B0 (nx167)
          ) ;
    inv01 ix168 (.Y (nx167), .A (BoothP[8])) ;
    mux21_ni ix67 (.Y (AdderBoothResult[8]), .A0 (BoothP[9]), .A1 (
             AdderResult_9_rename), .S0 (nx182)) ;
    mux21_ni ix75 (.Y (AdderBoothResult[9]), .A0 (BoothP[10]), .A1 (
             AdderResult_10_rename), .S0 (nx182)) ;
    mux21_ni ix83 (.Y (AdderBoothResult[10]), .A0 (BoothP[11]), .A1 (
             AdderResult_11_rename), .S0 (nx184)) ;
    mux21_ni ix91 (.Y (AdderBoothResult[11]), .A0 (BoothP[12]), .A1 (
             AdderResult_12_rename), .S0 (nx184)) ;
    mux21_ni ix99 (.Y (AdderBoothResult[12]), .A0 (BoothP[13]), .A1 (
             AdderResult_13_rename), .S0 (nx184)) ;
    mux21_ni ix107 (.Y (AdderBoothResult[13]), .A0 (BoothP[14]), .A1 (
             AdderResult_14_rename), .S0 (nx184)) ;
    mux21_ni ix115 (.Y (AdderBoothResult[14]), .A0 (BoothP[15]), .A1 (
             AdderResult_15_rename), .S0 (nx184)) ;
    mux21_ni ix123 (.Y (AdderBoothResult[15]), .A0 (BoothP[16]), .A1 (
             AdderResult_16_rename), .S0 (nx184)) ;
    nor02ii ix144 (.Y (nx143), .A0 (nx192), .A1 (nx184)) ;
    buf02 ix181 (.Y (nx182), .A (Operation)) ;
    buf02 ix183 (.Y (nx184), .A (Operation)) ;
    inv02 ix185 (.Y (nx186), .A (nx194)) ;
    inv02 ix187 (.Y (nx188), .A (nx153)) ;
    inv02 ix189 (.Y (nx190), .A (nx153)) ;
    inv02 ix191 (.Y (nx192), .A (nx153)) ;
    inv01 ix193 (.Y (nx194), .A (SelOperand)) ;
endmodule


module adder_17_unfolded1 ( A, B, Cin, Sum, Cout ) ;

    input [16:0]A ;
    input [16:0]B ;
    input Cin ;
    output [16:0]Sum ;
    output Cout ;

    wire nx2, nx16, nx18, nx32, nx34, nx48, nx93, nx95, nx98, nx101, nx105, 
         nx107, nx110, nx113, nx117, nx119, nx122, nx125, nx129, nx131;



    assign Sum[8] = B[8] ;
    assign Sum[7] = B[7] ;
    assign Sum[6] = B[6] ;
    assign Sum[5] = B[5] ;
    assign Sum[4] = B[4] ;
    assign Sum[3] = Cout ;
    assign Sum[2] = Cout ;
    assign Sum[1] = Cout ;
    assign Sum[0] = Cout ;
    fake_gnd ix68 (.Y (Cout)) ;
    xor2 ix71 (.Y (Sum[9]), .A0 (B[9]), .A1 (A[9])) ;
    xor2 ix65 (.Y (Sum[10]), .A0 (nx93), .A1 (nx95)) ;
    nand02 ix94 (.Y (nx93), .A0 (B[9]), .A1 (A[9])) ;
    xnor2 ix96 (.Y (nx95), .A0 (A[10]), .A1 (B[10])) ;
    xor2 ix63 (.Y (Sum[11]), .A0 (nx98), .A1 (nx101)) ;
    aoi32 ix99 (.Y (nx98), .A0 (B[9]), .A1 (A[9]), .A2 (nx2), .B0 (B[10]), .B1 (
          A[10])) ;
    xnor2 ix102 (.Y (nx101), .A0 (A[11]), .A1 (B[11])) ;
    xnor2 ix61 (.Y (Sum[12]), .A0 (nx16), .A1 (nx107)) ;
    oai21 ix17 (.Y (nx16), .A0 (nx98), .A1 (nx101), .B0 (nx105)) ;
    nand02 ix106 (.Y (nx105), .A0 (B[11]), .A1 (A[11])) ;
    xnor2 ix108 (.Y (nx107), .A0 (A[12]), .A1 (B[12])) ;
    xor2 ix59 (.Y (Sum[13]), .A0 (nx110), .A1 (nx113)) ;
    aoi22 ix111 (.Y (nx110), .A0 (B[12]), .A1 (A[12]), .B0 (nx16), .B1 (nx18)) ;
    xnor2 ix114 (.Y (nx113), .A0 (A[13]), .A1 (B[13])) ;
    xnor2 ix57 (.Y (Sum[14]), .A0 (nx32), .A1 (nx119)) ;
    oai21 ix33 (.Y (nx32), .A0 (nx110), .A1 (nx113), .B0 (nx117)) ;
    nand02 ix118 (.Y (nx117), .A0 (B[13]), .A1 (A[13])) ;
    xnor2 ix120 (.Y (nx119), .A0 (A[14]), .A1 (B[14])) ;
    xor2 ix55 (.Y (Sum[15]), .A0 (nx122), .A1 (nx125)) ;
    aoi22 ix123 (.Y (nx122), .A0 (B[14]), .A1 (A[14]), .B0 (nx32), .B1 (nx34)) ;
    xnor2 ix126 (.Y (nx125), .A0 (A[15]), .A1 (B[15])) ;
    xnor2 ix53 (.Y (Sum[16]), .A0 (nx48), .A1 (nx131)) ;
    oai21 ix49 (.Y (nx48), .A0 (nx122), .A1 (nx125), .B0 (nx129)) ;
    nand02 ix130 (.Y (nx129), .A0 (B[15]), .A1 (A[15])) ;
    xnor2 ix132 (.Y (nx131), .A0 (A[16]), .A1 (B[16])) ;
    inv01 ix35 (.Y (nx34), .A (nx119)) ;
    inv01 ix19 (.Y (nx18), .A (nx107)) ;
    inv01 ix3 (.Y (nx2), .A (nx95)) ;
endmodule


module booth_unit_17 ( CLK, RST, Start, Instr, LoopingAndResultNotReady, Filter, 
                       Window, AdderBoothResult, BoothXORCheck, BoothResult, 
                       BoothAddingOperand, BoothP, LargeWindowShifted ) ;

    input CLK ;
    input RST ;
    input Start ;
    input Instr ;
    input LoopingAndResultNotReady ;
    input [7:0]Filter ;
    input [7:0]Window ;
    input [16:0]AdderBoothResult ;
    output BoothXORCheck ;
    output [7:0]BoothResult ;
    output [16:0]BoothAddingOperand ;
    output [16:0]BoothP ;
    output [16:0]LargeWindowShifted ;

    wire RegisterPEN, RegisterPDin_16, RegisterPDin_15, RegisterPDin_14, 
         RegisterPDin_13, RegisterPDin_12, RegisterPDin_11, RegisterPDin_10, 
         RegisterPDin_9, RegisterPDin_8, RegisterPDin_7, RegisterPDin_6, 
         RegisterPDin_5, RegisterPDin_4, RegisterPDin_3, RegisterPDin_2, 
         RegisterPDin_1, RegisterPDin_0, RegisterSDout_10, nx12, nx20, 
         RegisterADout_10, RegisterSDout_11, nx52, nx60, RegisterADout_11, 
         RegisterSDout_12, nx92, nx100, RegisterADout_12, RegisterSDout_13, 
         nx132, nx140, RegisterADout_13, RegisterSDout_14, nx172, nx180, 
         RegisterADout_14, RegisterSDout_15, nx212, nx220, RegisterADout_15, 
         RegisterSDout_16, nx246, RegisterADout_16, nx69, nx79, nx89, nx99, 
         nx109, nx119, nx129, nx139, nx149, nx159, nx169, nx179, nx189, nx199, 
         nx209, nx224, nx226, nx235, nx249, nx261, nx273, nx286, nx299, nx320, 
         nx322, nx324, nx326, nx328;
    wire [14:0] \$dummy ;




    assign BoothResult[7] = LargeWindowShifted[16] ;
    assign BoothResult[6] = LargeWindowShifted[16] ;
    assign BoothResult[5] = LargeWindowShifted[16] ;
    assign BoothResult[4] = LargeWindowShifted[16] ;
    assign BoothResult[3] = LargeWindowShifted[16] ;
    assign BoothResult[2] = LargeWindowShifted[16] ;
    assign BoothResult[1] = LargeWindowShifted[16] ;
    assign BoothResult[0] = LargeWindowShifted[16] ;
    assign BoothAddingOperand[8] = LargeWindowShifted[16] ;
    assign BoothAddingOperand[7] = LargeWindowShifted[16] ;
    assign BoothAddingOperand[6] = LargeWindowShifted[16] ;
    assign BoothAddingOperand[5] = LargeWindowShifted[16] ;
    assign BoothAddingOperand[4] = LargeWindowShifted[16] ;
    assign BoothAddingOperand[3] = LargeWindowShifted[16] ;
    assign BoothAddingOperand[2] = LargeWindowShifted[16] ;
    assign BoothAddingOperand[1] = LargeWindowShifted[16] ;
    assign BoothAddingOperand[0] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[15] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[14] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[13] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[12] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[11] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[10] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[9] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[8] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[7] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[6] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[5] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[4] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[3] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[2] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[1] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[0] = LargeWindowShifted[16] ;
    register_edge_17 REGISTER_P (.CLK (CLK), .RST (RST), .EN (RegisterPEN), .Din (
                     {RegisterPDin_16,RegisterPDin_15,RegisterPDin_14,
                     RegisterPDin_13,RegisterPDin_12,RegisterPDin_11,
                     RegisterPDin_10,RegisterPDin_9,RegisterPDin_8,
                     RegisterPDin_7,RegisterPDin_6,RegisterPDin_5,RegisterPDin_4
                     ,RegisterPDin_3,RegisterPDin_2,RegisterPDin_1,
                     RegisterPDin_0}), .Dout ({BoothP[16],BoothP[15],BoothP[14],
                     BoothP[13],BoothP[12],BoothP[11],BoothP[10],BoothP[9],
                     BoothP[8],BoothP[7],BoothP[6],BoothP[5],BoothP[4],BoothP[3]
                     ,BoothP[2],BoothP[1],BoothP[0]})) ;
    mux_4x1_17 P_INPUT_DATA_MUX (.A ({LargeWindowShifted[16],
               AdderBoothResult[15],AdderBoothResult[14],AdderBoothResult[13],
               AdderBoothResult[12],AdderBoothResult[11],AdderBoothResult[10],
               AdderBoothResult[9],AdderBoothResult[8],AdderBoothResult[7],
               AdderBoothResult[6],AdderBoothResult[5],AdderBoothResult[4],
               AdderBoothResult[3],AdderBoothResult[2],AdderBoothResult[1],
               AdderBoothResult[0]}), .B ({LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16]}), .C ({
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],Window[7],Window[6]
               ,Window[5],Window[4],Window[3],Window[2],Window[1],Window[0],
               LargeWindowShifted[16]}), .D ({LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16]}), .S ({Start,Instr
               }), .Dout ({RegisterPDin_16,RegisterPDin_15,RegisterPDin_14,
               RegisterPDin_13,RegisterPDin_12,RegisterPDin_11,RegisterPDin_10,
               RegisterPDin_9,RegisterPDin_8,RegisterPDin_7,RegisterPDin_6,
               RegisterPDin_5,RegisterPDin_4,RegisterPDin_3,RegisterPDin_2,
               RegisterPDin_1,RegisterPDin_0})) ;
    fake_gnd ix43 (.Y (LargeWindowShifted[16])) ;
    dff REGISTER_A_reg_Dout_9 (.Q (BoothAddingOperand[9]), .QB (\$dummy [0]), .D (
        nx209), .CLK (CLK)) ;
    ao32 ix210 (.Y (nx209), .A0 (nx324), .A1 (Filter[0]), .A2 (Start), .B0 (
         BoothAddingOperand[9]), .B1 (nx326)) ;
    inv01 ix225 (.Y (nx224), .A (RST)) ;
    nor02_2x ix227 (.Y (nx226), .A0 (Start), .A1 (RST)) ;
    or02 ix287 (.Y (RegisterPEN), .A0 (Start), .A1 (LoopingAndResultNotReady)) ;
    mux21_ni ix46 (.Y (BoothAddingOperand[10]), .A0 (RegisterSDout_10), .A1 (
             RegisterADout_10), .S0 (nx320)) ;
    dff REGISTER_S_reg_Dout_10 (.Q (RegisterSDout_10), .QB (\$dummy [1]), .D (
        nx69), .CLK (CLK)) ;
    mux21_ni ix70 (.Y (nx69), .A0 (nx20), .A1 (RegisterSDout_10), .S0 (nx326)) ;
    aoi21 ix21 (.Y (nx20), .A0 (Filter[1]), .A1 (Filter[0]), .B0 (nx235)) ;
    or02 ix236 (.Y (nx235), .A0 (RST), .A1 (nx12)) ;
    nor02_2x ix13 (.Y (nx12), .A0 (Filter[0]), .A1 (Filter[1])) ;
    dff REGISTER_A_reg_Dout_10 (.Q (RegisterADout_10), .QB (\$dummy [2]), .D (
        nx79), .CLK (CLK)) ;
    ao32 ix80 (.Y (nx79), .A0 (nx324), .A1 (Filter[1]), .A2 (Start), .B0 (
         RegisterADout_10), .B1 (nx326)) ;
    mux21_ni ix85 (.Y (BoothAddingOperand[11]), .A0 (RegisterSDout_11), .A1 (
             RegisterADout_11), .S0 (nx320)) ;
    dff REGISTER_S_reg_Dout_11 (.Q (RegisterSDout_11), .QB (\$dummy [3]), .D (
        nx89), .CLK (CLK)) ;
    mux21_ni ix90 (.Y (nx89), .A0 (nx60), .A1 (RegisterSDout_11), .S0 (nx326)) ;
    nor03_2x ix61 (.Y (nx60), .A0 (nx249), .A1 (RST), .A2 (nx52)) ;
    nor02ii ix250 (.Y (nx249), .A0 (nx12), .A1 (Filter[2])) ;
    nor03_2x ix53 (.Y (nx52), .A0 (Filter[2]), .A1 (Filter[0]), .A2 (Filter[1])
             ) ;
    dff REGISTER_A_reg_Dout_11 (.Q (RegisterADout_11), .QB (\$dummy [4]), .D (
        nx99), .CLK (CLK)) ;
    ao32 ix100 (.Y (nx99), .A0 (nx324), .A1 (Filter[2]), .A2 (Start), .B0 (
         RegisterADout_11), .B1 (nx326)) ;
    mux21_ni ix125 (.Y (BoothAddingOperand[12]), .A0 (RegisterSDout_12), .A1 (
             RegisterADout_12), .S0 (nx320)) ;
    dff REGISTER_S_reg_Dout_12 (.Q (RegisterSDout_12), .QB (\$dummy [5]), .D (
        nx109), .CLK (CLK)) ;
    mux21_ni ix110 (.Y (nx109), .A0 (nx100), .A1 (RegisterSDout_12), .S0 (nx326)
             ) ;
    nor03_2x ix101 (.Y (nx100), .A0 (nx261), .A1 (RST), .A2 (nx92)) ;
    nor02ii ix262 (.Y (nx261), .A0 (nx52), .A1 (Filter[3])) ;
    nor04 ix93 (.Y (nx92), .A0 (Filter[3]), .A1 (Filter[2]), .A2 (Filter[0]), .A3 (
          Filter[1])) ;
    dff REGISTER_A_reg_Dout_12 (.Q (RegisterADout_12), .QB (\$dummy [6]), .D (
        nx119), .CLK (CLK)) ;
    ao32 ix120 (.Y (nx119), .A0 (nx324), .A1 (Filter[3]), .A2 (Start), .B0 (
         RegisterADout_12), .B1 (nx326)) ;
    mux21_ni ix165 (.Y (BoothAddingOperand[13]), .A0 (RegisterSDout_13), .A1 (
             RegisterADout_13), .S0 (nx320)) ;
    dff REGISTER_S_reg_Dout_13 (.Q (RegisterSDout_13), .QB (\$dummy [7]), .D (
        nx129), .CLK (CLK)) ;
    mux21_ni ix130 (.Y (nx129), .A0 (nx140), .A1 (RegisterSDout_13), .S0 (nx328)
             ) ;
    nor03_2x ix141 (.Y (nx140), .A0 (nx273), .A1 (RST), .A2 (nx132)) ;
    nor02ii ix274 (.Y (nx273), .A0 (nx92), .A1 (Filter[4])) ;
    nor02ii ix133 (.Y (nx132), .A0 (Filter[4]), .A1 (nx92)) ;
    dff REGISTER_A_reg_Dout_13 (.Q (RegisterADout_13), .QB (\$dummy [8]), .D (
        nx139), .CLK (CLK)) ;
    ao32 ix140 (.Y (nx139), .A0 (nx324), .A1 (Filter[4]), .A2 (Start), .B0 (
         RegisterADout_13), .B1 (nx328)) ;
    mux21_ni ix205 (.Y (BoothAddingOperand[14]), .A0 (RegisterSDout_14), .A1 (
             RegisterADout_14), .S0 (nx320)) ;
    dff REGISTER_S_reg_Dout_14 (.Q (RegisterSDout_14), .QB (\$dummy [9]), .D (
        nx149), .CLK (CLK)) ;
    mux21_ni ix150 (.Y (nx149), .A0 (nx180), .A1 (RegisterSDout_14), .S0 (nx328)
             ) ;
    nor03_2x ix181 (.Y (nx180), .A0 (nx286), .A1 (RST), .A2 (nx172)) ;
    nor02ii ix288 (.Y (nx286), .A0 (nx132), .A1 (Filter[5])) ;
    nor02ii ix173 (.Y (nx172), .A0 (Filter[5]), .A1 (nx132)) ;
    dff REGISTER_A_reg_Dout_14 (.Q (RegisterADout_14), .QB (\$dummy [10]), .D (
        nx159), .CLK (CLK)) ;
    ao32 ix160 (.Y (nx159), .A0 (nx324), .A1 (Filter[5]), .A2 (Start), .B0 (
         RegisterADout_14), .B1 (nx328)) ;
    mux21_ni ix245 (.Y (BoothAddingOperand[15]), .A0 (RegisterSDout_15), .A1 (
             RegisterADout_15), .S0 (nx320)) ;
    dff REGISTER_S_reg_Dout_15 (.Q (RegisterSDout_15), .QB (\$dummy [11]), .D (
        nx169), .CLK (CLK)) ;
    mux21_ni ix170 (.Y (nx169), .A0 (nx220), .A1 (RegisterSDout_15), .S0 (nx328)
             ) ;
    nor03_2x ix221 (.Y (nx220), .A0 (nx299), .A1 (RST), .A2 (nx212)) ;
    nor02ii ix300 (.Y (nx299), .A0 (nx172), .A1 (Filter[6])) ;
    nor02ii ix213 (.Y (nx212), .A0 (Filter[6]), .A1 (nx172)) ;
    dff REGISTER_A_reg_Dout_15 (.Q (RegisterADout_15), .QB (\$dummy [12]), .D (
        nx179), .CLK (CLK)) ;
    ao32 ix180 (.Y (nx179), .A0 (nx324), .A1 (Filter[6]), .A2 (Start), .B0 (
         RegisterADout_15), .B1 (nx328)) ;
    mux21_ni ix275 (.Y (BoothAddingOperand[16]), .A0 (RegisterSDout_16), .A1 (
             RegisterADout_16), .S0 (nx320)) ;
    dff REGISTER_S_reg_Dout_16 (.Q (RegisterSDout_16), .QB (\$dummy [13]), .D (
        nx189), .CLK (CLK)) ;
    ao32 ix190 (.Y (nx189), .A0 (nx224), .A1 (nx246), .A2 (Start), .B0 (
         RegisterSDout_16), .B1 (nx328)) ;
    xnor2 ix247 (.Y (nx246), .A0 (Filter[7]), .A1 (nx212)) ;
    dff REGISTER_A_reg_Dout_16 (.Q (RegisterADout_16), .QB (\$dummy [14]), .D (
        nx199), .CLK (CLK)) ;
    ao32 ix200 (.Y (nx199), .A0 (nx224), .A1 (Filter[7]), .A2 (Start), .B0 (
         RegisterADout_16), .B1 (nx226)) ;
    xor2 ix289 (.Y (BoothXORCheck), .A0 (BoothP[1]), .A1 (nx322)) ;
    buf02 ix319 (.Y (nx320), .A (BoothP[0])) ;
    buf02 ix321 (.Y (nx322), .A (BoothP[0])) ;
    inv01 ix323 (.Y (nx324), .A (RST)) ;
    nor02_2x ix325 (.Y (nx326), .A0 (Start), .A1 (RST)) ;
    nor02_2x ix327 (.Y (nx328), .A0 (Start), .A1 (RST)) ;
endmodule


module mux_4x1_17 ( A, B, C, D, S, Dout ) ;

    input [16:0]A ;
    input [16:0]B ;
    input [16:0]C ;
    input [16:0]D ;
    input [1:0]S ;
    output [16:0]Dout ;

    wire nx28, nx46, nx131, nx136, nx139, nx142, nx145, nx148, nx151, nx166, 
         nx168, nx170, nx172, nx178, nx180;



    fake_gnd ix85 (.Y (Dout[16])) ;
    ao22 ix37 (.Y (Dout[0]), .A0 (A[0]), .A1 (nx170), .B0 (C[1]), .B1 (nx166)) ;
    and02 ix29 (.Y (nx28), .A0 (S[0]), .A1 (S[1])) ;
    inv01 ix53 (.Y (Dout[1]), .A (nx131)) ;
    aoi222 ix132 (.Y (nx131), .A0 (A[1]), .A1 (nx170), .B0 (C[1]), .B1 (nx178), 
           .C0 (C[2]), .C1 (nx166)) ;
    inv01 ix65 (.Y (Dout[2]), .A (nx136)) ;
    aoi222 ix137 (.Y (nx136), .A0 (A[2]), .A1 (nx170), .B0 (C[2]), .B1 (nx178), 
           .C0 (C[3]), .C1 (nx166)) ;
    inv01 ix77 (.Y (Dout[3]), .A (nx139)) ;
    aoi222 ix140 (.Y (nx139), .A0 (A[3]), .A1 (nx170), .B0 (C[3]), .B1 (nx178), 
           .C0 (C[4]), .C1 (nx166)) ;
    inv01 ix89 (.Y (Dout[4]), .A (nx142)) ;
    aoi222 ix143 (.Y (nx142), .A0 (A[4]), .A1 (nx170), .B0 (C[4]), .B1 (nx178), 
           .C0 (C[5]), .C1 (nx166)) ;
    inv01 ix101 (.Y (Dout[5]), .A (nx145)) ;
    aoi222 ix146 (.Y (nx145), .A0 (A[5]), .A1 (nx170), .B0 (C[5]), .B1 (nx178), 
           .C0 (C[6]), .C1 (nx166)) ;
    inv01 ix113 (.Y (Dout[6]), .A (nx148)) ;
    aoi222 ix149 (.Y (nx148), .A0 (A[6]), .A1 (nx172), .B0 (C[6]), .B1 (nx178), 
           .C0 (C[7]), .C1 (nx166)) ;
    inv01 ix125 (.Y (Dout[7]), .A (nx151)) ;
    aoi222 ix152 (.Y (nx151), .A0 (A[7]), .A1 (nx172), .B0 (C[7]), .B1 (nx178), 
           .C0 (C[8]), .C1 (nx168)) ;
    ao22 ix133 (.Y (Dout[8]), .A0 (nx172), .A1 (A[8]), .B0 (C[8]), .B1 (nx180)
         ) ;
    nor02ii ix3 (.Y (Dout[9]), .A0 (S[1]), .A1 (A[9])) ;
    nor02ii ix7 (.Y (Dout[10]), .A0 (S[1]), .A1 (A[10])) ;
    nor02ii ix11 (.Y (Dout[11]), .A0 (S[1]), .A1 (A[11])) ;
    nor02ii ix15 (.Y (Dout[12]), .A0 (S[1]), .A1 (A[12])) ;
    nor02ii ix19 (.Y (Dout[13]), .A0 (S[1]), .A1 (A[13])) ;
    nor02ii ix23 (.Y (Dout[14]), .A0 (S[1]), .A1 (A[14])) ;
    nor02ii ix27 (.Y (Dout[15]), .A0 (S[1]), .A1 (A[15])) ;
    buf02 ix165 (.Y (nx166), .A (nx28)) ;
    buf02 ix167 (.Y (nx168), .A (nx28)) ;
    inv02 ix169 (.Y (nx170), .A (S[1])) ;
    inv02 ix171 (.Y (nx172), .A (S[1])) ;
    nor02ii ix47 (.Y (nx46), .A0 (S[0]), .A1 (S[1])) ;
    buf02 ix177 (.Y (nx178), .A (nx46)) ;
    buf02 ix179 (.Y (nx180), .A (nx46)) ;
endmodule


module register_edge_17 ( CLK, RST, EN, Din, Dout ) ;

    input CLK ;
    input RST ;
    input EN ;
    input [16:0]Din ;
    output [16:0]Dout ;

    wire nx402, nx412, nx422, nx432, nx442, nx452, nx462, nx472, nx482, nx492, 
         nx502, nx512, nx522, nx532, nx542, nx552, nx562, nx574, nx576, nx632, 
         nx634, nx636, nx638, nx644, nx646, nx648, nx650;
    wire [16:0] \$dummy ;




    dff reg_Dout_0 (.Q (Dout[0]), .QB (\$dummy [0]), .D (nx402), .CLK (CLK)) ;
    ao32 ix403 (.Y (nx402), .A0 (Din[0]), .A1 (nx632), .A2 (nx646), .B0 (Dout[0]
         ), .B1 (nx636)) ;
    inv01 ix575 (.Y (nx574), .A (RST)) ;
    nor02_2x ix577 (.Y (nx576), .A0 (RST), .A1 (nx646)) ;
    dff reg_Dout_1 (.Q (Dout[1]), .QB (\$dummy [1]), .D (nx412), .CLK (CLK)) ;
    ao32 ix413 (.Y (nx412), .A0 (Din[1]), .A1 (nx632), .A2 (nx646), .B0 (Dout[1]
         ), .B1 (nx636)) ;
    dff reg_Dout_2 (.Q (Dout[2]), .QB (\$dummy [2]), .D (nx422), .CLK (CLK)) ;
    ao32 ix423 (.Y (nx422), .A0 (Din[2]), .A1 (nx632), .A2 (nx646), .B0 (Dout[2]
         ), .B1 (nx636)) ;
    dff reg_Dout_3 (.Q (Dout[3]), .QB (\$dummy [3]), .D (nx432), .CLK (CLK)) ;
    ao32 ix433 (.Y (nx432), .A0 (Din[3]), .A1 (nx632), .A2 (nx646), .B0 (Dout[3]
         ), .B1 (nx636)) ;
    dff reg_Dout_4 (.Q (Dout[4]), .QB (\$dummy [4]), .D (nx442), .CLK (CLK)) ;
    ao32 ix443 (.Y (nx442), .A0 (Din[4]), .A1 (nx632), .A2 (nx646), .B0 (Dout[4]
         ), .B1 (nx636)) ;
    dff reg_Dout_5 (.Q (Dout[5]), .QB (\$dummy [5]), .D (nx452), .CLK (CLK)) ;
    ao32 ix453 (.Y (nx452), .A0 (Din[5]), .A1 (nx632), .A2 (nx646), .B0 (Dout[5]
         ), .B1 (nx636)) ;
    dff reg_Dout_6 (.Q (Dout[6]), .QB (\$dummy [6]), .D (nx462), .CLK (CLK)) ;
    ao32 ix463 (.Y (nx462), .A0 (Din[6]), .A1 (nx634), .A2 (nx648), .B0 (Dout[6]
         ), .B1 (nx636)) ;
    dff reg_Dout_7 (.Q (Dout[7]), .QB (\$dummy [7]), .D (nx472), .CLK (CLK)) ;
    ao32 ix473 (.Y (nx472), .A0 (Din[7]), .A1 (nx634), .A2 (nx648), .B0 (Dout[7]
         ), .B1 (nx638)) ;
    dff reg_Dout_8 (.Q (Dout[8]), .QB (\$dummy [8]), .D (nx482), .CLK (CLK)) ;
    ao32 ix483 (.Y (nx482), .A0 (Din[8]), .A1 (nx634), .A2 (nx648), .B0 (Dout[8]
         ), .B1 (nx638)) ;
    dff reg_Dout_9 (.Q (Dout[9]), .QB (\$dummy [9]), .D (nx492), .CLK (CLK)) ;
    ao32 ix493 (.Y (nx492), .A0 (Din[9]), .A1 (nx634), .A2 (nx648), .B0 (Dout[9]
         ), .B1 (nx638)) ;
    dff reg_Dout_10 (.Q (Dout[10]), .QB (\$dummy [10]), .D (nx502), .CLK (CLK)
        ) ;
    ao32 ix503 (.Y (nx502), .A0 (Din[10]), .A1 (nx634), .A2 (nx648), .B0 (
         Dout[10]), .B1 (nx638)) ;
    dff reg_Dout_11 (.Q (Dout[11]), .QB (\$dummy [11]), .D (nx512), .CLK (CLK)
        ) ;
    ao32 ix513 (.Y (nx512), .A0 (Din[11]), .A1 (nx634), .A2 (nx648), .B0 (
         Dout[11]), .B1 (nx638)) ;
    dff reg_Dout_12 (.Q (Dout[12]), .QB (\$dummy [12]), .D (nx522), .CLK (CLK)
        ) ;
    ao32 ix523 (.Y (nx522), .A0 (Din[12]), .A1 (nx574), .A2 (nx648), .B0 (
         Dout[12]), .B1 (nx638)) ;
    dff reg_Dout_13 (.Q (Dout[13]), .QB (\$dummy [13]), .D (nx532), .CLK (CLK)
        ) ;
    ao32 ix533 (.Y (nx532), .A0 (Din[13]), .A1 (nx574), .A2 (nx650), .B0 (
         Dout[13]), .B1 (nx638)) ;
    dff reg_Dout_14 (.Q (Dout[14]), .QB (\$dummy [14]), .D (nx542), .CLK (CLK)
        ) ;
    ao32 ix543 (.Y (nx542), .A0 (Din[14]), .A1 (nx574), .A2 (nx650), .B0 (
         Dout[14]), .B1 (nx576)) ;
    dff reg_Dout_15 (.Q (Dout[15]), .QB (\$dummy [15]), .D (nx552), .CLK (CLK)
        ) ;
    ao32 ix553 (.Y (nx552), .A0 (Din[15]), .A1 (nx574), .A2 (nx650), .B0 (
         Dout[15]), .B1 (nx576)) ;
    dff reg_Dout_16 (.Q (Dout[16]), .QB (\$dummy [16]), .D (nx562), .CLK (CLK)
        ) ;
    ao32 ix563 (.Y (nx562), .A0 (Din[16]), .A1 (nx574), .A2 (nx650), .B0 (
         Dout[16]), .B1 (nx576)) ;
    inv01 ix631 (.Y (nx632), .A (RST)) ;
    inv01 ix633 (.Y (nx634), .A (RST)) ;
    nor02_2x ix635 (.Y (nx636), .A0 (RST), .A1 (nx650)) ;
    nor02_2x ix637 (.Y (nx638), .A0 (RST), .A1 (nx650)) ;
    inv01 ix643 (.Y (nx644), .A (EN)) ;
    inv02 ix645 (.Y (nx646), .A (nx644)) ;
    inv02 ix647 (.Y (nx648), .A (nx644)) ;
    inv02 ix649 (.Y (nx650), .A (nx644)) ;
endmodule


module booth_adder_17 ( AdderFirstOperand, AdderSecondOperand, BoothOperand, 
                        BoothP, SelOperand, Operation, AdderResult, 
                        AdderBoothResult ) ;

    input [16:0]AdderFirstOperand ;
    input [16:0]AdderSecondOperand ;
    input [16:0]BoothOperand ;
    input [16:0]BoothP ;
    input SelOperand ;
    input Operation ;
    output [16:0]AdderResult ;
    output [16:0]AdderBoothResult ;

    wire FirstOperand_16, FirstOperand_15, FirstOperand_14, FirstOperand_13, 
         FirstOperand_12, FirstOperand_11, FirstOperand_10, FirstOperand_9, 
         FirstOperand_8, FirstOperand_7, FirstOperand_6, FirstOperand_5, 
         FirstOperand_4, FirstOperand_3, FirstOperand_2, FirstOperand_1, 
         FirstOperand_0, SecondOperand_16, SecondOperand_15, SecondOperand_14, 
         SecondOperand_13, SecondOperand_12, SecondOperand_11, SecondOperand_10, 
         SecondOperand_9, SecondOperand_8, SecondOperand_7, SecondOperand_6, 
         SecondOperand_5, SecondOperand_4, SecondOperand_3, SecondOperand_2, 
         SecondOperand_1, SecondOperand_0, nx224, nx227, nx229, nx231, nx233, 
         nx235, nx237, nx239, nx241, nx243;
    wire [0:0] \$dummy ;




    adder_17 ADDER (.A ({FirstOperand_16,FirstOperand_15,FirstOperand_14,
             FirstOperand_13,FirstOperand_12,FirstOperand_11,FirstOperand_10,
             FirstOperand_9,FirstOperand_8,FirstOperand_7,FirstOperand_6,
             FirstOperand_5,FirstOperand_4,FirstOperand_3,FirstOperand_2,
             FirstOperand_1,FirstOperand_0}), .B ({SecondOperand_16,
             SecondOperand_15,SecondOperand_14,SecondOperand_13,SecondOperand_12
             ,SecondOperand_11,SecondOperand_10,SecondOperand_9,SecondOperand_8,
             SecondOperand_7,SecondOperand_6,SecondOperand_5,SecondOperand_4,
             SecondOperand_3,SecondOperand_2,SecondOperand_1,SecondOperand_0}), 
             .Cin (AdderBoothResult[16]), .Sum ({AdderResult[16],AdderResult[15]
             ,AdderResult[14],AdderResult[13],AdderResult[12],AdderResult[11],
             AdderResult[10],AdderResult[9],AdderResult[8],AdderResult[7],
             AdderResult[6],AdderResult[5],AdderResult[4],AdderResult[3],
             AdderResult[2],AdderResult[1],AdderResult[0]}), .Cout (\$dummy [0])
             ) ;
    fake_gnd ix47 (.Y (AdderBoothResult[16])) ;
    mux21_ni ix137 (.Y (SecondOperand_0), .A0 (AdderSecondOperand[0]), .A1 (
             BoothP[0]), .S0 (nx235)) ;
    mux21_ni ix145 (.Y (SecondOperand_1), .A0 (AdderSecondOperand[1]), .A1 (
             BoothP[1]), .S0 (nx235)) ;
    mux21_ni ix153 (.Y (SecondOperand_2), .A0 (AdderSecondOperand[2]), .A1 (
             BoothP[2]), .S0 (nx235)) ;
    mux21_ni ix161 (.Y (SecondOperand_3), .A0 (AdderSecondOperand[3]), .A1 (
             BoothP[3]), .S0 (nx235)) ;
    mux21_ni ix169 (.Y (SecondOperand_4), .A0 (AdderSecondOperand[4]), .A1 (
             BoothP[4]), .S0 (nx235)) ;
    mux21_ni ix177 (.Y (SecondOperand_5), .A0 (AdderSecondOperand[5]), .A1 (
             BoothP[5]), .S0 (nx235)) ;
    mux21_ni ix185 (.Y (SecondOperand_6), .A0 (AdderSecondOperand[6]), .A1 (
             BoothP[6]), .S0 (nx235)) ;
    mux21_ni ix193 (.Y (SecondOperand_7), .A0 (AdderSecondOperand[7]), .A1 (
             BoothP[7]), .S0 (nx237)) ;
    mux21_ni ix201 (.Y (SecondOperand_8), .A0 (AdderSecondOperand[8]), .A1 (
             BoothP[8]), .S0 (nx237)) ;
    mux21_ni ix209 (.Y (SecondOperand_9), .A0 (AdderSecondOperand[9]), .A1 (
             BoothP[9]), .S0 (nx237)) ;
    mux21_ni ix217 (.Y (SecondOperand_10), .A0 (AdderSecondOperand[10]), .A1 (
             BoothP[10]), .S0 (nx237)) ;
    mux21_ni ix225 (.Y (SecondOperand_11), .A0 (AdderSecondOperand[11]), .A1 (
             BoothP[11]), .S0 (nx237)) ;
    mux21_ni ix233 (.Y (SecondOperand_12), .A0 (AdderSecondOperand[12]), .A1 (
             BoothP[12]), .S0 (nx237)) ;
    mux21_ni ix241 (.Y (SecondOperand_13), .A0 (AdderSecondOperand[13]), .A1 (
             BoothP[13]), .S0 (nx237)) ;
    mux21_ni ix249 (.Y (SecondOperand_14), .A0 (AdderSecondOperand[14]), .A1 (
             BoothP[14]), .S0 (nx239)) ;
    mux21_ni ix257 (.Y (SecondOperand_15), .A0 (AdderSecondOperand[15]), .A1 (
             BoothP[15]), .S0 (nx239)) ;
    nor02ii ix261 (.Y (FirstOperand_0), .A0 (nx239), .A1 (AdderFirstOperand[0])
            ) ;
    nor02ii ix265 (.Y (FirstOperand_1), .A0 (nx239), .A1 (AdderFirstOperand[1])
            ) ;
    nor02ii ix269 (.Y (FirstOperand_2), .A0 (nx239), .A1 (AdderFirstOperand[2])
            ) ;
    nor02ii ix273 (.Y (FirstOperand_3), .A0 (nx239), .A1 (AdderFirstOperand[3])
            ) ;
    nor02ii ix277 (.Y (FirstOperand_4), .A0 (nx239), .A1 (AdderFirstOperand[4])
            ) ;
    nor02ii ix281 (.Y (FirstOperand_5), .A0 (nx241), .A1 (AdderFirstOperand[5])
            ) ;
    nor02ii ix285 (.Y (FirstOperand_6), .A0 (nx241), .A1 (AdderFirstOperand[6])
            ) ;
    nor02ii ix289 (.Y (FirstOperand_7), .A0 (nx241), .A1 (AdderFirstOperand[7])
            ) ;
    nor02ii ix293 (.Y (FirstOperand_8), .A0 (nx241), .A1 (AdderFirstOperand[8])
            ) ;
    mux21_ni ix303 (.Y (FirstOperand_9), .A0 (AdderFirstOperand[9]), .A1 (
             BoothOperand[9]), .S0 (nx241)) ;
    mux21_ni ix311 (.Y (FirstOperand_10), .A0 (AdderFirstOperand[10]), .A1 (
             BoothOperand[10]), .S0 (nx241)) ;
    mux21_ni ix319 (.Y (FirstOperand_11), .A0 (AdderFirstOperand[11]), .A1 (
             BoothOperand[11]), .S0 (nx241)) ;
    mux21_ni ix327 (.Y (FirstOperand_12), .A0 (AdderFirstOperand[12]), .A1 (
             BoothOperand[12]), .S0 (nx243)) ;
    mux21_ni ix335 (.Y (FirstOperand_13), .A0 (AdderFirstOperand[13]), .A1 (
             BoothOperand[13]), .S0 (nx243)) ;
    mux21_ni ix343 (.Y (FirstOperand_14), .A0 (AdderFirstOperand[14]), .A1 (
             BoothOperand[14]), .S0 (nx243)) ;
    mux21_ni ix351 (.Y (FirstOperand_15), .A0 (AdderFirstOperand[15]), .A1 (
             BoothOperand[15]), .S0 (nx243)) ;
    mux21_ni ix7 (.Y (AdderBoothResult[0]), .A0 (BoothP[1]), .A1 (AdderResult[1]
             ), .S0 (nx227)) ;
    mux21_ni ix15 (.Y (AdderBoothResult[1]), .A0 (BoothP[2]), .A1 (
             AdderResult[2]), .S0 (nx227)) ;
    mux21_ni ix23 (.Y (AdderBoothResult[2]), .A0 (BoothP[3]), .A1 (
             AdderResult[3]), .S0 (nx227)) ;
    mux21_ni ix31 (.Y (AdderBoothResult[3]), .A0 (BoothP[4]), .A1 (
             AdderResult[4]), .S0 (nx227)) ;
    mux21_ni ix39 (.Y (AdderBoothResult[4]), .A0 (BoothP[5]), .A1 (
             AdderResult[5]), .S0 (nx227)) ;
    mux21_ni ix49 (.Y (AdderBoothResult[5]), .A0 (BoothP[6]), .A1 (
             AdderResult[6]), .S0 (nx227)) ;
    mux21_ni ix55 (.Y (AdderBoothResult[6]), .A0 (BoothP[7]), .A1 (
             AdderResult[7]), .S0 (nx227)) ;
    mux21_ni ix63 (.Y (AdderBoothResult[7]), .A0 (BoothP[8]), .A1 (
             AdderResult[8]), .S0 (nx229)) ;
    mux21_ni ix71 (.Y (AdderBoothResult[8]), .A0 (BoothP[9]), .A1 (
             AdderResult[9]), .S0 (nx229)) ;
    mux21_ni ix79 (.Y (AdderBoothResult[9]), .A0 (BoothP[10]), .A1 (
             AdderResult[10]), .S0 (nx229)) ;
    mux21_ni ix87 (.Y (AdderBoothResult[10]), .A0 (BoothP[11]), .A1 (
             AdderResult[11]), .S0 (nx229)) ;
    mux21_ni ix95 (.Y (AdderBoothResult[11]), .A0 (BoothP[12]), .A1 (
             AdderResult[12]), .S0 (nx229)) ;
    mux21_ni ix103 (.Y (AdderBoothResult[12]), .A0 (BoothP[13]), .A1 (
             AdderResult[13]), .S0 (nx229)) ;
    mux21_ni ix111 (.Y (AdderBoothResult[13]), .A0 (BoothP[14]), .A1 (
             AdderResult[14]), .S0 (nx229)) ;
    mux21_ni ix119 (.Y (AdderBoothResult[14]), .A0 (BoothP[15]), .A1 (
             AdderResult[15]), .S0 (nx231)) ;
    mux21_ni ix127 (.Y (AdderBoothResult[15]), .A0 (BoothP[16]), .A1 (
             AdderResult[16]), .S0 (nx231)) ;
    and02 ix129 (.Y (SecondOperand_16), .A0 (nx243), .A1 (BoothP[16])) ;
    and02 ix295 (.Y (FirstOperand_16), .A0 (nx243), .A1 (BoothOperand[16])) ;
    inv01 ix223 (.Y (nx224), .A (Operation)) ;
    inv02 ix226 (.Y (nx227), .A (nx224)) ;
    inv02 ix228 (.Y (nx229), .A (nx224)) ;
    inv02 ix230 (.Y (nx231), .A (nx224)) ;
    inv01 ix232 (.Y (nx233), .A (SelOperand)) ;
    inv02 ix234 (.Y (nx235), .A (nx233)) ;
    inv02 ix236 (.Y (nx237), .A (nx233)) ;
    inv02 ix238 (.Y (nx239), .A (nx233)) ;
    inv02 ix240 (.Y (nx241), .A (nx233)) ;
    inv02 ix242 (.Y (nx243), .A (nx233)) ;
endmodule


module adder_17 ( A, B, Cin, Sum, Cout ) ;

    input [16:0]A ;
    input [16:0]B ;
    input Cin ;
    output [16:0]Sum ;
    output Cout ;

    wire nx2, nx16, nx18, nx32, nx34, nx48, nx50, nx64, nx66, nx80, nx82, nx96, 
         nx98, nx112, nx114, nx122, nx105, nx107, nx111, nx115, nx121, nx123, 
         nx127, nx131, nx137, nx139, nx143, nx147, nx153, nx155, nx159, nx163, 
         nx167, nx169, nx172, nx175, nx179, nx181, nx184, nx187, nx191, nx193, 
         nx196, nx199, nx203, nx205, nx208;



    fake_gnd ix58 (.Y (Cout)) ;
    xor2 ix161 (.Y (Sum[0]), .A0 (B[0]), .A1 (A[0])) ;
    xor2 ix155 (.Y (Sum[1]), .A0 (nx105), .A1 (nx107)) ;
    nand02 ix106 (.Y (nx105), .A0 (B[0]), .A1 (A[0])) ;
    xnor2 ix108 (.Y (nx107), .A0 (A[1]), .A1 (B[1])) ;
    xor2 ix153 (.Y (Sum[2]), .A0 (nx111), .A1 (nx115)) ;
    aoi32 ix112 (.Y (nx111), .A0 (B[0]), .A1 (A[0]), .A2 (nx2), .B0 (B[1]), .B1 (
          A[1])) ;
    xnor2 ix116 (.Y (nx115), .A0 (A[2]), .A1 (B[2])) ;
    xnor2 ix151 (.Y (Sum[3]), .A0 (nx16), .A1 (nx123)) ;
    oai21 ix17 (.Y (nx16), .A0 (nx111), .A1 (nx115), .B0 (nx121)) ;
    nand02 ix122 (.Y (nx121), .A0 (B[2]), .A1 (A[2])) ;
    xnor2 ix124 (.Y (nx123), .A0 (A[3]), .A1 (B[3])) ;
    xor2 ix149 (.Y (Sum[4]), .A0 (nx127), .A1 (nx131)) ;
    aoi22 ix128 (.Y (nx127), .A0 (B[3]), .A1 (A[3]), .B0 (nx16), .B1 (nx18)) ;
    xnor2 ix132 (.Y (nx131), .A0 (A[4]), .A1 (B[4])) ;
    xnor2 ix147 (.Y (Sum[5]), .A0 (nx32), .A1 (nx139)) ;
    oai21 ix33 (.Y (nx32), .A0 (nx127), .A1 (nx131), .B0 (nx137)) ;
    nand02 ix138 (.Y (nx137), .A0 (B[4]), .A1 (A[4])) ;
    xnor2 ix140 (.Y (nx139), .A0 (A[5]), .A1 (B[5])) ;
    xor2 ix145 (.Y (Sum[6]), .A0 (nx143), .A1 (nx147)) ;
    aoi22 ix144 (.Y (nx143), .A0 (B[5]), .A1 (A[5]), .B0 (nx32), .B1 (nx34)) ;
    xnor2 ix148 (.Y (nx147), .A0 (A[6]), .A1 (B[6])) ;
    xnor2 ix143 (.Y (Sum[7]), .A0 (nx48), .A1 (nx155)) ;
    oai21 ix49 (.Y (nx48), .A0 (nx143), .A1 (nx147), .B0 (nx153)) ;
    nand02 ix154 (.Y (nx153), .A0 (B[6]), .A1 (A[6])) ;
    xnor2 ix156 (.Y (nx155), .A0 (A[7]), .A1 (B[7])) ;
    xor2 ix141 (.Y (Sum[8]), .A0 (nx159), .A1 (nx163)) ;
    aoi22 ix160 (.Y (nx159), .A0 (B[7]), .A1 (A[7]), .B0 (nx48), .B1 (nx50)) ;
    xnor2 ix164 (.Y (nx163), .A0 (A[8]), .A1 (B[8])) ;
    xnor2 ix139 (.Y (Sum[9]), .A0 (nx64), .A1 (nx169)) ;
    oai21 ix65 (.Y (nx64), .A0 (nx159), .A1 (nx163), .B0 (nx167)) ;
    nand02 ix168 (.Y (nx167), .A0 (B[8]), .A1 (A[8])) ;
    xnor2 ix170 (.Y (nx169), .A0 (A[9]), .A1 (B[9])) ;
    xor2 ix137 (.Y (Sum[10]), .A0 (nx172), .A1 (nx175)) ;
    aoi22 ix173 (.Y (nx172), .A0 (B[9]), .A1 (A[9]), .B0 (nx64), .B1 (nx66)) ;
    xnor2 ix176 (.Y (nx175), .A0 (A[10]), .A1 (B[10])) ;
    xnor2 ix135 (.Y (Sum[11]), .A0 (nx80), .A1 (nx181)) ;
    oai21 ix81 (.Y (nx80), .A0 (nx172), .A1 (nx175), .B0 (nx179)) ;
    nand02 ix180 (.Y (nx179), .A0 (B[10]), .A1 (A[10])) ;
    xnor2 ix182 (.Y (nx181), .A0 (A[11]), .A1 (B[11])) ;
    xor2 ix133 (.Y (Sum[12]), .A0 (nx184), .A1 (nx187)) ;
    aoi22 ix185 (.Y (nx184), .A0 (B[11]), .A1 (A[11]), .B0 (nx80), .B1 (nx82)) ;
    xnor2 ix188 (.Y (nx187), .A0 (A[12]), .A1 (B[12])) ;
    xnor2 ix131 (.Y (Sum[13]), .A0 (nx96), .A1 (nx193)) ;
    oai21 ix97 (.Y (nx96), .A0 (nx184), .A1 (nx187), .B0 (nx191)) ;
    nand02 ix192 (.Y (nx191), .A0 (B[12]), .A1 (A[12])) ;
    xnor2 ix194 (.Y (nx193), .A0 (A[13]), .A1 (B[13])) ;
    xor2 ix129 (.Y (Sum[14]), .A0 (nx196), .A1 (nx199)) ;
    aoi22 ix197 (.Y (nx196), .A0 (B[13]), .A1 (A[13]), .B0 (nx96), .B1 (nx98)) ;
    xnor2 ix200 (.Y (nx199), .A0 (A[14]), .A1 (B[14])) ;
    xnor2 ix127 (.Y (Sum[15]), .A0 (nx112), .A1 (nx205)) ;
    oai21 ix113 (.Y (nx112), .A0 (nx196), .A1 (nx199), .B0 (nx203)) ;
    nand02 ix204 (.Y (nx203), .A0 (B[14]), .A1 (A[14])) ;
    xnor2 ix206 (.Y (nx205), .A0 (A[15]), .A1 (B[15])) ;
    xnor2 ix125 (.Y (Sum[16]), .A0 (nx208), .A1 (nx122)) ;
    aoi22 ix209 (.Y (nx208), .A0 (B[15]), .A1 (A[15]), .B0 (nx112), .B1 (nx114)
          ) ;
    xor2 ix123 (.Y (nx122), .A0 (A[16]), .A1 (B[16])) ;
    inv01 ix115 (.Y (nx114), .A (nx205)) ;
    inv01 ix99 (.Y (nx98), .A (nx193)) ;
    inv01 ix83 (.Y (nx82), .A (nx181)) ;
    inv01 ix67 (.Y (nx66), .A (nx169)) ;
    inv01 ix51 (.Y (nx50), .A (nx155)) ;
    inv01 ix35 (.Y (nx34), .A (nx139)) ;
    inv01 ix19 (.Y (nx18), .A (nx123)) ;
    inv01 ix3 (.Y (nx2), .A (nx107)) ;
endmodule


module controller ( CLK, RST, Start, FilterSize, Stride, Instr, CalcFinished, 
                    Calc, MemRD, MemWR, MemAddr, CacheFilterWR, CacheWindowWR, 
                    FirstCycle, Done ) ;

    input CLK ;
    input RST ;
    input Start ;
    input FilterSize ;
    input Stride ;
    input Instr ;
    input CalcFinished ;
    output Calc ;
    output MemRD ;
    output MemWR ;
    output [17:0]MemAddr ;
    output CacheFilterWR ;
    output CacheWindowWR ;
    output FirstCycle ;
    output Done ;

    wire CurCol_5, nx487, CurRow_5, nx488, CurRow_4, CurRow_3, CurRow_2, nx14, 
         nx20, nx34, nx46, nx493, nx72, nx82, nx102, nx110, CurRow_7, CurRow_6, 
         nx118, nx138, nx162, nx164, nx178, nx188, nx196, nx224, nx230, nx246, 
         nx264, nx276, CurCol_4, CurCol_3, CurCol_2, CurCol_1, CurCol_0, nx497, 
         nx296, nx499, nx322, nx332, nx503, nx358, nx368, nx388, nx396, CurCol_7, 
         CurCol_6, nx410, nx422, nx448, nx456, nx462, nx472, nx478, nx500, nx522, 
         nx524, nx540, nx558, nx560, nx576, nx594, nx596, nx612, nx628, nx646, 
         nx662, nx668, nx690, nx696, nx718, nx515, nx525, nx535, nx545, nx555, 
         nx565, nx575, nx585, nx595, nx605, nx615, nx625, nx635, nx645, nx655, 
         nx665, nx683, nx695, nx697, nx703, nx707, nx709, nx711, nx721, nx727, 
         nx729, nx733, nx737, nx739, nx745, nx748, nx754, nx758, nx760, nx764, 
         nx768, nx771, nx775, nx777, nx780, nx784, nx787, nx796, nx800, nx802, 
         nx805, nx809, nx812, nx815, nx818, nx823, nx826, nx829, nx832, nx836, 
         nx838, nx842, nx844, nx850, nx852, nx856, nx858, nx861, nx865, nx867, 
         nx870, nx873, nx875, nx879, nx883, nx894, nx898, nx907, nx910, nx917, 
         nx920, nx923, nx925, nx928, nx932, nx935, nx938, nx942, nx946, nx949, 
         nx952, nx956, nx962, nx964, nx971, nx975, nx977, nx983, nx985, nx988, 
         nx998, nx1000, nx1002, nx1004, nx1006, nx1008, nx1010, nx1012, nx1014, 
         nx1016, nx1018, nx1020, nx1022, nx1028, nx1030, nx1032, nx1034, nx1036, 
         nx1042, nx1044, nx1046, nx1048, nx1050, nx1052, nx1054, nx1056, nx1058, 
         nx1060, nx1062;
    wire [5:0] \$dummy ;




    assign MemAddr[16] = MemWR ;
    and03 ix277 (.Y (nx276), .A0 (nx683), .A1 (CalcFinished), .A2 (Calc)) ;
    aoi21 ix684 (.Y (nx683), .A0 (Start), .A1 (nx487), .B0 (RST)) ;
    nor03_2x ix397 (.Y (nx396), .A0 (nx695), .A1 (nx1022), .A2 (nx388)) ;
    nand02 ix698 (.Y (nx697), .A0 (CurCol_4), .A1 (nx503)) ;
    oai21 ix636 (.Y (nx635), .A0 (nx703), .A1 (nx1010), .B0 (nx898)) ;
    dff COL_reg_Dout_4 (.Q (CurCol_4), .QB (nx703), .D (nx635), .CLK (CLK)) ;
    aoi21 ix708 (.Y (nx707), .A0 (nx709), .A1 (MemRD), .B0 (nx1022)) ;
    oai21 ix710 (.Y (nx709), .A0 (nx711), .A1 (nx894), .B0 (nx748)) ;
    dff ROW_reg_Dout_0 (.Q (\$dummy [0]), .QB (nx711), .D (nx515), .CLK (CLK)) ;
    oai21 ix15 (.Y (nx14), .A0 (nx721), .A1 (nx745), .B0 (nx683)) ;
    aoi22 ix728 (.Y (nx727), .A0 (nx729), .A1 (FirstCycle), .B0 (CacheFilterWR)
          , .B1 (nx188)) ;
    inv01 ix730 (.Y (nx729), .A (Instr)) ;
    nor04 ix213 (.Y (FirstCycle), .A0 (nx733), .A1 (Calc), .A2 (nx998), .A3 (
          MemRD)) ;
    inv01 ix734 (.Y (nx733), .A (Start)) ;
    dff STATE_reg_Dout_3 (.Q (Calc), .QB (\$dummy [1]), .D (nx264), .CLK (CLK)
        ) ;
    aoi22 ix738 (.Y (nx737), .A0 (nx739), .A1 (Calc), .B0 (CacheWindowWR), .B1 (
          nx224)) ;
    inv01 ix740 (.Y (nx739), .A (CalcFinished)) ;
    dff STATE_reg_Dout_1 (.Q (CacheWindowWR), .QB (\$dummy [2]), .D (nx246), .CLK (
        CLK)) ;
    aoi221 ix746 (.Y (nx745), .A0 (CacheFilterWR), .A1 (nx748), .B0 (nx998), .B1 (
           nx796), .C0 (nx230)) ;
    dff STATE_reg_Dout_0 (.Q (CacheFilterWR), .QB (nx721), .D (nx196), .CLK (CLK
        )) ;
    nand04 ix749 (.Y (nx748), .A0 (nx162), .A1 (nx178), .A2 (nx758), .A3 (nx764)
           ) ;
    nor03_2x ix111 (.Y (nx110), .A0 (nx754), .A1 (nx102), .A2 (nx1020)) ;
    aoi21 ix755 (.Y (nx754), .A0 (CurRow_4), .A1 (nx493), .B0 (CurRow_5)) ;
    oai21 ix556 (.Y (nx555), .A0 (nx758), .A1 (nx1008), .B0 (nx760)) ;
    dff ROW_reg_Dout_4 (.Q (CurRow_4), .QB (nx758), .D (nx555), .CLK (CLK)) ;
    nand04 ix761 (.Y (nx760), .A0 (nx82), .A1 (nx844), .A2 (nx1030), .A3 (nx1010
           )) ;
    or02 ix83 (.Y (nx82), .A0 (nx493), .A1 (CurRow_4)) ;
    nor03_2x ix73 (.Y (nx72), .A0 (nx768), .A1 (nx493), .A2 (nx1020)) ;
    dff ROW_reg_Dout_3 (.Q (CurRow_3), .QB (nx764), .D (nx545), .CLK (CLK)) ;
    oai21 ix536 (.Y (nx535), .A0 (nx775), .A1 (nx1008), .B0 (nx777)) ;
    dff ROW_reg_Dout_2 (.Q (CurRow_2), .QB (nx775), .D (nx535), .CLK (CLK)) ;
    nand04 ix778 (.Y (nx777), .A0 (nx46), .A1 (nx771), .A2 (nx1030), .A3 (nx1010
           )) ;
    nand02 ix47 (.Y (nx46), .A0 (nx780), .A1 (nx775)) ;
    oai21 ix785 (.Y (nx784), .A0 (nx1016), .A1 (nx1012), .B0 (nx34)) ;
    aoi21 ix35 (.Y (nx34), .A0 (nx1012), .A1 (nx1016), .B0 (nx1020)) ;
    dff ROW_reg_Dout_1 (.Q (\$dummy [3]), .QB (nx787), .D (nx525), .CLK (CLK)) ;
    nand04 ix797 (.Y (nx796), .A0 (CurCol_5), .A1 (CurCol_7), .A2 (CurCol_6), .A3 (
           nx456)) ;
    oai21 ix666 (.Y (nx665), .A0 (nx800), .A1 (nx1008), .B0 (nx802)) ;
    dff COL_reg_Dout_7 (.Q (CurCol_7), .QB (nx800), .D (nx665), .CLK (CLK)) ;
    nand03 ix803 (.Y (nx802), .A0 (nx1030), .A1 (nx422), .A2 (nx1008)) ;
    nand02 ix806 (.Y (nx805), .A0 (CurCol_6), .A1 (nx388)) ;
    oai21 ix810 (.Y (nx809), .A0 (nx388), .A1 (CurCol_6), .B0 (nx410)) ;
    dff COL_reg_Dout_5 (.Q (CurCol_5), .QB (nx812), .D (nx645), .CLK (CLK)) ;
    aoi21 ix411 (.Y (nx410), .A0 (CurCol_6), .A1 (nx388), .B0 (nx1020)) ;
    dff COL_reg_Dout_6 (.Q (CurCol_6), .QB (nx815), .D (nx655), .CLK (CLK)) ;
    nor03_2x ix457 (.Y (nx456), .A0 (nx818), .A1 (nx703), .A2 (nx875)) ;
    aoi32 ix819 (.Y (nx818), .A0 (CurCol_0), .A1 (FilterSize), .A2 (CurCol_1), .B0 (
          CurCol_2), .B1 (nx448)) ;
    dff COL_reg_Dout_0 (.Q (CurCol_0), .QB (nx852), .D (nx595), .CLK (CLK)) ;
    xnor2 ix824 (.Y (nx823), .A0 (nx138), .A1 (nx497)) ;
    oai21 ix586 (.Y (nx585), .A0 (nx826), .A1 (nx1008), .B0 (nx829)) ;
    nand02 ix833 (.Y (nx832), .A0 (CurRow_6), .A1 (nx102)) ;
    oai21 ix576 (.Y (nx575), .A0 (nx836), .A1 (nx1008), .B0 (nx838)) ;
    dff ROW_reg_Dout_6 (.Q (CurRow_6), .QB (nx836), .D (nx575), .CLK (CLK)) ;
    nand04 ix839 (.Y (nx838), .A0 (nx118), .A1 (nx832), .A2 (nx1030), .A3 (
           nx1008)) ;
    or02 ix119 (.Y (nx118), .A0 (nx102), .A1 (CurRow_6)) ;
    dff ROW_reg_Dout_5 (.Q (CurRow_5), .QB (nx842), .D (nx565), .CLK (CLK)) ;
    nand02 ix845 (.Y (nx844), .A0 (CurRow_4), .A1 (nx493)) ;
    dff ROW_reg_Dout_7 (.Q (CurRow_7), .QB (nx826), .D (nx585), .CLK (CLK)) ;
    nand02 ix851 (.Y (nx850), .A0 (Stride), .A1 (nx138)) ;
    nor03_2x ix323 (.Y (nx322), .A0 (nx856), .A1 (nx1020), .A2 (nx499)) ;
    oai21 ix859 (.Y (nx858), .A0 (CurCol_0), .A1 (Stride), .B0 (nx138)) ;
    dff COL_reg_Dout_1 (.Q (CurCol_1), .QB (nx861), .D (nx605), .CLK (CLK)) ;
    oai21 ix616 (.Y (nx615), .A0 (nx865), .A1 (nx1010), .B0 (nx867)) ;
    dff COL_reg_Dout_2 (.Q (CurCol_2), .QB (nx865), .D (nx615), .CLK (CLK)) ;
    nand04 ix868 (.Y (nx867), .A0 (nx332), .A1 (nx1030), .A2 (nx870), .A3 (
           nx1010)) ;
    or02 ix333 (.Y (nx332), .A0 (nx499), .A1 (CurCol_2)) ;
    nand02 ix871 (.Y (nx870), .A0 (CurCol_2), .A1 (nx499)) ;
    inv01 ix874 (.Y (nx873), .A (FilterSize)) ;
    nor03_2x ix359 (.Y (nx358), .A0 (nx879), .A1 (nx1020), .A2 (nx503)) ;
    dff COL_reg_Dout_3 (.Q (CurCol_3), .QB (nx875), .D (nx625), .CLK (CLK)) ;
    aoi22 ix884 (.Y (nx883), .A0 (Instr), .A1 (FirstCycle), .B0 (CacheWindowWR)
          , .B1 (nx709)) ;
    aoi21 ix179 (.Y (nx178), .A0 (nx873), .A1 (nx1012), .B0 (CurRow_2)) ;
    or02 ix205 (.Y (MemRD), .A0 (CacheFilterWR), .A1 (CacheWindowWR)) ;
    inv01 ix895 (.Y (nx894), .A (Stride)) ;
    dff STATE_reg_Dout_2 (.Q (MemWR), .QB (\$dummy [4]), .D (nx276), .CLK (CLK)
        ) ;
    nand04 ix899 (.Y (nx898), .A0 (nx368), .A1 (nx1030), .A2 (nx697), .A3 (
           nx1010)) ;
    or02 ix369 (.Y (nx368), .A0 (nx503), .A1 (CurCol_4)) ;
    dff STATE_reg_Dout_4 (.Q (Done), .QB (\$dummy [5]), .D (nx462), .CLK (CLK)
        ) ;
    nor03_2x ix463 (.Y (nx462), .A0 (nx796), .A1 (Start), .A2 (RST)) ;
    oai21 ix497 (.Y (MemAddr[0]), .A0 (nx852), .A1 (nx1034), .B0 (nx907)) ;
    aoi32 ix908 (.Y (nx907), .A0 (nx478), .A1 (nx998), .A2 (nx910), .B0 (nx1016)
          , .B1 (nx1004)) ;
    nand02 ix479 (.Y (nx478), .A0 (nx852), .A1 (FilterSize)) ;
    xor2 ix501 (.Y (nx500), .A0 (nx910), .A1 (nx917)) ;
    oai21 ix537 (.Y (MemAddr[2]), .A0 (nx865), .A1 (nx1034), .B0 (nx920)) ;
    aoi32 ix921 (.Y (nx920), .A0 (nx522), .A1 (nx1000), .A2 (nx925), .B0 (
          CurRow_2), .B1 (nx1004)) ;
    nand02 ix523 (.Y (nx522), .A0 (nx923), .A1 (nx865)) ;
    oai21 ix924 (.Y (nx923), .A0 (FilterSize), .A1 (CurCol_0), .B0 (CurCol_1)) ;
    oai21 ix555 (.Y (MemAddr[3]), .A0 (nx875), .A1 (nx1034), .B0 (nx928)) ;
    aoi32 ix929 (.Y (nx928), .A0 (nx540), .A1 (nx1000), .A2 (nx932), .B0 (
          CurRow_3), .B1 (nx1004)) ;
    or02 ix541 (.Y (nx540), .A0 (nx524), .A1 (CurCol_3)) ;
    nand02 ix933 (.Y (nx932), .A0 (CurCol_3), .A1 (nx524)) ;
    oai21 ix573 (.Y (MemAddr[4]), .A0 (nx703), .A1 (nx1034), .B0 (nx935)) ;
    aoi32 ix936 (.Y (nx935), .A0 (nx558), .A1 (nx1000), .A2 (nx938), .B0 (
          CurRow_4), .B1 (nx1004)) ;
    nand02 ix559 (.Y (nx558), .A0 (nx932), .A1 (nx703)) ;
    oai21 ix591 (.Y (MemAddr[5]), .A0 (nx812), .A1 (nx1034), .B0 (nx942)) ;
    aoi32 ix943 (.Y (nx942), .A0 (nx576), .A1 (nx1000), .A2 (nx946), .B0 (
          CurRow_5), .B1 (nx1004)) ;
    or02 ix577 (.Y (nx576), .A0 (nx560), .A1 (CurCol_5)) ;
    nand02 ix947 (.Y (nx946), .A0 (CurCol_5), .A1 (nx560)) ;
    oai21 ix609 (.Y (MemAddr[6]), .A0 (nx815), .A1 (nx1034), .B0 (nx949)) ;
    aoi32 ix950 (.Y (nx949), .A0 (nx594), .A1 (nx1000), .A2 (nx952), .B0 (
          CurRow_6), .B1 (nx1006)) ;
    nand02 ix595 (.Y (nx594), .A0 (nx946), .A1 (nx815)) ;
    oai21 ix625 (.Y (MemAddr[7]), .A0 (nx800), .A1 (nx1034), .B0 (nx956)) ;
    aoi32 ix957 (.Y (nx956), .A0 (nx612), .A1 (nx894), .A2 (nx1000), .B0 (
          CurRow_7), .B1 (nx1006)) ;
    ao32 ix643 (.Y (MemAddr[8]), .A0 (nx628), .A1 (nx1018), .A2 (nx962), .B0 (
         nx1002), .B1 (nx964)) ;
    xnor2 ix647 (.Y (nx646), .A0 (nx964), .A1 (nx164)) ;
    oai21 ix669 (.Y (nx668), .A0 (nx775), .A1 (nx971), .B0 (nx662)) ;
    aoi21 ix972 (.Y (nx971), .A0 (nx1018), .A1 (nx873), .B0 (nx1014)) ;
    nand02 ix663 (.Y (nx662), .A0 (nx971), .A1 (nx775)) ;
    oai22 ix689 (.Y (MemAddr[11]), .A0 (nx1058), .A1 (nx975), .B0 (nx764), .B1 (
          nx1036)) ;
    aoi21 ix976 (.Y (nx975), .A0 (CurRow_3), .A1 (nx662), .B0 (nx977)) ;
    oai21 ix697 (.Y (nx696), .A0 (nx758), .A1 (nx977), .B0 (nx690)) ;
    nand02 ix691 (.Y (nx690), .A0 (nx977), .A1 (nx758)) ;
    oai22 ix717 (.Y (MemAddr[13]), .A0 (nx1058), .A1 (nx983), .B0 (nx842), .B1 (
          nx1036)) ;
    aoi21 ix984 (.Y (nx983), .A0 (CurRow_5), .A1 (nx690), .B0 (nx985)) ;
    oai22 ix731 (.Y (MemAddr[14]), .A0 (nx1058), .A1 (nx988), .B0 (nx836), .B1 (
          nx1036)) ;
    nand02 ix719 (.Y (nx718), .A0 (nx985), .A1 (nx836)) ;
    inv01 ix953 (.Y (nx952), .A (nx596)) ;
    inv01 ix939 (.Y (nx938), .A (nx560)) ;
    inv01 ix926 (.Y (nx925), .A (nx524)) ;
    inv01 ix231 (.Y (nx230), .A (nx883)) ;
    inv01 ix225 (.Y (nx224), .A (nx709)) ;
    inv01 ix189 (.Y (nx188), .A (nx748)) ;
    inv01 ix459 (.Y (nx487), .A (nx796)) ;
    inv01 ix963 (.Y (nx962), .A (MemAddr[17])) ;
    inv02 ix997 (.Y (nx998), .A (nx1058)) ;
    inv02 ix999 (.Y (nx1000), .A (nx1058)) ;
    inv02 ix1001 (.Y (nx1002), .A (nx1058)) ;
    inv01 ix1003 (.Y (nx1004), .A (nx962)) ;
    inv01 ix1005 (.Y (nx1006), .A (nx962)) ;
    inv02 ix1007 (.Y (nx1008), .A (nx1028)) ;
    inv02 ix1009 (.Y (nx1010), .A (nx1028)) ;
    inv02 ix1011 (.Y (nx1012), .A (nx787)) ;
    inv02 ix1013 (.Y (nx1014), .A (nx787)) ;
    inv02 ix1015 (.Y (nx1016), .A (nx711)) ;
    inv02 ix1017 (.Y (nx1018), .A (nx711)) ;
    inv02 ix1019 (.Y (nx1020), .A (nx1032)) ;
    inv02 ix1021 (.Y (nx1022), .A (nx1032)) ;
    inv02 ix1027 (.Y (nx1028), .A (nx488)) ;
    inv02 ix1029 (.Y (nx1030), .A (nx14)) ;
    inv02 ix1031 (.Y (nx1032), .A (nx14)) ;
    inv02 ix1033 (.Y (nx1034), .A (nx472)) ;
    inv02 ix1035 (.Y (nx1036), .A (nx472)) ;
    nor02ii ix491 (.Y (MemAddr[17]), .A0 (CacheWindowWR), .A1 (nx1058)) ;
    mux21_ni ix646 (.Y (nx645), .A0 (CurCol_5), .A1 (nx396), .S0 (nx1054)) ;
    and02 ix696 (.Y (nx695), .A0 (nx812), .A1 (nx697)) ;
    mux21_ni ix516 (.Y (nx515), .A0 (nx1016), .A1 (nx20), .S0 (nx1054)) ;
    and02 ix21 (.Y (nx20), .A0 (nx711), .A1 (nx1032)) ;
    nor02ii ix197 (.Y (nx196), .A0 (nx727), .A1 (nx683)) ;
    nor02ii ix265 (.Y (nx264), .A0 (nx737), .A1 (nx683)) ;
    nor02ii ix247 (.Y (nx246), .A0 (nx745), .A1 (nx683)) ;
    and03 ix163 (.Y (nx162), .A0 (nx842), .A1 (nx826), .A2 (nx836)) ;
    mux21_ni ix566 (.Y (nx565), .A0 (CurRow_5), .A1 (nx110), .S0 (nx1054)) ;
    nor02ii ix81 (.Y (nx493), .A0 (nx771), .A1 (CurRow_3)) ;
    mux21_ni ix546 (.Y (nx545), .A0 (CurRow_3), .A1 (nx72), .S0 (nx1054)) ;
    and02 ix769 (.Y (nx768), .A0 (nx764), .A1 (nx771)) ;
    or03 ix772 (.Y (nx771), .A0 (nx775), .A1 (nx787), .A2 (nx711)) ;
    or02 ix781 (.Y (nx780), .A0 (nx787), .A1 (nx711)) ;
    mux21 ix526 (.Y (nx525), .A0 (nx787), .A1 (nx784), .S0 (nx1054)) ;
    nand02 ix790 (.Y (nx488), .A0 (nx1060), .A1 (nx707)) ;
    xor2 ix423 (.Y (nx422), .A0 (nx800), .A1 (nx805)) ;
    mux21 ix656 (.Y (nx655), .A0 (nx815), .A1 (nx809), .S0 (nx1054)) ;
    nor02ii ix389 (.Y (nx388), .A0 (nx697), .A1 (CurCol_5)) ;
    mux21_ni ix596 (.Y (nx595), .A0 (CurCol_0), .A1 (nx296), .S0 (nx1054)) ;
    nor02ii ix297 (.Y (nx296), .A0 (nx823), .A1 (nx1032)) ;
    nor02ii ix139 (.Y (nx138), .A0 (nx832), .A1 (CurRow_7)) ;
    or04 ix830 (.Y (nx829), .A0 (nx1042), .A1 (nx14), .A2 (nx138), .A3 (nx1028)
         ) ;
    nor02ii ix137 (.Y (nx1042), .A0 (CurRow_7), .A1 (nx832)) ;
    nor02ii ix103 (.Y (nx102), .A0 (nx844), .A1 (CurRow_5)) ;
    xor2 ix307 (.Y (nx497), .A0 (nx852), .A1 (nx850)) ;
    mux21_ni ix606 (.Y (nx605), .A0 (CurCol_1), .A1 (nx322), .S0 (nx1056)) ;
    and02 ix857 (.Y (nx856), .A0 (nx861), .A1 (nx858)) ;
    nor02ii ix331 (.Y (nx499), .A0 (nx858), .A1 (CurCol_1)) ;
    or03 ix449 (.Y (nx448), .A0 (CurCol_1), .A1 (FilterSize), .A2 (CurCol_0)) ;
    mux21_ni ix626 (.Y (nx625), .A0 (CurCol_3), .A1 (nx358), .S0 (nx1056)) ;
    and02 ix880 (.Y (nx879), .A0 (nx875), .A1 (nx870)) ;
    nor02ii ix367 (.Y (nx503), .A0 (nx870), .A1 (CurCol_3)) ;
    or02 ix911 (.Y (nx910), .A0 (FilterSize), .A1 (nx852)) ;
    oai222 ix914 (.Y (MemAddr[1]), .A0 (nx1060), .A1 (nx1044), .B0 (nx861), .B1 (
           nx1036), .C0 (nx787), .C1 (nx962)) ;
    inv01 ix1043 (.Y (nx1044), .A (nx500)) ;
    and02 ix473 (.Y (nx472), .A0 (nx1060), .A1 (CacheWindowWR)) ;
    xor2 ix918 (.Y (nx917), .A0 (FilterSize), .A1 (nx861)) ;
    nor02ii ix525 (.Y (nx524), .A0 (nx923), .A1 (CurCol_2)) ;
    nor02ii ix561 (.Y (nx560), .A0 (nx932), .A1 (CurCol_4)) ;
    xor2 ix613 (.Y (nx612), .A0 (nx596), .A1 (CurCol_7)) ;
    nor02ii ix597 (.Y (nx596), .A0 (nx946), .A1 (CurCol_6)) ;
    or02 ix629 (.Y (nx628), .A0 (nx1060), .A1 (FilterSize)) ;
    nor02ii ix965 (.Y (nx964), .A0 (FilterSize), .A1 (nx711)) ;
    oai22 ix651 (.Y (MemAddr[9]), .A0 (nx1060), .A1 (nx1046), .B0 (nx787), .B1 (
          nx1036)) ;
    inv01 ix1045 (.Y (nx1046), .A (nx646)) ;
    xor2 ix165 (.Y (nx164), .A0 (FilterSize), .A1 (nx787)) ;
    oai22 ix675 (.Y (MemAddr[10]), .A0 (nx1060), .A1 (nx1048), .B0 (nx775), .B1 (
          nx1036)) ;
    inv01 ix1047 (.Y (nx1048), .A (nx668)) ;
    nor02ii ix978 (.Y (nx977), .A0 (nx662), .A1 (nx764)) ;
    oai22 ix703 (.Y (MemAddr[12]), .A0 (nx1060), .A1 (nx1050), .B0 (nx758), .B1 (
          nx1036)) ;
    inv01 ix1049 (.Y (nx1050), .A (nx696)) ;
    nor02ii ix986 (.Y (nx985), .A0 (nx690), .A1 (nx842)) ;
    xor2 ix989 (.Y (nx988), .A0 (nx836), .A1 (nx985)) ;
    oai32 ix743 (.Y (MemAddr[15]), .A0 (nx1052), .A1 (Stride), .A2 (nx1062), .B0 (
          nx826), .B1 (nx1036)) ;
    xnor2 ix733 (.Y (nx1052), .A0 (nx826), .A1 (nx718)) ;
    inv02 ix1053 (.Y (nx1054), .A (nx1028)) ;
    inv02 ix1055 (.Y (nx1056), .A (nx1028)) ;
    inv02 ix1057 (.Y (nx1058), .A (MemWR)) ;
    inv02 ix1059 (.Y (nx1060), .A (MemWR)) ;
    inv02 ix1061 (.Y (nx1062), .A (MemWR)) ;
endmodule

