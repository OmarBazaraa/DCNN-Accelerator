//
// Verilog description for cell RAM, 
// Sat May 12 15:08:59 2018
//
// LeonardoSpectrum Level 3, 2017a.2 
//


module RAM ( CLK, WR, Address, Din, Dout ) ;

    input CLK ;
    input WR ;
    input [17:0]Address ;
    input [7:0]Din ;
    output [39:0]Dout ;

    wire Mem_2__0, nx2, nx14, nx22, nx28, nx32, nx44, nx60, nx64, nx74, nx80, 
         nx90, nx108, nx114, Mem_7__0, nx120, nx124, nx128, nx144, nx150, nx158, 
         nx166, nx180, nx184, nx188, nx198, nx204, nx212, nx224, nx228, Mem_3__0, 
         nx258, nx270, Mem_6__0, nx286, nx308, Mem_5__0, nx318, nx326, nx334, 
         nx346, nx354, nx366, nx376, Mem_1__0, nx404, nx416, Mem_0__0, nx422, 
         nx430, nx436, nx446, nx458, nx464, nx476, Mem_4__0, nx504, nx514, 
         Mem_2__1, Mem_7__1, Mem_3__1, Mem_6__1, Mem_5__1, Mem_1__1, Mem_0__1, 
         Mem_4__1, Mem_2__2, Mem_7__2, Mem_3__2, Mem_6__2, Mem_5__2, Mem_1__2, 
         Mem_0__2, Mem_4__2, Mem_2__3, Mem_7__3, Mem_3__3, Mem_6__3, Mem_5__3, 
         Mem_1__3, Mem_0__3, Mem_4__3, Mem_2__4, Mem_7__4, Mem_3__4, Mem_6__4, 
         Mem_5__4, Mem_1__4, Mem_0__4, Mem_4__4, Mem_2__5, Mem_7__5, Mem_3__5, 
         Mem_6__5, Mem_5__5, Mem_1__5, Mem_0__5, Mem_4__5, Mem_2__6, Mem_7__6, 
         Mem_3__6, Mem_6__6, Mem_5__6, Mem_1__6, Mem_0__6, Mem_4__6, Mem_2__7, 
         Mem_7__7, Mem_3__7, Mem_6__7, Mem_5__7, Mem_1__7, Mem_0__7, Mem_4__7, 
         nx1084, nx1092, nx1102, nx1108, Mem_8__0, nx1122, nx1130, nx1138, 
         nx1152, nx1162, nx1176, nx1188, nx1200, nx1210, Mem_8__1, Mem_8__2, 
         Mem_8__3, Mem_8__4, Mem_8__5, Mem_8__6, Mem_8__7, Mem_21__0, nx1472, 
         nx1480, nx1488, nx1502, nx1522, nx1534, nx1540, nx1546, nx1552, nx1558, 
         nx1572, Mem_22__0, nx1584, nx1594, nx1616, nx1626, Mem_20__0, nx1632, 
         nx1664, nx1674, nx1680, nx1692, nx1704, nx1718, nx1730, Mem_27__0, 
         nx1744, nx1756, nx1762, nx1770, nx1794, Mem_25__0, nx1824, nx1834, 
         Mem_26__0, nx1852, nx1872, Mem_11__0, nx1904, nx1916, Mem_30__0, nx1932, 
         nx1944, nx1950, nx1972, Mem_31__0, nx1988, nx2010, nx2018, Mem_29__0, 
         nx2046, nx2056, Mem_18__0, nx2066, nx2096, nx2114, nx2122, Mem_9__0, 
         nx2150, nx2160, Mem_15__0, nx2170, nx2180, nx2196, nx2204, nx2216, 
         nx2220, Mem_10__0, nx2236, nx2258, Mem_19__0, nx2288, nx2298, Mem_13__0, 
         nx2326, nx2336, Mem_12__0, nx2360, Mem_14__0, nx2396, nx2422, Mem_23__0, 
         nx2448, nx2458, Mem_16__0, nx2486, nx2496, Mem_28__0, nx2516, nx2538, 
         Mem_24__0, nx2554, nx2576, Mem_17__0, nx2604, nx2614, Mem_21__1, 
         Mem_22__1, Mem_20__1, nx2658, nx2664, nx2670, Mem_27__1, Mem_25__1, 
         Mem_26__1, Mem_11__1, Mem_30__1, Mem_31__1, nx2736, Mem_29__1, 
         Mem_18__1, Mem_9__1, Mem_15__1, Mem_10__1, Mem_19__1, Mem_13__1, 
         Mem_12__1, Mem_14__1, nx2828, Mem_23__1, Mem_16__1, Mem_28__1, 
         Mem_24__1, Mem_17__1, Mem_21__2, Mem_22__2, Mem_20__2, nx2914, nx2920, 
         nx2926, Mem_27__2, Mem_25__2, Mem_26__2, Mem_11__2, Mem_30__2, 
         Mem_31__2, nx2992, Mem_29__2, Mem_18__2, Mem_9__2, Mem_15__2, Mem_10__2, 
         Mem_19__2, Mem_13__2, Mem_12__2, Mem_14__2, nx3084, Mem_23__2, 
         Mem_16__2, Mem_28__2, Mem_24__2, Mem_17__2, Mem_21__3, Mem_22__3, 
         Mem_20__3, nx3170, nx3176, nx3182, Mem_27__3, Mem_25__3, Mem_26__3, 
         Mem_11__3, Mem_30__3, Mem_31__3, nx3248, Mem_29__3, Mem_18__3, Mem_9__3, 
         Mem_15__3, Mem_10__3, Mem_19__3, Mem_13__3, Mem_12__3, Mem_14__3, 
         nx3340, Mem_23__3, Mem_16__3, Mem_28__3, Mem_24__3, Mem_17__3, 
         Mem_21__4, Mem_22__4, Mem_20__4, nx3426, nx3432, nx3438, Mem_27__4, 
         Mem_25__4, Mem_26__4, Mem_11__4, Mem_30__4, Mem_31__4, nx3504, 
         Mem_29__4, Mem_18__4, Mem_9__4, Mem_15__4, Mem_10__4, Mem_19__4, 
         Mem_13__4, Mem_12__4, Mem_14__4, nx3596, Mem_23__4, Mem_16__4, 
         Mem_28__4, Mem_24__4, Mem_17__4, Mem_21__5, Mem_22__5, Mem_20__5, 
         nx3682, nx3688, nx3694, Mem_27__5, Mem_25__5, Mem_26__5, Mem_11__5, 
         Mem_30__5, Mem_31__5, nx3760, Mem_29__5, Mem_18__5, Mem_9__5, Mem_15__5, 
         Mem_10__5, Mem_19__5, Mem_13__5, Mem_12__5, Mem_14__5, nx3852, 
         Mem_23__5, Mem_16__5, Mem_28__5, Mem_24__5, Mem_17__5, Mem_21__6, 
         Mem_22__6, Mem_20__6, nx3938, nx3944, nx3950, Mem_27__6, Mem_25__6, 
         Mem_26__6, Mem_11__6, Mem_30__6, Mem_31__6, nx4016, Mem_29__6, 
         Mem_18__6, Mem_9__6, Mem_15__6, Mem_10__6, Mem_19__6, Mem_13__6, 
         Mem_12__6, Mem_14__6, nx4108, Mem_23__6, Mem_16__6, Mem_28__6, 
         Mem_24__6, Mem_17__6, Mem_21__7, Mem_22__7, Mem_20__7, nx4194, nx4200, 
         nx4206, Mem_27__7, Mem_25__7, Mem_26__7, Mem_11__7, Mem_30__7, 
         Mem_31__7, nx4272, Mem_29__7, Mem_18__7, Mem_9__7, Mem_15__7, Mem_10__7, 
         Mem_19__7, Mem_13__7, Mem_12__7, Mem_14__7, nx4364, Mem_23__7, 
         Mem_16__7, Mem_28__7, Mem_24__7, Mem_17__7, nx4420, nx4428, nx4430, 
         nx4436, nx4444, nx4454, nx4470, nx4476, nx4482, nx4490, nx4498, nx4504, 
         nx4514, nx4530, nx4534, nx4540, nx4544, nx4548, nx4554, nx4558, nx4566, 
         nx4576, nx4584, nx4586, nx4594, nx4606, nx4610, nx4616, nx4620, nx4628, 
         nx4632, nx4636, nx4646, nx4650, nx4664, nx4668, nx4672, nx4676, nx4694, 
         nx4700, nx4716, nx4744, nx4784, nx4808, nx4814, nx4830, nx4858, nx4898, 
         nx4922, nx4928, nx4944, nx4972, nx5012, nx5036, nx5042, nx5058, nx5086, 
         nx5126, nx5150, nx5156, nx5172, nx5200, nx5240, nx5264, nx5270, nx5286, 
         nx5314, nx5354, nx5378, nx5384, nx5400, nx5428, nx5468, nx5494, nx5496, 
         nx5502, nx5504, nx5510, nx5512, nx5522, nx5532, nx5538, nx5552, nx5562, 
         nx5566, nx5582, nx5592, nx5604, nx5608, nx5616, nx5620, nx5624, nx5640, 
         nx5650, nx5652, nx5656, nx5664, nx5668, nx5672, nx5690, nx5692, nx5696, 
         nx5704, nx5708, nx5712, nx5736, nx5784, nx5810, nx5846, nx5894, nx5920, 
         nx5956, nx6004, nx6030, nx6066, nx6114, nx6140, nx6176, nx6224, nx6250, 
         nx6286, nx6334, nx6360, nx6396, nx6444, nx6470, nx12614, nx12624, 
         nx12634, nx12644, nx12654, nx12664, nx12674, nx12684, nx12694, nx12704, 
         nx12714, nx12724, nx12734, nx12744, nx12754, nx12764, nx12774, nx12784, 
         nx12794, nx12804, nx12814, nx12824, nx12834, nx12844, nx12854, nx12864, 
         nx12874, nx12884, nx12894, nx12904, nx12914, nx12924, nx12934, nx12944, 
         nx12954, nx12964, nx12974, nx12984, nx12994, nx13004, nx13014, nx13024, 
         nx13034, nx13044, nx13054, nx13064, nx13074, nx13084, nx13094, nx13104, 
         nx13114, nx13124, nx13134, nx13144, nx13154, nx13164, nx13174, nx13184, 
         nx13194, nx13204, nx13214, nx13224, nx13234, nx13244, nx13254, nx13264, 
         nx13274, nx13284, nx13294, nx13304, nx13314, nx13324, nx13334, nx13344, 
         nx13354, nx13364, nx13374, nx13384, nx13394, nx13404, nx13414, nx13424, 
         nx13434, nx13444, nx13454, nx13464, nx13474, nx13484, nx13494, nx13504, 
         nx13514, nx13524, nx13534, nx13544, nx13554, nx13564, nx13574, nx13584, 
         nx13594, nx13604, nx13614, nx13624, nx13634, nx13644, nx13654, nx13664, 
         nx13674, nx13684, nx13694, nx13704, nx13714, nx13724, nx13734, nx13744, 
         nx13754, nx13764, nx13774, nx13784, nx13794, nx13804, nx13814, nx13824, 
         nx13834, nx13844, nx13854, nx13864, nx13874, nx13884, nx13894, nx13904, 
         nx13914, nx13924, nx13934, nx13944, nx13954, nx13964, nx13974, nx13984, 
         nx13994, nx14004, nx14014, nx14024, nx14034, nx14044, nx14054, nx14064, 
         nx14074, nx14084, nx14094, nx14104, nx14114, nx14124, nx14134, nx14144, 
         nx14154, nx14164, nx14174, nx14184, nx14194, nx14204, nx14214, nx14224, 
         nx14234, nx14244, nx14254, nx14264, nx14274, nx14284, nx14294, nx14304, 
         nx14314, nx14324, nx14334, nx14344, nx14354, nx14364, nx14374, nx14384, 
         nx14394, nx14404, nx14414, nx14424, nx14434, nx14444, nx14454, nx14464, 
         nx14474, nx14484, nx14494, nx14504, nx14514, nx14524, nx14534, nx14544, 
         nx14554, nx14564, nx14574, nx14584, nx14594, nx14604, nx14614, nx14624, 
         nx14634, nx14644, nx14654, nx14664, nx14674, nx14684, nx14694, nx14704, 
         nx14714, nx14724, nx14734, nx14744, nx14754, nx14764, nx14774, nx14784, 
         nx14794, nx14804, nx14814, nx14824, nx14834, nx14844, nx14854, nx14864, 
         nx14874, nx14884, nx14894, nx14904, nx14914, nx14924, nx14934, nx14944, 
         nx14954, nx14964, nx14974, nx14984, nx14994, nx15004, nx15014, nx15024, 
         nx15034, nx15044, nx15054, nx15064, nx15074, nx15084, nx15094, nx15104, 
         nx15114, nx15124, nx15134, nx15144, nx15154, nx15164, nx15175, nx15180, 
         nx15182, nx15184, nx15186, nx15188, nx15192, nx15196, nx15198, nx15200, 
         nx15203, nx15206, nx15208, nx15210, nx15214, nx15226, nx15230, nx15234, 
         nx15236, nx15240, nx15242, nx15244, nx15246, nx15255, nx15258, nx15260, 
         nx15262, nx15270, nx15272, nx15274, nx15281, nx15283, nx15286, nx15291, 
         nx15296, nx15301, nx15306, nx15308, nx15314, nx15316, nx15318, nx15320, 
         nx15322, nx15324, nx15326, nx15329, nx15334, nx15337, nx15341, nx15343, 
         nx15348, nx15350, nx15355, nx15362, nx15363, nx15370, nx15371, nx15375, 
         nx15378, nx15379, nx15383, nx15388, nx15395, nx15396, nx15403, nx15404, 
         nx15408, nx15411, nx15412, nx15416, nx15421, nx15428, nx15429, nx15436, 
         nx15437, nx15441, nx15444, nx15445, nx15449, nx15454, nx15461, nx15462, 
         nx15469, nx15470, nx15474, nx15477, nx15478, nx15482, nx15487, nx15494, 
         nx15495, nx15502, nx15503, nx15507, nx15510, nx15511, nx15515, nx15520, 
         nx15527, nx15528, nx15535, nx15536, nx15540, nx15543, nx15544, nx15548, 
         nx15553, nx15560, nx15561, nx15568, nx15569, nx15573, nx15576, nx15577, 
         nx15581, nx15586, nx15590, nx15596, nx15598, nx15600, nx15605, nx15609, 
         nx15614, nx15616, nx15621, nx15623, nx15626, nx15628, nx15633, nx15635, 
         nx15638, nx15640, nx15645, nx15647, nx15650, nx15652, nx15657, nx15659, 
         nx15662, nx15664, nx15669, nx15671, nx15674, nx15676, nx15681, nx15683, 
         nx15686, nx15688, nx15693, nx15695, nx15698, nx15702, nx15704, nx15708, 
         nx15711, nx15713, nx15715, nx15717, nx15720, nx15723, nx15727, nx15731, 
         nx15733, nx15736, nx15740, nx15744, nx15746, nx15754, nx15756, nx15758, 
         nx15765, nx15767, nx15769, nx15771, nx15774, nx15780, nx15782, nx15786, 
         nx15791, nx15793, nx15795, nx15798, nx15807, nx15811, nx15813, nx15817, 
         nx15819, nx15821, nx15824, nx15828, nx15833, nx15836, nx15838, nx15840, 
         nx15846, nx15848, nx15853, nx15855, nx15865, nx15869, nx15873, nx15875, 
         nx15877, nx15881, nx15887, nx15891, nx15895, nx15901, nx15907, nx15912, 
         nx15914, nx15916, nx15921, nx15923, nx15929, nx15932, nx15936, nx15939, 
         nx15942, nx15944, nx15946, nx15950, nx15953, nx15956, nx15963, nx15967, 
         nx15971, nx15979, nx15981, nx15985, nx15989, nx15991, nx15997, nx16000, 
         nx16003, nx16006, nx16008, nx16011, nx16013, nx16018, nx16020, nx16022, 
         nx16025, nx16031, nx16033, nx16038, nx16043, nx16047, nx16053, nx16054, 
         nx16058, nx16063, nx16067, nx16071, nx16073, nx16077, nx16081, nx16089, 
         nx16094, nx16098, nx16102, nx16105, nx16109, nx16116, nx16124, nx16132, 
         nx16136, nx16140, nx16145, nx16149, nx16155, nx16156, nx16160, nx16165, 
         nx16169, nx16173, nx16175, nx16179, nx16183, nx16191, nx16196, nx16200, 
         nx16204, nx16207, nx16211, nx16218, nx16226, nx16234, nx16238, nx16242, 
         nx16247, nx16251, nx16257, nx16258, nx16262, nx16267, nx16271, nx16275, 
         nx16277, nx16281, nx16285, nx16293, nx16298, nx16302, nx16306, nx16309, 
         nx16313, nx16320, nx16328, nx16336, nx16340, nx16344, nx16349, nx16353, 
         nx16359, nx16360, nx16364, nx16369, nx16373, nx16377, nx16379, nx16383, 
         nx16387, nx16395, nx16400, nx16404, nx16408, nx16411, nx16415, nx16422, 
         nx16430, nx16438, nx16442, nx16446, nx16451, nx16455, nx16461, nx16462, 
         nx16466, nx16471, nx16475, nx16479, nx16481, nx16485, nx16489, nx16497, 
         nx16502, nx16506, nx16510, nx16513, nx16517, nx16524, nx16532, nx16540, 
         nx16544, nx16548, nx16553, nx16557, nx16563, nx16564, nx16568, nx16573, 
         nx16577, nx16581, nx16583, nx16587, nx16591, nx16599, nx16604, nx16608, 
         nx16612, nx16615, nx16619, nx16626, nx16634, nx16642, nx16646, nx16650, 
         nx16655, nx16659, nx16665, nx16666, nx16670, nx16675, nx16679, nx16683, 
         nx16685, nx16689, nx16693, nx16701, nx16706, nx16710, nx16714, nx16717, 
         nx16721, nx16728, nx16736, nx16744, nx16748, nx16752, nx16757, nx16760, 
         nx16762, nx16764, nx16767, nx16770, nx16776, nx16778, nx16784, nx16786, 
         nx16794, nx16797, nx16800, nx16802, nx16805, nx16811, nx16817, nx16823, 
         nx16826, nx16833, nx16836, nx16839, nx16846, nx16848, nx16851, nx16856, 
         nx16858, nx16861, nx16863, nx16866, nx16868, nx16871, nx16873, nx16875, 
         nx16877, nx16879, nx16882, nx16884, nx16886, nx16889, nx16894, nx16896, 
         nx16899, nx16901, nx16903, nx16905, nx16907, nx16910, nx16912, nx16914, 
         nx16917, nx16922, nx16924, nx16927, nx16929, nx16931, nx16933, nx16935, 
         nx16938, nx16940, nx16942, nx16945, nx16950, nx16952, nx16955, nx16957, 
         nx16959, nx16961, nx16963, nx16966, nx16968, nx16970, nx16973, nx16978, 
         nx16980, nx16983, nx16985, nx16987, nx16989, nx16991, nx16994, nx16996, 
         nx16998, nx17001, nx17006, nx17008, nx17011, nx17013, nx17015, nx17017, 
         nx17019, nx17022, nx17024, nx17026, nx17029, nx17034, nx17036, nx17039, 
         nx17041, nx17043, nx17045, nx17047, nx17050, nx17052, nx17054, nx17057, 
         nx17062, nx17064, nx17067, nx17069, nx17072, nx17075, nx17078, nx17081, 
         nx17087, nx17093, nx17096, nx17103, nx17106, nx17109, nx17112, nx17115, 
         nx17118, nx17120, nx17126, nx17130, nx17134, nx17143, nx17149, nx17152, 
         nx17155, nx17157, nx17159, nx17162, nx17164, nx17167, nx17169, nx17171, 
         nx17173, nx17175, nx17177, nx17181, nx17183, nx17185, nx17188, nx17190, 
         nx17193, nx17195, nx17197, nx17199, nx17201, nx17203, nx17207, nx17209, 
         nx17211, nx17214, nx17216, nx17219, nx17221, nx17223, nx17225, nx17227, 
         nx17229, nx17233, nx17235, nx17237, nx17240, nx17242, nx17245, nx17247, 
         nx17249, nx17251, nx17253, nx17255, nx17259, nx17261, nx17263, nx17266, 
         nx17268, nx17271, nx17273, nx17275, nx17277, nx17279, nx17281, nx17285, 
         nx17287, nx17289, nx17292, nx17294, nx17297, nx17299, nx17301, nx17303, 
         nx17305, nx17307, nx17311, nx17313, nx17315, nx17318, nx17320, nx17323, 
         nx17325, nx17327, nx17329, nx17331, nx17333, nx17341, nx17343, nx17347, 
         nx17349, nx17351, nx17353, nx17355, nx17357, nx17359, nx17361, nx17363, 
         nx17365, nx17367, nx17369, nx17371, nx17373, nx17375, nx17377, nx17379, 
         nx17381, nx17383, nx17385, nx17387, nx17389, nx17391, nx17393, nx17395, 
         nx17397, nx17399, nx17401, nx17403, nx17405, nx17407, nx17409, nx17411, 
         nx17413, nx17415, nx17417, nx17419, nx17421, nx17423, nx17425, nx17427, 
         nx17429, nx17431, nx17433, nx17435, nx17437, nx17439, nx17441, nx17443, 
         nx17445, nx17447, nx17449, nx17451, nx17453, nx17455, nx17457, nx17459, 
         nx17461, nx17463, nx17465, nx17467, nx17469, nx17471, nx17473, nx17475, 
         nx17477, nx17479, nx17481, nx17483, nx17485, nx17487, nx17489, nx17491, 
         nx17493, nx17495, nx17497, nx17499, nx17501, nx17503, nx17505, nx17507, 
         nx17509, nx17511, nx17513, nx17515, nx17517, nx17519, nx17521, nx17523, 
         nx17525, nx17527, nx17529, nx17531, nx17533, nx17535, nx17537, nx17539, 
         nx17541, nx17543, nx17545, nx17547, nx17549, nx17551, nx17553, nx17555, 
         nx17557, nx17559, nx17561, nx17563, nx17565, nx17567, nx17569, nx17571, 
         nx17573, nx17575, nx17577, nx17579, nx17581, nx17583, nx17585, nx17587, 
         nx17589, nx17591, nx17593, nx17595, nx17597, nx17599, nx17601, nx17603, 
         nx17605, nx17607, nx17609, nx17611, nx17613, nx17615, nx17617, nx17619, 
         nx17621, nx17623, nx17625, nx17627, nx17629, nx17631, nx17633, nx17635, 
         nx17637, nx17641, nx17643, nx17645, nx17649, nx17651, nx17653, nx17655, 
         nx17665, nx17669, nx17671, nx17673, nx17675, nx17679, nx17681, nx17683, 
         nx17685, nx17687, nx17689, nx17691, nx17693, nx17695, nx17697, nx17699, 
         nx17701, nx17703, nx17705, nx17707, nx17709, nx17711, nx17713, nx17715, 
         nx17717, nx17719, nx17721, nx17723, nx17725, nx17727, nx17729, nx17731, 
         nx17733, nx17735, nx17737, nx17739, nx17741, nx17743, nx17745, nx17747, 
         nx17749, nx17751, nx17753, nx17755, nx17757, nx17759, nx17761, nx17763, 
         nx17765, nx17767, nx17769, nx17771, nx17773, nx17775, nx17779, nx17781, 
         nx17783, nx17787, nx17789, nx17791, nx17793, nx17795, nx17797, nx17799, 
         nx17801, nx17803, nx17805, nx17807, nx17809, nx17811, nx17813, nx17815, 
         nx17817, nx17821, nx17823, nx17825, nx17827, nx17829, nx17831, nx17833, 
         nx17835, nx17837, nx17839, nx17841, nx17843, nx17845, nx17847, nx17849, 
         nx17851, nx17853, nx18049, nx18051, nx18053, nx18055, nx18057, nx18059, 
         nx18061, nx18063, nx18065, nx18067, nx18069, nx18071, nx18073, nx18075, 
         nx18077, nx18079, nx18081, nx18083, nx18085, nx18087, nx18089, nx18091, 
         nx18093, nx18095, nx18097, nx18099, nx18101, nx18103, nx18105, nx18107, 
         nx18109, nx18111, nx18113, nx18115, nx18117, nx18119, nx18121, nx18123, 
         nx18125, nx18127, nx18129, nx18131, nx18133, nx18135, nx18137, nx18139, 
         nx18141, nx18143, nx18145, nx18147, nx18149, nx18151, nx18153, nx18155, 
         nx18157, nx18159, nx18161, nx18163, nx18165, nx18167;
    wire [135:0] \$dummy ;




    nand04 ix523 (.Y (Dout[0]), .A0 (nx15175), .A1 (nx15246), .A2 (nx15274), .A3 (
           nx15329)) ;
    aoi22 ix15176 (.Y (nx15175), .A0 (Mem_0__0), .A1 (nx476), .B0 (Mem_4__0), .B1 (
          nx514)) ;
    dff reg_Mem_0__0 (.Q (Mem_0__0), .QB (\$dummy [0]), .D (nx12674), .CLK (CLK)
        ) ;
    mux21_ni ix12675 (.Y (nx12674), .A0 (Mem_0__0), .A1 (Din[0]), .S0 (nx17363)
             ) ;
    oai321 ix465 (.Y (nx464), .A0 (Address[14]), .A1 (Address[13]), .A2 (nx15180
           ), .B0 (nx15186), .B1 (nx15192), .C0 (nx15198)) ;
    nand03 ix15181 (.Y (nx15180), .A0 (nx15182), .A1 (nx15184), .A2 (WR)) ;
    nor02_2x ix15183 (.Y (nx15182), .A0 (Address[15]), .A1 (Address[16])) ;
    inv02 ix15185 (.Y (nx15184), .A (Address[17])) ;
    inv01 ix15189 (.Y (nx15188), .A (Address[3])) ;
    nor02_2x ix15197 (.Y (nx15196), .A0 (Address[0]), .A1 (Address[1])) ;
    aoi222 ix15199 (.Y (nx15198), .A0 (nx15200), .A1 (nx17691), .B0 (nx15203), .B1 (
           nx14), .C0 (nx15210), .C1 (nx32)) ;
    nor02_2x ix15201 (.Y (nx15200), .A0 (Address[5]), .A1 (Address[4])) ;
    nor02_2x ix15204 (.Y (nx15203), .A0 (Address[2]), .A1 (Address[1])) ;
    nor03_2x ix15 (.Y (nx14), .A0 (nx15206), .A1 (Address[4]), .A2 (Address[3])
             ) ;
    nand02 ix15207 (.Y (nx15206), .A0 (nx15208), .A1 (WR)) ;
    inv02 ix15209 (.Y (nx15208), .A (Address[5])) ;
    nor02_2x ix15211 (.Y (nx15210), .A0 (Address[8]), .A1 (Address[9])) ;
    inv02 ix15215 (.Y (nx15214), .A (WR)) ;
    nor03_2x ix477 (.Y (nx476), .A0 (Address[17]), .A1 (Address[15]), .A2 (
             Address[16])) ;
    dff reg_Mem_4__0 (.Q (Mem_4__0), .QB (nx15244), .D (nx12684), .CLK (CLK)) ;
    nor02_2x ix15231 (.Y (nx15230), .A0 (Address[14]), .A1 (Address[13])) ;
    inv02 ix15235 (.Y (nx15234), .A (Address[16])) ;
    nand02 ix15237 (.Y (nx15236), .A0 (nx15184), .A1 (WR)) ;
    nor03_2x ix167 (.Y (nx166), .A0 (nx18129), .A1 (Address[12]), .A2 (nx15214)
             ) ;
    inv01 ix15241 (.Y (nx15240), .A (Address[11])) ;
    nor03_2x ix515 (.Y (nx514), .A0 (nx15184), .A1 (Address[15]), .A2 (
             Address[16])) ;
    aoi22 ix15247 (.Y (nx15246), .A0 (Mem_1__0), .A1 (nx17687), .B0 (Mem_5__0), 
          .B1 (nx376)) ;
    dff reg_Mem_1__0 (.Q (Mem_1__0), .QB (\$dummy [1]), .D (nx12664), .CLK (CLK)
        ) ;
    mux21_ni ix12665 (.Y (nx12664), .A0 (Mem_1__0), .A1 (Din[0]), .S0 (nx17359)
             ) ;
    oai321 ix405 (.Y (nx404), .A0 (nx15186), .A1 (Address[4]), .A2 (nx354), .B0 (
           nx318), .B1 (nx15180), .C0 (nx15255)) ;
    nand02 ix355 (.Y (nx354), .A0 (Address[0]), .A1 (nx17545)) ;
    nand02 ix319 (.Y (nx318), .A0 (nx17549), .A1 (Address[13])) ;
    aoi222 ix15256 (.Y (nx15255), .A0 (nx15200), .A1 (nx334), .B0 (nx15258), .B1 (
           nx14), .C0 (nx17815), .C1 (nx32)) ;
    inv01 ix15263 (.Y (nx15262), .A (Address[8])) ;
    dff reg_Mem_5__0 (.Q (Mem_5__0), .QB (nx15272), .D (nx12654), .CLK (CLK)) ;
    oai321 ix367 (.Y (nx366), .A0 (nx18131), .A1 (Address[4]), .A2 (nx354), .B0 (
           nx346), .B1 (nx15226), .C0 (nx15270)) ;
    nand02 ix347 (.Y (nx346), .A0 (nx17533), .A1 (Address[1])) ;
    aoi332 ix15271 (.Y (nx15270), .A0 (nx15208), .A1 (Address[4]), .A2 (nx334), 
           .B0 (nx17549), .B1 (Address[13]), .B2 (nx188), .C0 (nx17815), .C1 (
           nx166)) ;
    aoi22 ix15275 (.Y (nx15274), .A0 (Mem_3__0), .A1 (nx270), .B0 (Mem_6__0), .B1 (
          nx17683)) ;
    dff reg_Mem_3__0 (.Q (Mem_3__0), .QB (nx15291), .D (nx12634), .CLK (CLK)) ;
    oai221 ix259 (.Y (nx258), .A0 (nx180), .A1 (nx15180), .B0 (nx198), .B1 (
           nx15281), .C0 (nx15283)) ;
    nand02 ix181 (.Y (nx180), .A0 (Address[14]), .A1 (Address[13])) ;
    nand02 ix199 (.Y (nx198), .A0 (Address[2]), .A1 (Address[1])) ;
    aoi332 ix15284 (.Y (nx15283), .A0 (nx15208), .A1 (nx17537), .A2 (nx128), .B0 (
           Address[8]), .B1 (Address[9]), .B2 (nx32), .C0 (nx17341), .C1 (nx150)
           ) ;
    nand03 ix15287 (.Y (nx15286), .A0 (WR), .A1 (Address[3]), .A2 (Address[2])
           ) ;
    nor03_2x ix45 (.Y (nx44), .A0 (nx15214), .A1 (Address[3]), .A2 (Address[2])
             ) ;
    nor02_2x ix151 (.Y (nx150), .A0 (Address[4]), .A1 (nx144)) ;
    nand02 ix145 (.Y (nx144), .A0 (Address[0]), .A1 (Address[1])) ;
    nor02_2x ix271 (.Y (nx270), .A0 (Address[17]), .A1 (nx224)) ;
    nand02 ix225 (.Y (nx224), .A0 (Address[15]), .A1 (Address[16])) ;
    dff reg_Mem_6__0 (.Q (Mem_6__0), .QB (nx15326), .D (nx12644), .CLK (CLK)) ;
    aoi221 ix15297 (.Y (nx15296), .A0 (nx17813), .A1 (nx90), .B0 (nx15301), .B1 (
           nx204), .C0 (nx286)) ;
    nor03_2x ix205 (.Y (nx204), .A0 (nx15206), .A1 (Address[4]), .A2 (nx15188)
             ) ;
    oai222 ix287 (.Y (nx286), .A0 (nx22), .A1 (nx15306), .B0 (nx64), .B1 (
           nx15316), .C0 (nx18131), .C1 (nx15322)) ;
    nand02_2x ix23 (.Y (nx22), .A0 (nx15262), .A1 (Address[9])) ;
    inv01 ix15315 (.Y (nx15314), .A (Address[13])) ;
    nand03 ix15317 (.Y (nx15316), .A0 (nx15318), .A1 (nx15184), .A2 (WR)) ;
    inv02 ix15321 (.Y (nx15320), .A (Address[15])) ;
    nand02 ix15323 (.Y (nx15322), .A0 (nx17537), .A1 (nx17821)) ;
    nand02 ix109 (.Y (nx108), .A0 (nx15320), .A1 (Address[16])) ;
    aoi22 ix15330 (.Y (nx15329), .A0 (Mem_7__0), .A1 (nx17679), .B0 (Mem_2__0), 
          .B1 (nx114)) ;
    dff reg_Mem_7__0 (.Q (Mem_7__0), .QB (nx15337), .D (nx12624), .CLK (CLK)) ;
    oai221 ix213 (.Y (nx212), .A0 (nx198), .A1 (nx15226), .B0 (nx180), .B1 (
           nx15316), .C0 (nx15334)) ;
    aoi332 ix15335 (.Y (nx15334), .A0 (nx15208), .A1 (Address[4]), .A2 (nx128), 
           .B0 (Address[8]), .B1 (Address[9]), .B2 (nx166), .C0 (nx17675), .C1 (
           nx150)) ;
    dff reg_Mem_2__0 (.Q (Mem_2__0), .QB (\$dummy [2]), .D (nx12614), .CLK (CLK)
        ) ;
    mux21_ni ix12615 (.Y (nx12614), .A0 (Din[0]), .A1 (Mem_2__0), .S0 (nx17561)
             ) ;
    aoi221 ix15342 (.Y (nx15341), .A0 (nx15343), .A1 (nx74), .B0 (nx15200), .B1 (
           nx90), .C0 (nx60)) ;
    oai222 ix61 (.Y (nx60), .A0 (nx15186), .A1 (nx15322), .B0 (nx2), .B1 (
           nx15281), .C0 (nx22), .C1 (nx15348)) ;
    nand02 ix15349 (.Y (nx15348), .A0 (nx17823), .A1 (nx28)) ;
    nor02_2x ix15351 (.Y (nx15350), .A0 (Address[11]), .A1 (Address[10])) ;
    nor02_2x ix115 (.Y (nx114), .A0 (Address[17]), .A1 (nx108)) ;
    nand04 ix601 (.Y (Dout[1]), .A0 (nx15355), .A1 (nx15363), .A2 (nx15371), .A3 (
           nx15379)) ;
    aoi22 ix15356 (.Y (nx15355), .A0 (Mem_0__1), .A1 (nx476), .B0 (Mem_4__1), .B1 (
          nx514)) ;
    dff reg_Mem_0__1 (.Q (Mem_0__1), .QB (\$dummy [3]), .D (nx12754), .CLK (CLK)
        ) ;
    mux21_ni ix12755 (.Y (nx12754), .A0 (Mem_0__1), .A1 (Din[1]), .S0 (nx17363)
             ) ;
    dff reg_Mem_4__1 (.Q (Mem_4__1), .QB (nx15362), .D (nx12764), .CLK (CLK)) ;
    aoi22 ix15364 (.Y (nx15363), .A0 (Mem_1__1), .A1 (nx17687), .B0 (Mem_5__1), 
          .B1 (nx376)) ;
    dff reg_Mem_1__1 (.Q (Mem_1__1), .QB (\$dummy [4]), .D (nx12744), .CLK (CLK)
        ) ;
    mux21_ni ix12745 (.Y (nx12744), .A0 (Mem_1__1), .A1 (Din[1]), .S0 (nx17359)
             ) ;
    dff reg_Mem_5__1 (.Q (Mem_5__1), .QB (nx15370), .D (nx12734), .CLK (CLK)) ;
    aoi22 ix15372 (.Y (nx15371), .A0 (Mem_3__1), .A1 (nx270), .B0 (Mem_6__1), .B1 (
          nx17683)) ;
    dff reg_Mem_3__1 (.Q (Mem_3__1), .QB (nx15375), .D (nx12714), .CLK (CLK)) ;
    dff reg_Mem_6__1 (.Q (Mem_6__1), .QB (nx15378), .D (nx12724), .CLK (CLK)) ;
    aoi22 ix15380 (.Y (nx15379), .A0 (Mem_7__1), .A1 (nx17679), .B0 (Mem_2__1), 
          .B1 (nx114)) ;
    dff reg_Mem_7__1 (.Q (Mem_7__1), .QB (nx15383), .D (nx12704), .CLK (CLK)) ;
    dff reg_Mem_2__1 (.Q (Mem_2__1), .QB (\$dummy [5]), .D (nx12694), .CLK (CLK)
        ) ;
    mux21_ni ix12695 (.Y (nx12694), .A0 (Din[1]), .A1 (Mem_2__1), .S0 (nx17561)
             ) ;
    nand04 ix679 (.Y (Dout[2]), .A0 (nx15388), .A1 (nx15396), .A2 (nx15404), .A3 (
           nx15412)) ;
    aoi22 ix15389 (.Y (nx15388), .A0 (Mem_0__2), .A1 (nx476), .B0 (Mem_4__2), .B1 (
          nx514)) ;
    dff reg_Mem_0__2 (.Q (Mem_0__2), .QB (\$dummy [6]), .D (nx12834), .CLK (CLK)
        ) ;
    mux21_ni ix12835 (.Y (nx12834), .A0 (Mem_0__2), .A1 (Din[2]), .S0 (nx17363)
             ) ;
    dff reg_Mem_4__2 (.Q (Mem_4__2), .QB (nx15395), .D (nx12844), .CLK (CLK)) ;
    aoi22 ix15397 (.Y (nx15396), .A0 (Mem_1__2), .A1 (nx17687), .B0 (Mem_5__2), 
          .B1 (nx376)) ;
    dff reg_Mem_1__2 (.Q (Mem_1__2), .QB (\$dummy [7]), .D (nx12824), .CLK (CLK)
        ) ;
    mux21_ni ix12825 (.Y (nx12824), .A0 (Mem_1__2), .A1 (Din[2]), .S0 (nx17359)
             ) ;
    dff reg_Mem_5__2 (.Q (Mem_5__2), .QB (nx15403), .D (nx12814), .CLK (CLK)) ;
    aoi22 ix15405 (.Y (nx15404), .A0 (Mem_3__2), .A1 (nx270), .B0 (Mem_6__2), .B1 (
          nx17683)) ;
    dff reg_Mem_3__2 (.Q (Mem_3__2), .QB (nx15408), .D (nx12794), .CLK (CLK)) ;
    dff reg_Mem_6__2 (.Q (Mem_6__2), .QB (nx15411), .D (nx12804), .CLK (CLK)) ;
    aoi22 ix15413 (.Y (nx15412), .A0 (Mem_7__2), .A1 (nx17679), .B0 (Mem_2__2), 
          .B1 (nx114)) ;
    dff reg_Mem_7__2 (.Q (Mem_7__2), .QB (nx15416), .D (nx12784), .CLK (CLK)) ;
    dff reg_Mem_2__2 (.Q (Mem_2__2), .QB (\$dummy [8]), .D (nx12774), .CLK (CLK)
        ) ;
    mux21_ni ix12775 (.Y (nx12774), .A0 (Din[2]), .A1 (Mem_2__2), .S0 (nx17561)
             ) ;
    nand04 ix757 (.Y (Dout[3]), .A0 (nx15421), .A1 (nx15429), .A2 (nx15437), .A3 (
           nx15445)) ;
    aoi22 ix15422 (.Y (nx15421), .A0 (Mem_0__3), .A1 (nx476), .B0 (Mem_4__3), .B1 (
          nx514)) ;
    dff reg_Mem_0__3 (.Q (Mem_0__3), .QB (\$dummy [9]), .D (nx12914), .CLK (CLK)
        ) ;
    mux21_ni ix12915 (.Y (nx12914), .A0 (Mem_0__3), .A1 (Din[3]), .S0 (nx17363)
             ) ;
    dff reg_Mem_4__3 (.Q (Mem_4__3), .QB (nx15428), .D (nx12924), .CLK (CLK)) ;
    aoi22 ix15430 (.Y (nx15429), .A0 (Mem_1__3), .A1 (nx17687), .B0 (Mem_5__3), 
          .B1 (nx376)) ;
    dff reg_Mem_1__3 (.Q (Mem_1__3), .QB (\$dummy [10]), .D (nx12904), .CLK (CLK
        )) ;
    mux21_ni ix12905 (.Y (nx12904), .A0 (Mem_1__3), .A1 (Din[3]), .S0 (nx17359)
             ) ;
    dff reg_Mem_5__3 (.Q (Mem_5__3), .QB (nx15436), .D (nx12894), .CLK (CLK)) ;
    aoi22 ix15438 (.Y (nx15437), .A0 (Mem_3__3), .A1 (nx270), .B0 (Mem_6__3), .B1 (
          nx17683)) ;
    dff reg_Mem_3__3 (.Q (Mem_3__3), .QB (nx15441), .D (nx12874), .CLK (CLK)) ;
    dff reg_Mem_6__3 (.Q (Mem_6__3), .QB (nx15444), .D (nx12884), .CLK (CLK)) ;
    aoi22 ix15446 (.Y (nx15445), .A0 (Mem_7__3), .A1 (nx17679), .B0 (Mem_2__3), 
          .B1 (nx114)) ;
    dff reg_Mem_7__3 (.Q (Mem_7__3), .QB (nx15449), .D (nx12864), .CLK (CLK)) ;
    dff reg_Mem_2__3 (.Q (Mem_2__3), .QB (\$dummy [11]), .D (nx12854), .CLK (CLK
        )) ;
    mux21_ni ix12855 (.Y (nx12854), .A0 (Din[3]), .A1 (Mem_2__3), .S0 (nx17561)
             ) ;
    nand04 ix835 (.Y (Dout[4]), .A0 (nx15454), .A1 (nx15462), .A2 (nx15470), .A3 (
           nx15478)) ;
    aoi22 ix15455 (.Y (nx15454), .A0 (Mem_0__4), .A1 (nx476), .B0 (Mem_4__4), .B1 (
          nx514)) ;
    dff reg_Mem_0__4 (.Q (Mem_0__4), .QB (\$dummy [12]), .D (nx12994), .CLK (CLK
        )) ;
    mux21_ni ix12995 (.Y (nx12994), .A0 (Mem_0__4), .A1 (Din[4]), .S0 (nx17363)
             ) ;
    dff reg_Mem_4__4 (.Q (Mem_4__4), .QB (nx15461), .D (nx13004), .CLK (CLK)) ;
    aoi22 ix15463 (.Y (nx15462), .A0 (Mem_1__4), .A1 (nx17687), .B0 (Mem_5__4), 
          .B1 (nx376)) ;
    dff reg_Mem_1__4 (.Q (Mem_1__4), .QB (\$dummy [13]), .D (nx12984), .CLK (CLK
        )) ;
    mux21_ni ix12985 (.Y (nx12984), .A0 (Mem_1__4), .A1 (Din[4]), .S0 (nx17359)
             ) ;
    dff reg_Mem_5__4 (.Q (Mem_5__4), .QB (nx15469), .D (nx12974), .CLK (CLK)) ;
    aoi22 ix15471 (.Y (nx15470), .A0 (Mem_3__4), .A1 (nx270), .B0 (Mem_6__4), .B1 (
          nx17683)) ;
    dff reg_Mem_3__4 (.Q (Mem_3__4), .QB (nx15474), .D (nx12954), .CLK (CLK)) ;
    dff reg_Mem_6__4 (.Q (Mem_6__4), .QB (nx15477), .D (nx12964), .CLK (CLK)) ;
    aoi22 ix15479 (.Y (nx15478), .A0 (Mem_7__4), .A1 (nx17679), .B0 (Mem_2__4), 
          .B1 (nx114)) ;
    dff reg_Mem_7__4 (.Q (Mem_7__4), .QB (nx15482), .D (nx12944), .CLK (CLK)) ;
    dff reg_Mem_2__4 (.Q (Mem_2__4), .QB (\$dummy [14]), .D (nx12934), .CLK (CLK
        )) ;
    mux21_ni ix12935 (.Y (nx12934), .A0 (Din[4]), .A1 (Mem_2__4), .S0 (nx17561)
             ) ;
    nand04 ix913 (.Y (Dout[5]), .A0 (nx15487), .A1 (nx15495), .A2 (nx15503), .A3 (
           nx15511)) ;
    aoi22 ix15488 (.Y (nx15487), .A0 (Mem_0__5), .A1 (nx476), .B0 (Mem_4__5), .B1 (
          nx514)) ;
    dff reg_Mem_0__5 (.Q (Mem_0__5), .QB (\$dummy [15]), .D (nx13074), .CLK (CLK
        )) ;
    mux21_ni ix13075 (.Y (nx13074), .A0 (Mem_0__5), .A1 (Din[5]), .S0 (nx17363)
             ) ;
    dff reg_Mem_4__5 (.Q (Mem_4__5), .QB (nx15494), .D (nx13084), .CLK (CLK)) ;
    aoi22 ix15496 (.Y (nx15495), .A0 (Mem_1__5), .A1 (nx17687), .B0 (Mem_5__5), 
          .B1 (nx376)) ;
    dff reg_Mem_1__5 (.Q (Mem_1__5), .QB (\$dummy [16]), .D (nx13064), .CLK (CLK
        )) ;
    mux21_ni ix13065 (.Y (nx13064), .A0 (Mem_1__5), .A1 (Din[5]), .S0 (nx17359)
             ) ;
    dff reg_Mem_5__5 (.Q (Mem_5__5), .QB (nx15502), .D (nx13054), .CLK (CLK)) ;
    aoi22 ix15504 (.Y (nx15503), .A0 (Mem_3__5), .A1 (nx270), .B0 (Mem_6__5), .B1 (
          nx17683)) ;
    dff reg_Mem_3__5 (.Q (Mem_3__5), .QB (nx15507), .D (nx13034), .CLK (CLK)) ;
    dff reg_Mem_6__5 (.Q (Mem_6__5), .QB (nx15510), .D (nx13044), .CLK (CLK)) ;
    aoi22 ix15512 (.Y (nx15511), .A0 (Mem_7__5), .A1 (nx17679), .B0 (Mem_2__5), 
          .B1 (nx114)) ;
    dff reg_Mem_7__5 (.Q (Mem_7__5), .QB (nx15515), .D (nx13024), .CLK (CLK)) ;
    dff reg_Mem_2__5 (.Q (Mem_2__5), .QB (\$dummy [17]), .D (nx13014), .CLK (CLK
        )) ;
    mux21_ni ix13015 (.Y (nx13014), .A0 (Din[5]), .A1 (Mem_2__5), .S0 (nx17561)
             ) ;
    nand04 ix991 (.Y (Dout[6]), .A0 (nx15520), .A1 (nx15528), .A2 (nx15536), .A3 (
           nx15544)) ;
    aoi22 ix15521 (.Y (nx15520), .A0 (Mem_0__6), .A1 (nx476), .B0 (Mem_4__6), .B1 (
          nx514)) ;
    dff reg_Mem_0__6 (.Q (Mem_0__6), .QB (\$dummy [18]), .D (nx13154), .CLK (CLK
        )) ;
    mux21_ni ix13155 (.Y (nx13154), .A0 (Mem_0__6), .A1 (Din[6]), .S0 (nx17363)
             ) ;
    dff reg_Mem_4__6 (.Q (Mem_4__6), .QB (nx15527), .D (nx13164), .CLK (CLK)) ;
    aoi22 ix15529 (.Y (nx15528), .A0 (Mem_1__6), .A1 (nx17687), .B0 (Mem_5__6), 
          .B1 (nx376)) ;
    dff reg_Mem_1__6 (.Q (Mem_1__6), .QB (\$dummy [19]), .D (nx13144), .CLK (CLK
        )) ;
    mux21_ni ix13145 (.Y (nx13144), .A0 (Mem_1__6), .A1 (Din[6]), .S0 (nx17359)
             ) ;
    dff reg_Mem_5__6 (.Q (Mem_5__6), .QB (nx15535), .D (nx13134), .CLK (CLK)) ;
    aoi22 ix15537 (.Y (nx15536), .A0 (Mem_3__6), .A1 (nx270), .B0 (Mem_6__6), .B1 (
          nx17683)) ;
    dff reg_Mem_3__6 (.Q (Mem_3__6), .QB (nx15540), .D (nx13114), .CLK (CLK)) ;
    dff reg_Mem_6__6 (.Q (Mem_6__6), .QB (nx15543), .D (nx13124), .CLK (CLK)) ;
    aoi22 ix15545 (.Y (nx15544), .A0 (Mem_7__6), .A1 (nx17679), .B0 (Mem_2__6), 
          .B1 (nx114)) ;
    dff reg_Mem_7__6 (.Q (Mem_7__6), .QB (nx15548), .D (nx13104), .CLK (CLK)) ;
    dff reg_Mem_2__6 (.Q (Mem_2__6), .QB (\$dummy [20]), .D (nx13094), .CLK (CLK
        )) ;
    mux21_ni ix13095 (.Y (nx13094), .A0 (Din[6]), .A1 (Mem_2__6), .S0 (nx17561)
             ) ;
    nand04 ix1069 (.Y (Dout[7]), .A0 (nx15553), .A1 (nx15561), .A2 (nx15569), .A3 (
           nx15577)) ;
    aoi22 ix15554 (.Y (nx15553), .A0 (Mem_0__7), .A1 (nx476), .B0 (Mem_4__7), .B1 (
          nx514)) ;
    dff reg_Mem_0__7 (.Q (Mem_0__7), .QB (\$dummy [21]), .D (nx13234), .CLK (CLK
        )) ;
    mux21_ni ix13235 (.Y (nx13234), .A0 (Mem_0__7), .A1 (Din[7]), .S0 (nx17365)
             ) ;
    dff reg_Mem_4__7 (.Q (Mem_4__7), .QB (nx15560), .D (nx13244), .CLK (CLK)) ;
    aoi22 ix15562 (.Y (nx15561), .A0 (Mem_1__7), .A1 (nx17689), .B0 (Mem_5__7), 
          .B1 (nx376)) ;
    dff reg_Mem_1__7 (.Q (Mem_1__7), .QB (\$dummy [22]), .D (nx13224), .CLK (CLK
        )) ;
    mux21_ni ix13225 (.Y (nx13224), .A0 (Mem_1__7), .A1 (Din[7]), .S0 (nx17361)
             ) ;
    dff reg_Mem_5__7 (.Q (Mem_5__7), .QB (nx15568), .D (nx13214), .CLK (CLK)) ;
    aoi22 ix15570 (.Y (nx15569), .A0 (Mem_3__7), .A1 (nx270), .B0 (Mem_6__7), .B1 (
          nx17685)) ;
    dff reg_Mem_3__7 (.Q (Mem_3__7), .QB (nx15573), .D (nx13194), .CLK (CLK)) ;
    dff reg_Mem_6__7 (.Q (Mem_6__7), .QB (nx15576), .D (nx13204), .CLK (CLK)) ;
    aoi22 ix15578 (.Y (nx15577), .A0 (Mem_7__7), .A1 (nx17681), .B0 (Mem_2__7), 
          .B1 (nx114)) ;
    dff reg_Mem_7__7 (.Q (Mem_7__7), .QB (nx15581), .D (nx13184), .CLK (CLK)) ;
    dff reg_Mem_2__7 (.Q (Mem_2__7), .QB (\$dummy [23]), .D (nx13174), .CLK (CLK
        )) ;
    mux21_ni ix13175 (.Y (nx13174), .A0 (Din[7]), .A1 (Mem_2__7), .S0 (nx17563)
             ) ;
    nand04 ix1219 (.Y (Dout[8]), .A0 (nx15586), .A1 (nx15590), .A2 (nx15605), .A3 (
           nx15609)) ;
    aoi22 ix15587 (.Y (nx15586), .A0 (Mem_3__0), .A1 (nx1200), .B0 (Mem_5__0), .B1 (
          nx1210)) ;
    nor03_2x ix1201 (.Y (nx1200), .A0 (Address[16]), .A1 (Address[14]), .A2 (
             nx15320)) ;
    nor03_2x ix1211 (.Y (nx1210), .A0 (nx15234), .A1 (Address[14]), .A2 (
             Address[15])) ;
    aoi22 ix15591 (.Y (nx15590), .A0 (Mem_1__0), .A1 (nx1188), .B0 (Mem_8__0), .B1 (
          nx1176)) ;
    nor03_2x ix1189 (.Y (nx1188), .A0 (Address[16]), .A1 (Address[14]), .A2 (
             Address[15])) ;
    dff reg_Mem_8__0 (.Q (Mem_8__0), .QB (\$dummy [24]), .D (nx13254), .CLK (CLK
        )) ;
    mux21_ni ix13255 (.Y (nx13254), .A0 (Mem_8__0), .A1 (Din[0]), .S0 (nx17371)
             ) ;
    aoi332 ix15599 (.Y (nx15598), .A0 (nx15210), .A1 (nx17825), .A2 (nx28), .B0 (
           Address[5]), .B1 (nx17537), .B2 (nx17691), .C0 (nx15230), .C1 (nx1138
           )) ;
    nor02_2x ix1139 (.Y (nx1138), .A0 (nx108), .A1 (nx15236)) ;
    and03 ix1177 (.Y (nx1176), .A0 (Address[16]), .A1 (Address[14]), .A2 (
          Address[15])) ;
    aoi22 ix15606 (.Y (nx15605), .A0 (Mem_6__0), .A1 (nx1108), .B0 (Mem_7__0), .B1 (
          nx1102)) ;
    nor03_2x ix1109 (.Y (nx1108), .A0 (nx15234), .A1 (nx17549), .A2 (Address[15]
             )) ;
    nor03_2x ix1103 (.Y (nx1102), .A0 (nx15234), .A1 (Address[14]), .A2 (nx15320
             )) ;
    aoi22 ix15610 (.Y (nx15609), .A0 (Mem_2__0), .A1 (nx1092), .B0 (Mem_4__0), .B1 (
          nx1084)) ;
    nor03_2x ix1093 (.Y (nx1092), .A0 (Address[16]), .A1 (nx17549), .A2 (
             Address[15])) ;
    nor03_2x ix1085 (.Y (nx1084), .A0 (Address[16]), .A1 (nx17549), .A2 (nx15320
             )) ;
    nand04 ix1255 (.Y (Dout[9]), .A0 (nx15614), .A1 (nx15616), .A2 (nx15621), .A3 (
           nx15623)) ;
    aoi22 ix15615 (.Y (nx15614), .A0 (Mem_3__1), .A1 (nx1200), .B0 (Mem_5__1), .B1 (
          nx1210)) ;
    aoi22 ix15617 (.Y (nx15616), .A0 (Mem_1__1), .A1 (nx1188), .B0 (Mem_8__1), .B1 (
          nx1176)) ;
    dff reg_Mem_8__1 (.Q (Mem_8__1), .QB (\$dummy [25]), .D (nx13264), .CLK (CLK
        )) ;
    mux21_ni ix13265 (.Y (nx13264), .A0 (Mem_8__1), .A1 (Din[1]), .S0 (nx17371)
             ) ;
    aoi22 ix15622 (.Y (nx15621), .A0 (Mem_6__1), .A1 (nx1108), .B0 (Mem_7__1), .B1 (
          nx1102)) ;
    aoi22 ix15624 (.Y (nx15623), .A0 (Mem_2__1), .A1 (nx1092), .B0 (Mem_4__1), .B1 (
          nx1084)) ;
    nand04 ix1291 (.Y (Dout[10]), .A0 (nx15626), .A1 (nx15628), .A2 (nx15633), .A3 (
           nx15635)) ;
    aoi22 ix15627 (.Y (nx15626), .A0 (Mem_3__2), .A1 (nx1200), .B0 (Mem_5__2), .B1 (
          nx1210)) ;
    aoi22 ix15629 (.Y (nx15628), .A0 (Mem_1__2), .A1 (nx1188), .B0 (Mem_8__2), .B1 (
          nx1176)) ;
    dff reg_Mem_8__2 (.Q (Mem_8__2), .QB (\$dummy [26]), .D (nx13274), .CLK (CLK
        )) ;
    mux21_ni ix13275 (.Y (nx13274), .A0 (Mem_8__2), .A1 (Din[2]), .S0 (nx17371)
             ) ;
    aoi22 ix15634 (.Y (nx15633), .A0 (Mem_6__2), .A1 (nx1108), .B0 (Mem_7__2), .B1 (
          nx1102)) ;
    aoi22 ix15636 (.Y (nx15635), .A0 (Mem_2__2), .A1 (nx1092), .B0 (Mem_4__2), .B1 (
          nx1084)) ;
    nand04 ix1327 (.Y (Dout[11]), .A0 (nx15638), .A1 (nx15640), .A2 (nx15645), .A3 (
           nx15647)) ;
    aoi22 ix15639 (.Y (nx15638), .A0 (Mem_3__3), .A1 (nx1200), .B0 (Mem_5__3), .B1 (
          nx1210)) ;
    aoi22 ix15641 (.Y (nx15640), .A0 (Mem_1__3), .A1 (nx1188), .B0 (Mem_8__3), .B1 (
          nx1176)) ;
    dff reg_Mem_8__3 (.Q (Mem_8__3), .QB (\$dummy [27]), .D (nx13284), .CLK (CLK
        )) ;
    mux21_ni ix13285 (.Y (nx13284), .A0 (Mem_8__3), .A1 (Din[3]), .S0 (nx17371)
             ) ;
    aoi22 ix15646 (.Y (nx15645), .A0 (Mem_6__3), .A1 (nx1108), .B0 (Mem_7__3), .B1 (
          nx1102)) ;
    aoi22 ix15648 (.Y (nx15647), .A0 (Mem_2__3), .A1 (nx1092), .B0 (Mem_4__3), .B1 (
          nx1084)) ;
    nand04 ix1363 (.Y (Dout[12]), .A0 (nx15650), .A1 (nx15652), .A2 (nx15657), .A3 (
           nx15659)) ;
    aoi22 ix15651 (.Y (nx15650), .A0 (Mem_3__4), .A1 (nx1200), .B0 (Mem_5__4), .B1 (
          nx1210)) ;
    aoi22 ix15653 (.Y (nx15652), .A0 (Mem_1__4), .A1 (nx1188), .B0 (Mem_8__4), .B1 (
          nx1176)) ;
    dff reg_Mem_8__4 (.Q (Mem_8__4), .QB (\$dummy [28]), .D (nx13294), .CLK (CLK
        )) ;
    mux21_ni ix13295 (.Y (nx13294), .A0 (Mem_8__4), .A1 (Din[4]), .S0 (nx17371)
             ) ;
    aoi22 ix15658 (.Y (nx15657), .A0 (Mem_6__4), .A1 (nx1108), .B0 (Mem_7__4), .B1 (
          nx1102)) ;
    aoi22 ix15660 (.Y (nx15659), .A0 (Mem_2__4), .A1 (nx1092), .B0 (Mem_4__4), .B1 (
          nx1084)) ;
    nand04 ix1399 (.Y (Dout[13]), .A0 (nx15662), .A1 (nx15664), .A2 (nx15669), .A3 (
           nx15671)) ;
    aoi22 ix15663 (.Y (nx15662), .A0 (Mem_3__5), .A1 (nx1200), .B0 (Mem_5__5), .B1 (
          nx1210)) ;
    aoi22 ix15665 (.Y (nx15664), .A0 (Mem_1__5), .A1 (nx1188), .B0 (Mem_8__5), .B1 (
          nx1176)) ;
    dff reg_Mem_8__5 (.Q (Mem_8__5), .QB (\$dummy [29]), .D (nx13304), .CLK (CLK
        )) ;
    mux21_ni ix13305 (.Y (nx13304), .A0 (Mem_8__5), .A1 (Din[5]), .S0 (nx17371)
             ) ;
    aoi22 ix15670 (.Y (nx15669), .A0 (Mem_6__5), .A1 (nx1108), .B0 (Mem_7__5), .B1 (
          nx1102)) ;
    aoi22 ix15672 (.Y (nx15671), .A0 (Mem_2__5), .A1 (nx1092), .B0 (Mem_4__5), .B1 (
          nx1084)) ;
    nand04 ix1435 (.Y (Dout[14]), .A0 (nx15674), .A1 (nx15676), .A2 (nx15681), .A3 (
           nx15683)) ;
    aoi22 ix15675 (.Y (nx15674), .A0 (Mem_3__6), .A1 (nx1200), .B0 (Mem_5__6), .B1 (
          nx1210)) ;
    aoi22 ix15677 (.Y (nx15676), .A0 (Mem_1__6), .A1 (nx1188), .B0 (Mem_8__6), .B1 (
          nx1176)) ;
    dff reg_Mem_8__6 (.Q (Mem_8__6), .QB (\$dummy [30]), .D (nx13314), .CLK (CLK
        )) ;
    mux21_ni ix13315 (.Y (nx13314), .A0 (Mem_8__6), .A1 (Din[6]), .S0 (nx17371)
             ) ;
    aoi22 ix15682 (.Y (nx15681), .A0 (Mem_6__6), .A1 (nx1108), .B0 (Mem_7__6), .B1 (
          nx1102)) ;
    aoi22 ix15684 (.Y (nx15683), .A0 (Mem_2__6), .A1 (nx1092), .B0 (Mem_4__6), .B1 (
          nx1084)) ;
    nand04 ix1471 (.Y (Dout[15]), .A0 (nx15686), .A1 (nx15688), .A2 (nx15693), .A3 (
           nx15695)) ;
    aoi22 ix15687 (.Y (nx15686), .A0 (Mem_3__7), .A1 (nx1200), .B0 (Mem_5__7), .B1 (
          nx1210)) ;
    aoi22 ix15689 (.Y (nx15688), .A0 (Mem_1__7), .A1 (nx1188), .B0 (Mem_8__7), .B1 (
          nx1176)) ;
    dff reg_Mem_8__7 (.Q (Mem_8__7), .QB (\$dummy [31]), .D (nx13324), .CLK (CLK
        )) ;
    mux21_ni ix13325 (.Y (nx13324), .A0 (Mem_8__7), .A1 (Din[7]), .S0 (nx17373)
             ) ;
    aoi22 ix15694 (.Y (nx15693), .A0 (Mem_6__7), .A1 (nx1108), .B0 (Mem_7__7), .B1 (
          nx1102)) ;
    aoi22 ix15696 (.Y (nx15695), .A0 (Mem_2__7), .A1 (nx1092), .B0 (Mem_4__7), .B1 (
          nx1084)) ;
    nand04 ix2627 (.Y (Dout[16]), .A0 (nx15698), .A1 (nx15774), .A2 (nx15838), .A3 (
           nx15929)) ;
    aoi222 ix15699 (.Y (nx15698), .A0 (Mem_28__0), .A1 (nx17441), .B0 (Mem_24__0
           ), .B1 (nx17835), .C0 (Mem_17__0), .C1 (nx17837)) ;
    dff reg_Mem_28__0 (.Q (Mem_28__0), .QB (nx15717), .D (nx13534), .CLK (CLK)
        ) ;
    aoi321 ix15703 (.Y (nx15702), .A0 (nx15704), .A1 (Address[6]), .A2 (nx17341)
           , .B0 (nx15210), .B1 (nx1950), .C0 (nx2516)) ;
    nand02 ix1535 (.Y (nx1534), .A0 (Address[11]), .A1 (Address[10])) ;
    nand02 ix15709 (.Y (nx15708), .A0 (Address[12]), .A1 (WR)) ;
    oai222 ix2517 (.Y (nx2516), .A0 (nx17553), .A1 (nx15711), .B0 (nx422), .B1 (
           nx15713), .C0 (nx224), .C1 (nx15715)) ;
    nand02 ix15712 (.Y (nx15711), .A0 (Address[4]), .A1 (nx15196)) ;
    nand04 ix15714 (.Y (nx15713), .A0 (Address[5]), .A1 (WR), .A2 (Address[4]), 
           .A3 (Address[3])) ;
    nand03 ix15716 (.Y (nx15715), .A0 (nx15230), .A1 (Address[17]), .A2 (WR)) ;
    nand03 ix15721 (.Y (nx15720), .A0 (nx1540), .A1 (nx1546), .A2 (nx1552)) ;
    xnor2 ix1541 (.Y (nx1540), .A0 (Address[14]), .A1 (nx15723)) ;
    nand03 ix15724 (.Y (nx15723), .A0 (Address[13]), .A1 (Address[12]), .A2 (
           Address[11])) ;
    xnor2 ix1553 (.Y (nx1552), .A0 (Address[13]), .A1 (nx15727)) ;
    nand02 ix15728 (.Y (nx15727), .A0 (Address[12]), .A1 (Address[11])) ;
    dff reg_Mem_24__0 (.Q (Mem_24__0), .QB (\$dummy [32]), .D (nx13544), .CLK (
        CLK)) ;
    mux21_ni ix13545 (.Y (nx13544), .A0 (Din[0]), .A1 (Mem_24__0), .S0 (nx17569)
             ) ;
    aoi321 ix15732 (.Y (nx15731), .A0 (nx15733), .A1 (Address[6]), .A2 (nx17341)
           , .B0 (nx15203), .B1 (nx1762), .C0 (nx2554)) ;
    nor03_2x ix1763 (.Y (nx1762), .A0 (nx15736), .A1 (nx17537), .A2 (Address[3])
             ) ;
    nand02 ix15737 (.Y (nx15736), .A0 (Address[5]), .A1 (WR)) ;
    oai222 ix2555 (.Y (nx2554), .A0 (nx436), .A1 (nx15740), .B0 (nx18133), .B1 (
           nx15711), .C0 (nx108), .C1 (nx15715)) ;
    nand03 ix15741 (.Y (nx15740), .A0 (nx17825), .A1 (Address[12]), .A2 (WR)) ;
    nand03 ix15745 (.Y (nx15744), .A0 (nx1540), .A1 (nx17573), .A2 (nx1552)) ;
    oai21 ix15747 (.Y (nx15746), .A0 (Address[11]), .A1 (Address[12]), .B0 (
          nx15727)) ;
    dff reg_Mem_17__0 (.Q (Mem_17__0), .QB (nx15767), .D (nx13554), .CLK (CLK)
        ) ;
    oai221 ix2605 (.Y (nx2604), .A0 (nx326), .A1 (nx15754), .B0 (nx346), .B1 (
           nx15756), .C0 (nx15758)) ;
    nand03 ix15755 (.Y (nx15754), .A0 (nx17823), .A1 (Address[12]), .A2 (WR)) ;
    aoi222 ix15759 (.Y (nx15758), .A0 (nx17341), .A1 (nx17693), .B0 (nx15200), .B1 (
           nx1472), .C0 (nx15182), .C1 (nx1502)) ;
    nor02_2x ix1503 (.Y (nx1502), .A0 (nx318), .A1 (nx15765)) ;
    nand02 ix15766 (.Y (nx15765), .A0 (Address[17]), .A1 (WR)) ;
    nand03 ix15770 (.Y (nx15769), .A0 (nx1540), .A1 (nx17573), .A2 (nx15771)) ;
    aoi221 ix15775 (.Y (nx15774), .A0 (Mem_16__0), .A1 (nx17737), .B0 (Mem_23__0
           ), .B1 (nx17733), .C0 (nx2422)) ;
    dff reg_Mem_16__0 (.Q (Mem_16__0), .QB (nx15786), .D (nx13524), .CLK (CLK)
        ) ;
    oai221 ix2487 (.Y (nx2486), .A0 (nx80), .A1 (nx15780), .B0 (nx436), .B1 (
           nx15754), .C0 (nx15782)) ;
    nand02 ix15781 (.Y (nx15780), .A0 (Address[6]), .A1 (nx17341)) ;
    aoi322 ix15783 (.Y (nx15782), .A0 (nx17341), .A1 (Address[4]), .A2 (nx15196)
           , .B0 (nx15182), .B1 (nx1632), .C0 (nx15203), .C1 (nx2066)) ;
    nor03_2x ix2067 (.Y (nx2066), .A0 (nx15736), .A1 (Address[4]), .A2 (
             Address[3])) ;
    dff reg_Mem_23__0 (.Q (Mem_23__0), .QB (\$dummy [33]), .D (nx13514), .CLK (
        CLK)) ;
    mux21_ni ix13515 (.Y (nx13514), .A0 (Mem_23__0), .A1 (Din[0]), .S0 (nx17433)
             ) ;
    oai221 ix2449 (.Y (nx2448), .A0 (nx184), .A1 (nx15791), .B0 (nx198), .B1 (
           nx15793), .C0 (nx15795)) ;
    nand04 ix15794 (.Y (nx15793), .A0 (Address[5]), .A1 (WR), .A2 (nx17537), .A3 (
           Address[3])) ;
    aoi332 ix15796 (.Y (nx15795), .A0 (nx17813), .A1 (Address[6]), .A2 (nx17673)
           , .B0 (Address[8]), .B1 (Address[9]), .B2 (nx17695), .C0 (nx17675), .C1 (
           nx1744)) ;
    nand02 ix15799 (.Y (nx15798), .A0 (Address[3]), .A1 (Address[2])) ;
    oai22 ix2423 (.Y (nx2422), .A0 (nx15807), .A1 (nx15821), .B0 (nx15824), .B1 (
          nx17583)) ;
    dff reg_Mem_14__0 (.Q (Mem_14__0), .QB (nx15807), .D (nx13504), .CLK (CLK)
        ) ;
    aoi221 ix15812 (.Y (nx15811), .A0 (nx15704), .A1 (nx90), .B0 (nx15813), .B1 (
           nx2196), .C0 (nx2396)) ;
    nor03_2x ix2197 (.Y (nx2196), .A0 (nx17379), .A1 (Address[12]), .A2 (nx15214
             )) ;
    oai222 ix2397 (.Y (nx2396), .A0 (nx17553), .A1 (nx15322), .B0 (nx64), .B1 (
           nx15817), .C0 (nx2), .C1 (nx15819)) ;
    nand04 ix15820 (.Y (nx15819), .A0 (nx15208), .A1 (WR), .A2 (Address[4]), .A3 (
           Address[3])) ;
    nand02 ix15822 (.Y (nx15821), .A0 (nx17823), .A1 (nx2216)) ;
    nor03_2x ix2217 (.Y (nx2216), .A0 (nx1540), .A1 (nx17573), .A2 (nx15771)) ;
    dff reg_Mem_12__0 (.Q (Mem_12__0), .QB (nx15824), .D (nx13494), .CLK (CLK)
        ) ;
    aoi221 ix15829 (.Y (nx15828), .A0 (nx17673), .A1 (nx458), .B0 (nx15210), .B1 (
           nx2196), .C0 (nx2360)) ;
    nor03_2x ix459 (.Y (nx458), .A0 (Address[4]), .A1 (Address[0]), .A2 (
             Address[1])) ;
    oai222 ix2361 (.Y (nx2360), .A0 (nx1932), .A1 (nx15833), .B0 (nx446), .B1 (
           nx15817), .C0 (nx422), .C1 (nx15819)) ;
    nand02_2x ix1933 (.Y (nx1932), .A0 (Address[5]), .A1 (Address[4])) ;
    nand02 ix15837 (.Y (nx15836), .A0 (nx17825), .A1 (nx2216)) ;
    and04 ix15839 (.Y (nx15838), .A0 (nx15840), .A1 (nx15865), .A2 (nx15895), .A3 (
          nx15907)) ;
    aoi22 ix15841 (.Y (nx15840), .A0 (Mem_19__0), .A1 (nx17729), .B0 (Mem_13__0)
          , .B1 (nx2336)) ;
    dff reg_Mem_19__0 (.Q (Mem_19__0), .QB (nx15848), .D (nx13474), .CLK (CLK)
        ) ;
    oai321 ix2289 (.Y (nx2288), .A0 (Address[15]), .A1 (Address[16]), .A2 (
           nx15791), .B0 (nx158), .B1 (nx15754), .C0 (nx15846)) ;
    nand02 ix159 (.Y (nx158), .A0 (Address[8]), .A1 (Address[9])) ;
    aoi332 ix15847 (.Y (nx15846), .A0 (nx15200), .A1 (Address[6]), .A2 (nx17673)
           , .B0 (Address[2]), .B1 (Address[1]), .B2 (nx2066), .C0 (nx17341), .C1 (
           nx1744)) ;
    dff reg_Mem_13__0 (.Q (Mem_13__0), .QB (\$dummy [34]), .D (nx13484), .CLK (
        CLK)) ;
    mux21_ni ix13485 (.Y (nx13484), .A0 (Mem_13__0), .A1 (Din[0]), .S0 (nx17429)
             ) ;
    oai321 ix2327 (.Y (nx2326), .A0 (nx1932), .A1 (Address[6]), .A2 (nx18131), .B0 (
           nx17553), .B1 (nx15853), .C0 (nx15855)) ;
    nand03 ix15854 (.Y (nx15853), .A0 (nx17539), .A1 (Address[0]), .A2 (nx17545)
           ) ;
    aoi322 ix15856 (.Y (nx15855), .A0 (nx17549), .A1 (Address[13]), .A2 (nx2180)
           , .B0 (nx15258), .B1 (nx2170), .C0 (nx17815), .C1 (nx2196)) ;
    nor02_2x ix2181 (.Y (nx2180), .A0 (nx224), .A1 (nx15236)) ;
    aoi22 ix15866 (.Y (nx15865), .A0 (Mem_10__0), .A1 (nx17725), .B0 (Mem_15__0)
          , .B1 (nx2220)) ;
    dff reg_Mem_10__0 (.Q (Mem_10__0), .QB (\$dummy [35]), .D (nx13464), .CLK (
        CLK)) ;
    mux21_ni ix13465 (.Y (nx13464), .A0 (Din[0]), .A1 (Mem_10__0), .S0 (nx17587)
             ) ;
    aoi221 ix15870 (.Y (nx15869), .A0 (nx15733), .A1 (nx90), .B0 (nx15301), .B1 (
           nx1152), .C0 (nx2236)) ;
    nor03_2x ix1153 (.Y (nx1152), .A0 (nx15206), .A1 (nx17539), .A2 (Address[3])
             ) ;
    oai222 ix2237 (.Y (nx2236), .A0 (nx18133), .A1 (nx15322), .B0 (nx22), .B1 (
           nx15873), .C0 (nx64), .C1 (nx15875)) ;
    nand02 ix15874 (.Y (nx15873), .A0 (nx17825), .A1 (nx28)) ;
    nand02 ix15882 (.Y (nx15881), .A0 (nx1552), .A1 (nx1692)) ;
    dff reg_Mem_15__0 (.Q (Mem_15__0), .QB (\$dummy [36]), .D (nx13454), .CLK (
        CLK)) ;
    mux21_ni ix13455 (.Y (nx13454), .A0 (Mem_15__0), .A1 (Din[0]), .S0 (nx17421)
             ) ;
    oai321 ix2205 (.Y (nx2204), .A0 (nx1932), .A1 (Address[6]), .A2 (nx17553), .B0 (
           nx158), .B1 (nx15887), .C0 (nx15891)) ;
    aoi332 ix15892 (.Y (nx15891), .A0 (Address[14]), .A1 (Address[13]), .A2 (
           nx2180), .B0 (Address[2]), .B1 (Address[1]), .B2 (nx2170), .C0 (
           nx17673), .C1 (nx150)) ;
    aoi22 ix15896 (.Y (nx15895), .A0 (Mem_9__0), .A1 (nx17721), .B0 (Mem_8__0), 
          .B1 (nx17717)) ;
    dff reg_Mem_9__0 (.Q (Mem_9__0), .QB (\$dummy [37]), .D (nx13444), .CLK (CLK
        )) ;
    mux21_ni ix13445 (.Y (nx13444), .A0 (Mem_9__0), .A1 (Din[0]), .S0 (nx17417)
             ) ;
    oai321 ix2151 (.Y (nx2150), .A0 (nx1130), .A1 (Address[6]), .A2 (nx18131), .B0 (
           nx18133), .B1 (nx15853), .C0 (nx15901)) ;
    nand02 ix1131 (.Y (nx1130), .A0 (Address[5]), .A1 (nx17539)) ;
    aoi332 ix15902 (.Y (nx15901), .A0 (nx17551), .A1 (Address[13]), .A2 (nx1138)
           , .B0 (nx17533), .B1 (Address[1]), .B2 (nx1152), .C0 (nx17815), .C1 (
           nx1122)) ;
    aoi22 ix15908 (.Y (nx15907), .A0 (Mem_29__0), .A1 (nx17709), .B0 (Mem_18__0)
          , .B1 (nx17713)) ;
    dff reg_Mem_29__0 (.Q (Mem_29__0), .QB (nx15916), .D (nx13424), .CLK (CLK)
        ) ;
    oai221 ix2047 (.Y (nx2046), .A0 (nx326), .A1 (nx15912), .B0 (nx346), .B1 (
           nx15713), .C0 (nx15914)) ;
    aoi332 ix15915 (.Y (nx15914), .A0 (Address[15]), .A1 (Address[16]), .A2 (
           nx1502), .B0 (Address[5]), .B1 (Address[4]), .B2 (nx1472), .C0 (
           nx17673), .C1 (nx17693)) ;
    dff reg_Mem_18__0 (.Q (Mem_18__0), .QB (\$dummy [38]), .D (nx13434), .CLK (
        CLK)) ;
    mux21_ni ix13435 (.Y (nx13434), .A0 (Mem_18__0), .A1 (Din[0]), .S0 (nx17413)
             ) ;
    oai221 ix2097 (.Y (nx2096), .A0 (nx15186), .A1 (nx15921), .B0 (nx22), .B1 (
           nx15754), .C0 (nx15923)) ;
    nand02 ix15922 (.Y (nx15921), .A0 (Address[4]), .A1 (nx17821)) ;
    aoi222 ix15924 (.Y (nx15923), .A0 (nx15182), .A1 (nx1584), .B0 (nx15200), .B1 (
           nx1594), .C0 (nx15301), .C1 (nx2066)) ;
    nor04 ix15930 (.Y (nx15929), .A0 (nx2018), .A1 (nx1718), .A2 (nx1704), .A3 (
          nx1680)) ;
    nand03 ix2019 (.Y (nx2018), .A0 (nx15932), .A1 (nx15967), .A2 (nx15985)) ;
    aoi222 ix15933 (.Y (nx15932), .A0 (Mem_31__0), .A1 (nx17405), .B0 (Mem_30__0
           ), .B1 (nx17833), .C0 (Mem_11__0), .C1 (nx17831)) ;
    dff reg_Mem_31__0 (.Q (Mem_31__0), .QB (nx15946), .D (nx13414), .CLK (CLK)
        ) ;
    aoi321 ix15937 (.Y (nx15936), .A0 (Address[15]), .A1 (Address[16]), .A2 (
           nx1770), .B0 (nx15939), .B1 (nx1950), .C0 (nx1988)) ;
    nor02_2x ix1771 (.Y (nx1770), .A0 (nx180), .A1 (nx15765)) ;
    oai222 ix1989 (.Y (nx1988), .A0 (nx1932), .A1 (nx15942), .B0 (nx198), .B1 (
           nx15713), .C0 (nx17553), .C1 (nx15944)) ;
    nand02 ix15943 (.Y (nx15942), .A0 (Address[6]), .A1 (nx17673)) ;
    nand03 ix15945 (.Y (nx15944), .A0 (Address[4]), .A1 (Address[0]), .A2 (
           Address[1])) ;
    dff reg_Mem_30__0 (.Q (Mem_30__0), .QB (\$dummy [39]), .D (nx13404), .CLK (
        CLK)) ;
    mux21_ni ix13405 (.Y (nx13404), .A0 (Din[0]), .A1 (Mem_30__0), .S0 (nx17595)
             ) ;
    aoi321 ix15951 (.Y (nx15950), .A0 (nx124), .A1 (Address[4]), .A2 (nx17821), 
           .B0 (nx15813), .B1 (nx1950), .C0 (nx1944)) ;
    oai222 ix1945 (.Y (nx1944), .A0 (nx1932), .A1 (nx15953), .B0 (nx224), .B1 (
           nx15956), .C0 (nx2), .C1 (nx15713)) ;
    nand03 ix15957 (.Y (nx15956), .A0 (nx15343), .A1 (Address[17]), .A2 (WR)) ;
    dff reg_Mem_11__0 (.Q (Mem_11__0), .QB (\$dummy [40]), .D (nx13394), .CLK (
        CLK)) ;
    mux21_ni ix13395 (.Y (nx13394), .A0 (Mem_11__0), .A1 (Din[0]), .S0 (nx17397)
             ) ;
    oai321 ix1905 (.Y (nx1904), .A0 (nx1130), .A1 (Address[6]), .A2 (nx17553), .B0 (
           nx198), .B1 (nx15596), .C0 (nx15963)) ;
    aoi332 ix15964 (.Y (nx15963), .A0 (Address[14]), .A1 (Address[13]), .A2 (
           nx1138), .B0 (Address[8]), .B1 (Address[9]), .B2 (nx1122), .C0 (
           nx17671), .C1 (nx150)) ;
    aoi22 ix15968 (.Y (nx15967), .A0 (Mem_26__0), .A1 (nx17705), .B0 (Mem_25__0)
          , .B1 (nx17701)) ;
    dff reg_Mem_26__0 (.Q (Mem_26__0), .QB (\$dummy [41]), .D (nx13384), .CLK (
        CLK)) ;
    mux21_ni ix13385 (.Y (nx13384), .A0 (Din[0]), .A1 (Mem_26__0), .S0 (nx17599)
             ) ;
    aoi321 ix15972 (.Y (nx15971), .A0 (nx17671), .A1 (Address[4]), .A2 (nx17821)
           , .B0 (nx15301), .B1 (nx1762), .C0 (nx1852)) ;
    oai222 ix1853 (.Y (nx1852), .A0 (nx1130), .A1 (nx15953), .B0 (nx108), .B1 (
           nx15956), .C0 (nx22), .C1 (nx15740)) ;
    dff reg_Mem_25__0 (.Q (Mem_25__0), .QB (\$dummy [42]), .D (nx13374), .CLK (
        CLK)) ;
    mux21_ni ix13375 (.Y (nx13374), .A0 (Mem_25__0), .A1 (Din[0]), .S0 (nx17393)
             ) ;
    oai221 ix1825 (.Y (nx1824), .A0 (nx346), .A1 (nx15979), .B0 (nx326), .B1 (
           nx15740), .C0 (nx15981)) ;
    aoi332 ix15982 (.Y (nx15981), .A0 (nx15320), .A1 (Address[16]), .A2 (nx1502)
           , .B0 (Address[5]), .B1 (nx17539), .B2 (nx1472), .C0 (nx17671), .C1 (
           nx17693)) ;
    aoi22 ix15986 (.Y (nx15985), .A0 (Mem_27__0), .A1 (nx17697), .B0 (Mem_2__0)
          , .B1 (nx17389)) ;
    dff reg_Mem_27__0 (.Q (Mem_27__0), .QB (\$dummy [43]), .D (nx13364), .CLK (
        CLK)) ;
    mux21_ni ix13365 (.Y (nx13364), .A0 (Din[0]), .A1 (Mem_27__0), .S0 (nx17603)
             ) ;
    aoi221 ix15990 (.Y (nx15989), .A0 (nx15877), .A1 (nx1770), .B0 (nx15991), .B1 (
           nx1762), .C0 (nx1756)) ;
    oai222 ix1757 (.Y (nx1756), .A0 (nx1130), .A1 (nx15942), .B0 (nx18133), .B1 (
           nx15944), .C0 (nx158), .C1 (nx15740)) ;
    nor04 ix1731 (.Y (nx1730), .A0 (nx15997), .A1 (Address[11]), .A2 (
          Address[10]), .A3 (Address[13])) ;
    oai22 ix1719 (.Y (nx1718), .A0 (nx15337), .A1 (nx16000), .B0 (nx15272), .B1 (
          nx17607)) ;
    nand02 ix16001 (.Y (nx16000), .A0 (nx17817), .A1 (nx1572)) ;
    nor03_2x ix1573 (.Y (nx1572), .A0 (nx1540), .A1 (nx17573), .A2 (nx1552)) ;
    nand02 ix16004 (.Y (nx16003), .A0 (nx17829), .A1 (nx1572)) ;
    oai22 ix1705 (.Y (nx1704), .A0 (nx15244), .A1 (nx16006), .B0 (nx15291), .B1 (
          nx16008)) ;
    nand02 ix16007 (.Y (nx16006), .A0 (nx17825), .A1 (nx1572)) ;
    nand04 ix16009 (.Y (nx16008), .A0 (nx1692), .A1 (nx15240), .A2 (Address[10])
           , .A3 (nx15314)) ;
    oai221 ix1681 (.Y (nx1680), .A0 (nx15326), .A1 (nx17611), .B0 (nx16013), .B1 (
           nx17613), .C0 (nx16025)) ;
    nand02 ix16012 (.Y (nx16011), .A0 (nx17823), .A1 (nx1572)) ;
    dff reg_Mem_21__0 (.Q (Mem_21__0), .QB (nx16013), .D (nx13334), .CLK (CLK)
        ) ;
    oai221 ix1523 (.Y (nx1522), .A0 (nx346), .A1 (nx15793), .B0 (nx184), .B1 (
           nx16018), .C0 (nx16020)) ;
    aoi222 ix16021 (.Y (nx16020), .A0 (nx17815), .A1 (nx17695), .B0 (nx17675), .B1 (
           nx17693), .C0 (nx17813), .C1 (nx1472)) ;
    nand02 ix16023 (.Y (nx16022), .A0 (nx17829), .A1 (nx1558)) ;
    aoi22 ix16026 (.Y (nx16025), .A0 (Mem_20__0), .A1 (nx1674), .B0 (Mem_22__0)
          , .B1 (nx1626)) ;
    dff reg_Mem_20__0 (.Q (Mem_20__0), .QB (nx16033), .D (nx13354), .CLK (CLK)
        ) ;
    oai221 ix1665 (.Y (nx1664), .A0 (nx120), .A1 (nx15780), .B0 (nx422), .B1 (
           nx15793), .C0 (nx16031)) ;
    aoi332 ix16032 (.Y (nx16031), .A0 (nx17675), .A1 (Address[4]), .A2 (nx15196)
           , .B0 (Address[15]), .B1 (nx15234), .B2 (nx1632), .C0 (nx15210), .C1 (
           nx17695)) ;
    and02 ix1675 (.Y (nx1674), .A0 (nx17825), .A1 (nx1558)) ;
    dff reg_Mem_22__0 (.Q (Mem_22__0), .QB (\$dummy [44]), .D (nx13344), .CLK (
        CLK)) ;
    mux21_ni ix13345 (.Y (nx13344), .A0 (Mem_22__0), .A1 (Din[0]), .S0 (nx17381)
             ) ;
    oai221 ix1617 (.Y (nx1616), .A0 (nx17543), .A1 (nx15921), .B0 (nx2), .B1 (
           nx15793), .C0 (nx16038)) ;
    aoi222 ix16039 (.Y (nx16038), .A0 (nx15813), .A1 (nx17695), .B0 (nx17813), .B1 (
           nx1594), .C0 (nx15318), .C1 (nx1584)) ;
    and02 ix1627 (.Y (nx1626), .A0 (nx17823), .A1 (nx1558)) ;
    nand04 ix2883 (.Y (Dout[17]), .A0 (nx16043), .A1 (nx16054), .A2 (nx16071), .A3 (
           nx16102)) ;
    aoi222 ix16044 (.Y (nx16043), .A0 (Mem_28__1), .A1 (nx17441), .B0 (Mem_24__1
           ), .B1 (nx17835), .C0 (Mem_17__1), .C1 (nx17837)) ;
    dff reg_Mem_28__1 (.Q (Mem_28__1), .QB (nx16047), .D (nx13764), .CLK (CLK)
        ) ;
    dff reg_Mem_24__1 (.Q (Mem_24__1), .QB (\$dummy [45]), .D (nx13774), .CLK (
        CLK)) ;
    mux21_ni ix13775 (.Y (nx13774), .A0 (Din[1]), .A1 (Mem_24__1), .S0 (nx17569)
             ) ;
    dff reg_Mem_17__1 (.Q (Mem_17__1), .QB (nx16053), .D (nx13784), .CLK (CLK)
        ) ;
    aoi221 ix16055 (.Y (nx16054), .A0 (Mem_16__1), .A1 (nx17737), .B0 (Mem_23__1
           ), .B1 (nx17733), .C0 (nx2828)) ;
    dff reg_Mem_16__1 (.Q (Mem_16__1), .QB (nx16058), .D (nx13754), .CLK (CLK)
        ) ;
    dff reg_Mem_23__1 (.Q (Mem_23__1), .QB (\$dummy [46]), .D (nx13744), .CLK (
        CLK)) ;
    mux21_ni ix13745 (.Y (nx13744), .A0 (Mem_23__1), .A1 (Din[1]), .S0 (nx17433)
             ) ;
    oai22 ix2829 (.Y (nx2828), .A0 (nx16063), .A1 (nx15821), .B0 (nx16067), .B1 (
          nx17583)) ;
    dff reg_Mem_14__1 (.Q (Mem_14__1), .QB (nx16063), .D (nx13734), .CLK (CLK)
        ) ;
    dff reg_Mem_12__1 (.Q (Mem_12__1), .QB (nx16067), .D (nx13724), .CLK (CLK)
        ) ;
    and04 ix16072 (.Y (nx16071), .A0 (nx16073), .A1 (nx16081), .A2 (nx16089), .A3 (
          nx16094)) ;
    aoi22 ix16074 (.Y (nx16073), .A0 (Mem_19__1), .A1 (nx17729), .B0 (Mem_13__1)
          , .B1 (nx2336)) ;
    dff reg_Mem_19__1 (.Q (Mem_19__1), .QB (nx16077), .D (nx13704), .CLK (CLK)
        ) ;
    dff reg_Mem_13__1 (.Q (Mem_13__1), .QB (\$dummy [47]), .D (nx13714), .CLK (
        CLK)) ;
    mux21_ni ix13715 (.Y (nx13714), .A0 (Mem_13__1), .A1 (Din[1]), .S0 (nx17429)
             ) ;
    aoi22 ix16082 (.Y (nx16081), .A0 (Mem_10__1), .A1 (nx17725), .B0 (Mem_15__1)
          , .B1 (nx2220)) ;
    dff reg_Mem_10__1 (.Q (Mem_10__1), .QB (\$dummy [48]), .D (nx13694), .CLK (
        CLK)) ;
    mux21_ni ix13695 (.Y (nx13694), .A0 (Din[1]), .A1 (Mem_10__1), .S0 (nx17587)
             ) ;
    dff reg_Mem_15__1 (.Q (Mem_15__1), .QB (\$dummy [49]), .D (nx13684), .CLK (
        CLK)) ;
    mux21_ni ix13685 (.Y (nx13684), .A0 (Mem_15__1), .A1 (Din[1]), .S0 (nx17421)
             ) ;
    aoi22 ix16090 (.Y (nx16089), .A0 (Mem_9__1), .A1 (nx17721), .B0 (Mem_8__1), 
          .B1 (nx17717)) ;
    dff reg_Mem_9__1 (.Q (Mem_9__1), .QB (\$dummy [50]), .D (nx13674), .CLK (CLK
        )) ;
    mux21_ni ix13675 (.Y (nx13674), .A0 (Mem_9__1), .A1 (Din[1]), .S0 (nx17417)
             ) ;
    aoi22 ix16095 (.Y (nx16094), .A0 (Mem_29__1), .A1 (nx17709), .B0 (Mem_18__1)
          , .B1 (nx17713)) ;
    dff reg_Mem_29__1 (.Q (Mem_29__1), .QB (nx16098), .D (nx13654), .CLK (CLK)
        ) ;
    dff reg_Mem_18__1 (.Q (Mem_18__1), .QB (\$dummy [51]), .D (nx13664), .CLK (
        CLK)) ;
    mux21_ni ix13665 (.Y (nx13664), .A0 (Mem_18__1), .A1 (Din[1]), .S0 (nx17413)
             ) ;
    nor04 ix16103 (.Y (nx16102), .A0 (nx2736), .A1 (nx2670), .A2 (nx2664), .A3 (
          nx2658)) ;
    nand03 ix2737 (.Y (nx2736), .A0 (nx16105), .A1 (nx16116), .A2 (nx16124)) ;
    aoi222 ix16106 (.Y (nx16105), .A0 (Mem_31__1), .A1 (nx17405), .B0 (Mem_30__1
           ), .B1 (nx17833), .C0 (Mem_11__1), .C1 (nx17831)) ;
    dff reg_Mem_31__1 (.Q (Mem_31__1), .QB (nx16109), .D (nx13644), .CLK (CLK)
        ) ;
    dff reg_Mem_30__1 (.Q (Mem_30__1), .QB (\$dummy [52]), .D (nx13634), .CLK (
        CLK)) ;
    mux21_ni ix13635 (.Y (nx13634), .A0 (Din[1]), .A1 (Mem_30__1), .S0 (nx17595)
             ) ;
    dff reg_Mem_11__1 (.Q (Mem_11__1), .QB (\$dummy [53]), .D (nx13624), .CLK (
        CLK)) ;
    mux21_ni ix13625 (.Y (nx13624), .A0 (Mem_11__1), .A1 (Din[1]), .S0 (nx17397)
             ) ;
    aoi22 ix16117 (.Y (nx16116), .A0 (Mem_26__1), .A1 (nx17705), .B0 (Mem_25__1)
          , .B1 (nx17701)) ;
    dff reg_Mem_26__1 (.Q (Mem_26__1), .QB (\$dummy [54]), .D (nx13614), .CLK (
        CLK)) ;
    mux21_ni ix13615 (.Y (nx13614), .A0 (Din[1]), .A1 (Mem_26__1), .S0 (nx17599)
             ) ;
    dff reg_Mem_25__1 (.Q (Mem_25__1), .QB (\$dummy [55]), .D (nx13604), .CLK (
        CLK)) ;
    mux21_ni ix13605 (.Y (nx13604), .A0 (Mem_25__1), .A1 (Din[1]), .S0 (nx17393)
             ) ;
    aoi22 ix16125 (.Y (nx16124), .A0 (Mem_27__1), .A1 (nx17697), .B0 (Mem_2__1)
          , .B1 (nx17389)) ;
    dff reg_Mem_27__1 (.Q (Mem_27__1), .QB (\$dummy [56]), .D (nx13594), .CLK (
        CLK)) ;
    mux21_ni ix13595 (.Y (nx13594), .A0 (Din[1]), .A1 (Mem_27__1), .S0 (nx17603)
             ) ;
    oai22 ix2671 (.Y (nx2670), .A0 (nx15383), .A1 (nx16000), .B0 (nx15370), .B1 (
          nx17607)) ;
    oai22 ix2665 (.Y (nx2664), .A0 (nx15362), .A1 (nx16006), .B0 (nx15375), .B1 (
          nx16008)) ;
    oai221 ix2659 (.Y (nx2658), .A0 (nx15378), .A1 (nx17611), .B0 (nx16132), .B1 (
           nx17613), .C0 (nx16136)) ;
    dff reg_Mem_21__1 (.Q (Mem_21__1), .QB (nx16132), .D (nx13564), .CLK (CLK)
        ) ;
    aoi22 ix16137 (.Y (nx16136), .A0 (Mem_20__1), .A1 (nx1674), .B0 (Mem_22__1)
          , .B1 (nx1626)) ;
    dff reg_Mem_20__1 (.Q (Mem_20__1), .QB (nx16140), .D (nx13584), .CLK (CLK)
        ) ;
    dff reg_Mem_22__1 (.Q (Mem_22__1), .QB (\$dummy [57]), .D (nx13574), .CLK (
        CLK)) ;
    mux21_ni ix13575 (.Y (nx13574), .A0 (Mem_22__1), .A1 (Din[1]), .S0 (nx17381)
             ) ;
    nand04 ix3139 (.Y (Dout[18]), .A0 (nx16145), .A1 (nx16156), .A2 (nx16173), .A3 (
           nx16204)) ;
    aoi222 ix16146 (.Y (nx16145), .A0 (Mem_28__2), .A1 (nx17441), .B0 (Mem_24__2
           ), .B1 (nx17835), .C0 (Mem_17__2), .C1 (nx17837)) ;
    dff reg_Mem_28__2 (.Q (Mem_28__2), .QB (nx16149), .D (nx13994), .CLK (CLK)
        ) ;
    dff reg_Mem_24__2 (.Q (Mem_24__2), .QB (\$dummy [58]), .D (nx14004), .CLK (
        CLK)) ;
    mux21_ni ix14005 (.Y (nx14004), .A0 (Din[2]), .A1 (Mem_24__2), .S0 (nx17569)
             ) ;
    dff reg_Mem_17__2 (.Q (Mem_17__2), .QB (nx16155), .D (nx14014), .CLK (CLK)
        ) ;
    aoi221 ix16157 (.Y (nx16156), .A0 (Mem_16__2), .A1 (nx17737), .B0 (Mem_23__2
           ), .B1 (nx17733), .C0 (nx3084)) ;
    dff reg_Mem_16__2 (.Q (Mem_16__2), .QB (nx16160), .D (nx13984), .CLK (CLK)
        ) ;
    dff reg_Mem_23__2 (.Q (Mem_23__2), .QB (\$dummy [59]), .D (nx13974), .CLK (
        CLK)) ;
    mux21_ni ix13975 (.Y (nx13974), .A0 (Mem_23__2), .A1 (Din[2]), .S0 (nx17433)
             ) ;
    oai22 ix3085 (.Y (nx3084), .A0 (nx16165), .A1 (nx15821), .B0 (nx16169), .B1 (
          nx17583)) ;
    dff reg_Mem_14__2 (.Q (Mem_14__2), .QB (nx16165), .D (nx13964), .CLK (CLK)
        ) ;
    dff reg_Mem_12__2 (.Q (Mem_12__2), .QB (nx16169), .D (nx13954), .CLK (CLK)
        ) ;
    and04 ix16174 (.Y (nx16173), .A0 (nx16175), .A1 (nx16183), .A2 (nx16191), .A3 (
          nx16196)) ;
    aoi22 ix16176 (.Y (nx16175), .A0 (Mem_19__2), .A1 (nx17729), .B0 (Mem_13__2)
          , .B1 (nx2336)) ;
    dff reg_Mem_19__2 (.Q (Mem_19__2), .QB (nx16179), .D (nx13934), .CLK (CLK)
        ) ;
    dff reg_Mem_13__2 (.Q (Mem_13__2), .QB (\$dummy [60]), .D (nx13944), .CLK (
        CLK)) ;
    mux21_ni ix13945 (.Y (nx13944), .A0 (Mem_13__2), .A1 (Din[2]), .S0 (nx17429)
             ) ;
    aoi22 ix16184 (.Y (nx16183), .A0 (Mem_10__2), .A1 (nx17725), .B0 (Mem_15__2)
          , .B1 (nx2220)) ;
    dff reg_Mem_10__2 (.Q (Mem_10__2), .QB (\$dummy [61]), .D (nx13924), .CLK (
        CLK)) ;
    mux21_ni ix13925 (.Y (nx13924), .A0 (Din[2]), .A1 (Mem_10__2), .S0 (nx17587)
             ) ;
    dff reg_Mem_15__2 (.Q (Mem_15__2), .QB (\$dummy [62]), .D (nx13914), .CLK (
        CLK)) ;
    mux21_ni ix13915 (.Y (nx13914), .A0 (Mem_15__2), .A1 (Din[2]), .S0 (nx17421)
             ) ;
    aoi22 ix16192 (.Y (nx16191), .A0 (Mem_9__2), .A1 (nx17721), .B0 (Mem_8__2), 
          .B1 (nx17717)) ;
    dff reg_Mem_9__2 (.Q (Mem_9__2), .QB (\$dummy [63]), .D (nx13904), .CLK (CLK
        )) ;
    mux21_ni ix13905 (.Y (nx13904), .A0 (Mem_9__2), .A1 (Din[2]), .S0 (nx17417)
             ) ;
    aoi22 ix16197 (.Y (nx16196), .A0 (Mem_29__2), .A1 (nx17709), .B0 (Mem_18__2)
          , .B1 (nx17713)) ;
    dff reg_Mem_29__2 (.Q (Mem_29__2), .QB (nx16200), .D (nx13884), .CLK (CLK)
        ) ;
    dff reg_Mem_18__2 (.Q (Mem_18__2), .QB (\$dummy [64]), .D (nx13894), .CLK (
        CLK)) ;
    mux21_ni ix13895 (.Y (nx13894), .A0 (Mem_18__2), .A1 (Din[2]), .S0 (nx17413)
             ) ;
    nor04 ix16205 (.Y (nx16204), .A0 (nx2992), .A1 (nx2926), .A2 (nx2920), .A3 (
          nx2914)) ;
    nand03 ix2993 (.Y (nx2992), .A0 (nx16207), .A1 (nx16218), .A2 (nx16226)) ;
    aoi222 ix16208 (.Y (nx16207), .A0 (Mem_31__2), .A1 (nx17405), .B0 (Mem_30__2
           ), .B1 (nx17833), .C0 (Mem_11__2), .C1 (nx17831)) ;
    dff reg_Mem_31__2 (.Q (Mem_31__2), .QB (nx16211), .D (nx13874), .CLK (CLK)
        ) ;
    dff reg_Mem_30__2 (.Q (Mem_30__2), .QB (\$dummy [65]), .D (nx13864), .CLK (
        CLK)) ;
    mux21_ni ix13865 (.Y (nx13864), .A0 (Din[2]), .A1 (Mem_30__2), .S0 (nx17595)
             ) ;
    dff reg_Mem_11__2 (.Q (Mem_11__2), .QB (\$dummy [66]), .D (nx13854), .CLK (
        CLK)) ;
    mux21_ni ix13855 (.Y (nx13854), .A0 (Mem_11__2), .A1 (Din[2]), .S0 (nx17397)
             ) ;
    aoi22 ix16219 (.Y (nx16218), .A0 (Mem_26__2), .A1 (nx17705), .B0 (Mem_25__2)
          , .B1 (nx17701)) ;
    dff reg_Mem_26__2 (.Q (Mem_26__2), .QB (\$dummy [67]), .D (nx13844), .CLK (
        CLK)) ;
    mux21_ni ix13845 (.Y (nx13844), .A0 (Din[2]), .A1 (Mem_26__2), .S0 (nx17599)
             ) ;
    dff reg_Mem_25__2 (.Q (Mem_25__2), .QB (\$dummy [68]), .D (nx13834), .CLK (
        CLK)) ;
    mux21_ni ix13835 (.Y (nx13834), .A0 (Mem_25__2), .A1 (Din[2]), .S0 (nx17393)
             ) ;
    aoi22 ix16227 (.Y (nx16226), .A0 (Mem_27__2), .A1 (nx17697), .B0 (Mem_2__2)
          , .B1 (nx17389)) ;
    dff reg_Mem_27__2 (.Q (Mem_27__2), .QB (\$dummy [69]), .D (nx13824), .CLK (
        CLK)) ;
    mux21_ni ix13825 (.Y (nx13824), .A0 (Din[2]), .A1 (Mem_27__2), .S0 (nx17603)
             ) ;
    oai22 ix2927 (.Y (nx2926), .A0 (nx15416), .A1 (nx16000), .B0 (nx15403), .B1 (
          nx17607)) ;
    oai22 ix2921 (.Y (nx2920), .A0 (nx15395), .A1 (nx16006), .B0 (nx15408), .B1 (
          nx16008)) ;
    oai221 ix2915 (.Y (nx2914), .A0 (nx15411), .A1 (nx17611), .B0 (nx16234), .B1 (
           nx17613), .C0 (nx16238)) ;
    dff reg_Mem_21__2 (.Q (Mem_21__2), .QB (nx16234), .D (nx13794), .CLK (CLK)
        ) ;
    aoi22 ix16239 (.Y (nx16238), .A0 (Mem_20__2), .A1 (nx1674), .B0 (Mem_22__2)
          , .B1 (nx1626)) ;
    dff reg_Mem_20__2 (.Q (Mem_20__2), .QB (nx16242), .D (nx13814), .CLK (CLK)
        ) ;
    dff reg_Mem_22__2 (.Q (Mem_22__2), .QB (\$dummy [70]), .D (nx13804), .CLK (
        CLK)) ;
    mux21_ni ix13805 (.Y (nx13804), .A0 (Mem_22__2), .A1 (Din[2]), .S0 (nx17381)
             ) ;
    nand04 ix3395 (.Y (Dout[19]), .A0 (nx16247), .A1 (nx16258), .A2 (nx16275), .A3 (
           nx16306)) ;
    aoi222 ix16248 (.Y (nx16247), .A0 (Mem_28__3), .A1 (nx17441), .B0 (Mem_24__3
           ), .B1 (nx17835), .C0 (Mem_17__3), .C1 (nx17837)) ;
    dff reg_Mem_28__3 (.Q (Mem_28__3), .QB (nx16251), .D (nx14224), .CLK (CLK)
        ) ;
    dff reg_Mem_24__3 (.Q (Mem_24__3), .QB (\$dummy [71]), .D (nx14234), .CLK (
        CLK)) ;
    mux21_ni ix14235 (.Y (nx14234), .A0 (Din[3]), .A1 (Mem_24__3), .S0 (nx17569)
             ) ;
    dff reg_Mem_17__3 (.Q (Mem_17__3), .QB (nx16257), .D (nx14244), .CLK (CLK)
        ) ;
    aoi221 ix16259 (.Y (nx16258), .A0 (Mem_16__3), .A1 (nx17737), .B0 (Mem_23__3
           ), .B1 (nx17733), .C0 (nx3340)) ;
    dff reg_Mem_16__3 (.Q (Mem_16__3), .QB (nx16262), .D (nx14214), .CLK (CLK)
        ) ;
    dff reg_Mem_23__3 (.Q (Mem_23__3), .QB (\$dummy [72]), .D (nx14204), .CLK (
        CLK)) ;
    mux21_ni ix14205 (.Y (nx14204), .A0 (Mem_23__3), .A1 (Din[3]), .S0 (nx17433)
             ) ;
    oai22 ix3341 (.Y (nx3340), .A0 (nx16267), .A1 (nx15821), .B0 (nx16271), .B1 (
          nx17583)) ;
    dff reg_Mem_14__3 (.Q (Mem_14__3), .QB (nx16267), .D (nx14194), .CLK (CLK)
        ) ;
    dff reg_Mem_12__3 (.Q (Mem_12__3), .QB (nx16271), .D (nx14184), .CLK (CLK)
        ) ;
    and04 ix16276 (.Y (nx16275), .A0 (nx16277), .A1 (nx16285), .A2 (nx16293), .A3 (
          nx16298)) ;
    aoi22 ix16278 (.Y (nx16277), .A0 (Mem_19__3), .A1 (nx17729), .B0 (Mem_13__3)
          , .B1 (nx2336)) ;
    dff reg_Mem_19__3 (.Q (Mem_19__3), .QB (nx16281), .D (nx14164), .CLK (CLK)
        ) ;
    dff reg_Mem_13__3 (.Q (Mem_13__3), .QB (\$dummy [73]), .D (nx14174), .CLK (
        CLK)) ;
    mux21_ni ix14175 (.Y (nx14174), .A0 (Mem_13__3), .A1 (Din[3]), .S0 (nx17429)
             ) ;
    aoi22 ix16286 (.Y (nx16285), .A0 (Mem_10__3), .A1 (nx17725), .B0 (Mem_15__3)
          , .B1 (nx2220)) ;
    dff reg_Mem_10__3 (.Q (Mem_10__3), .QB (\$dummy [74]), .D (nx14154), .CLK (
        CLK)) ;
    mux21_ni ix14155 (.Y (nx14154), .A0 (Din[3]), .A1 (Mem_10__3), .S0 (nx17587)
             ) ;
    dff reg_Mem_15__3 (.Q (Mem_15__3), .QB (\$dummy [75]), .D (nx14144), .CLK (
        CLK)) ;
    mux21_ni ix14145 (.Y (nx14144), .A0 (Mem_15__3), .A1 (Din[3]), .S0 (nx17421)
             ) ;
    aoi22 ix16294 (.Y (nx16293), .A0 (Mem_9__3), .A1 (nx17721), .B0 (Mem_8__3), 
          .B1 (nx17717)) ;
    dff reg_Mem_9__3 (.Q (Mem_9__3), .QB (\$dummy [76]), .D (nx14134), .CLK (CLK
        )) ;
    mux21_ni ix14135 (.Y (nx14134), .A0 (Mem_9__3), .A1 (Din[3]), .S0 (nx17417)
             ) ;
    aoi22 ix16299 (.Y (nx16298), .A0 (Mem_29__3), .A1 (nx17709), .B0 (Mem_18__3)
          , .B1 (nx17713)) ;
    dff reg_Mem_29__3 (.Q (Mem_29__3), .QB (nx16302), .D (nx14114), .CLK (CLK)
        ) ;
    dff reg_Mem_18__3 (.Q (Mem_18__3), .QB (\$dummy [77]), .D (nx14124), .CLK (
        CLK)) ;
    mux21_ni ix14125 (.Y (nx14124), .A0 (Mem_18__3), .A1 (Din[3]), .S0 (nx17413)
             ) ;
    nor04 ix16307 (.Y (nx16306), .A0 (nx3248), .A1 (nx3182), .A2 (nx3176), .A3 (
          nx3170)) ;
    nand03 ix3249 (.Y (nx3248), .A0 (nx16309), .A1 (nx16320), .A2 (nx16328)) ;
    aoi222 ix16310 (.Y (nx16309), .A0 (Mem_31__3), .A1 (nx17405), .B0 (Mem_30__3
           ), .B1 (nx17833), .C0 (Mem_11__3), .C1 (nx17831)) ;
    dff reg_Mem_31__3 (.Q (Mem_31__3), .QB (nx16313), .D (nx14104), .CLK (CLK)
        ) ;
    dff reg_Mem_30__3 (.Q (Mem_30__3), .QB (\$dummy [78]), .D (nx14094), .CLK (
        CLK)) ;
    mux21_ni ix14095 (.Y (nx14094), .A0 (Din[3]), .A1 (Mem_30__3), .S0 (nx17595)
             ) ;
    dff reg_Mem_11__3 (.Q (Mem_11__3), .QB (\$dummy [79]), .D (nx14084), .CLK (
        CLK)) ;
    mux21_ni ix14085 (.Y (nx14084), .A0 (Mem_11__3), .A1 (Din[3]), .S0 (nx17397)
             ) ;
    aoi22 ix16321 (.Y (nx16320), .A0 (Mem_26__3), .A1 (nx17705), .B0 (Mem_25__3)
          , .B1 (nx17701)) ;
    dff reg_Mem_26__3 (.Q (Mem_26__3), .QB (\$dummy [80]), .D (nx14074), .CLK (
        CLK)) ;
    mux21_ni ix14075 (.Y (nx14074), .A0 (Din[3]), .A1 (Mem_26__3), .S0 (nx17599)
             ) ;
    dff reg_Mem_25__3 (.Q (Mem_25__3), .QB (\$dummy [81]), .D (nx14064), .CLK (
        CLK)) ;
    mux21_ni ix14065 (.Y (nx14064), .A0 (Mem_25__3), .A1 (Din[3]), .S0 (nx17393)
             ) ;
    aoi22 ix16329 (.Y (nx16328), .A0 (Mem_27__3), .A1 (nx17697), .B0 (Mem_2__3)
          , .B1 (nx17389)) ;
    dff reg_Mem_27__3 (.Q (Mem_27__3), .QB (\$dummy [82]), .D (nx14054), .CLK (
        CLK)) ;
    mux21_ni ix14055 (.Y (nx14054), .A0 (Din[3]), .A1 (Mem_27__3), .S0 (nx17603)
             ) ;
    oai22 ix3183 (.Y (nx3182), .A0 (nx15449), .A1 (nx16000), .B0 (nx15436), .B1 (
          nx17607)) ;
    oai22 ix3177 (.Y (nx3176), .A0 (nx15428), .A1 (nx16006), .B0 (nx15441), .B1 (
          nx16008)) ;
    oai221 ix3171 (.Y (nx3170), .A0 (nx15444), .A1 (nx17611), .B0 (nx16336), .B1 (
           nx17613), .C0 (nx16340)) ;
    dff reg_Mem_21__3 (.Q (Mem_21__3), .QB (nx16336), .D (nx14024), .CLK (CLK)
        ) ;
    aoi22 ix16341 (.Y (nx16340), .A0 (Mem_20__3), .A1 (nx1674), .B0 (Mem_22__3)
          , .B1 (nx1626)) ;
    dff reg_Mem_20__3 (.Q (Mem_20__3), .QB (nx16344), .D (nx14044), .CLK (CLK)
        ) ;
    dff reg_Mem_22__3 (.Q (Mem_22__3), .QB (\$dummy [83]), .D (nx14034), .CLK (
        CLK)) ;
    mux21_ni ix14035 (.Y (nx14034), .A0 (Mem_22__3), .A1 (Din[3]), .S0 (nx17381)
             ) ;
    nand04 ix3651 (.Y (Dout[20]), .A0 (nx16349), .A1 (nx16360), .A2 (nx16377), .A3 (
           nx16408)) ;
    aoi222 ix16350 (.Y (nx16349), .A0 (Mem_28__4), .A1 (nx17441), .B0 (Mem_24__4
           ), .B1 (nx17835), .C0 (Mem_17__4), .C1 (nx17837)) ;
    dff reg_Mem_28__4 (.Q (Mem_28__4), .QB (nx16353), .D (nx14454), .CLK (CLK)
        ) ;
    dff reg_Mem_24__4 (.Q (Mem_24__4), .QB (\$dummy [84]), .D (nx14464), .CLK (
        CLK)) ;
    mux21_ni ix14465 (.Y (nx14464), .A0 (Din[4]), .A1 (Mem_24__4), .S0 (nx17569)
             ) ;
    dff reg_Mem_17__4 (.Q (Mem_17__4), .QB (nx16359), .D (nx14474), .CLK (CLK)
        ) ;
    aoi221 ix16361 (.Y (nx16360), .A0 (Mem_16__4), .A1 (nx17737), .B0 (Mem_23__4
           ), .B1 (nx17733), .C0 (nx3596)) ;
    dff reg_Mem_16__4 (.Q (Mem_16__4), .QB (nx16364), .D (nx14444), .CLK (CLK)
        ) ;
    dff reg_Mem_23__4 (.Q (Mem_23__4), .QB (\$dummy [85]), .D (nx14434), .CLK (
        CLK)) ;
    mux21_ni ix14435 (.Y (nx14434), .A0 (Mem_23__4), .A1 (Din[4]), .S0 (nx17433)
             ) ;
    oai22 ix3597 (.Y (nx3596), .A0 (nx16369), .A1 (nx15821), .B0 (nx16373), .B1 (
          nx17583)) ;
    dff reg_Mem_14__4 (.Q (Mem_14__4), .QB (nx16369), .D (nx14424), .CLK (CLK)
        ) ;
    dff reg_Mem_12__4 (.Q (Mem_12__4), .QB (nx16373), .D (nx14414), .CLK (CLK)
        ) ;
    and04 ix16378 (.Y (nx16377), .A0 (nx16379), .A1 (nx16387), .A2 (nx16395), .A3 (
          nx16400)) ;
    aoi22 ix16380 (.Y (nx16379), .A0 (Mem_19__4), .A1 (nx17729), .B0 (Mem_13__4)
          , .B1 (nx2336)) ;
    dff reg_Mem_19__4 (.Q (Mem_19__4), .QB (nx16383), .D (nx14394), .CLK (CLK)
        ) ;
    dff reg_Mem_13__4 (.Q (Mem_13__4), .QB (\$dummy [86]), .D (nx14404), .CLK (
        CLK)) ;
    mux21_ni ix14405 (.Y (nx14404), .A0 (Mem_13__4), .A1 (Din[4]), .S0 (nx17429)
             ) ;
    aoi22 ix16388 (.Y (nx16387), .A0 (Mem_10__4), .A1 (nx17725), .B0 (Mem_15__4)
          , .B1 (nx2220)) ;
    dff reg_Mem_10__4 (.Q (Mem_10__4), .QB (\$dummy [87]), .D (nx14384), .CLK (
        CLK)) ;
    mux21_ni ix14385 (.Y (nx14384), .A0 (Din[4]), .A1 (Mem_10__4), .S0 (nx17587)
             ) ;
    dff reg_Mem_15__4 (.Q (Mem_15__4), .QB (\$dummy [88]), .D (nx14374), .CLK (
        CLK)) ;
    mux21_ni ix14375 (.Y (nx14374), .A0 (Mem_15__4), .A1 (Din[4]), .S0 (nx17421)
             ) ;
    aoi22 ix16396 (.Y (nx16395), .A0 (Mem_9__4), .A1 (nx17721), .B0 (Mem_8__4), 
          .B1 (nx17717)) ;
    dff reg_Mem_9__4 (.Q (Mem_9__4), .QB (\$dummy [89]), .D (nx14364), .CLK (CLK
        )) ;
    mux21_ni ix14365 (.Y (nx14364), .A0 (Mem_9__4), .A1 (Din[4]), .S0 (nx17417)
             ) ;
    aoi22 ix16401 (.Y (nx16400), .A0 (Mem_29__4), .A1 (nx17709), .B0 (Mem_18__4)
          , .B1 (nx17713)) ;
    dff reg_Mem_29__4 (.Q (Mem_29__4), .QB (nx16404), .D (nx14344), .CLK (CLK)
        ) ;
    dff reg_Mem_18__4 (.Q (Mem_18__4), .QB (\$dummy [90]), .D (nx14354), .CLK (
        CLK)) ;
    mux21_ni ix14355 (.Y (nx14354), .A0 (Mem_18__4), .A1 (Din[4]), .S0 (nx17413)
             ) ;
    nor04 ix16409 (.Y (nx16408), .A0 (nx3504), .A1 (nx3438), .A2 (nx3432), .A3 (
          nx3426)) ;
    nand03 ix3505 (.Y (nx3504), .A0 (nx16411), .A1 (nx16422), .A2 (nx16430)) ;
    aoi222 ix16412 (.Y (nx16411), .A0 (Mem_31__4), .A1 (nx17405), .B0 (Mem_30__4
           ), .B1 (nx17833), .C0 (Mem_11__4), .C1 (nx17831)) ;
    dff reg_Mem_31__4 (.Q (Mem_31__4), .QB (nx16415), .D (nx14334), .CLK (CLK)
        ) ;
    dff reg_Mem_30__4 (.Q (Mem_30__4), .QB (\$dummy [91]), .D (nx14324), .CLK (
        CLK)) ;
    mux21_ni ix14325 (.Y (nx14324), .A0 (Din[4]), .A1 (Mem_30__4), .S0 (nx17595)
             ) ;
    dff reg_Mem_11__4 (.Q (Mem_11__4), .QB (\$dummy [92]), .D (nx14314), .CLK (
        CLK)) ;
    mux21_ni ix14315 (.Y (nx14314), .A0 (Mem_11__4), .A1 (Din[4]), .S0 (nx17397)
             ) ;
    aoi22 ix16423 (.Y (nx16422), .A0 (Mem_26__4), .A1 (nx17705), .B0 (Mem_25__4)
          , .B1 (nx17701)) ;
    dff reg_Mem_26__4 (.Q (Mem_26__4), .QB (\$dummy [93]), .D (nx14304), .CLK (
        CLK)) ;
    mux21_ni ix14305 (.Y (nx14304), .A0 (Din[4]), .A1 (Mem_26__4), .S0 (nx17599)
             ) ;
    dff reg_Mem_25__4 (.Q (Mem_25__4), .QB (\$dummy [94]), .D (nx14294), .CLK (
        CLK)) ;
    mux21_ni ix14295 (.Y (nx14294), .A0 (Mem_25__4), .A1 (Din[4]), .S0 (nx17393)
             ) ;
    aoi22 ix16431 (.Y (nx16430), .A0 (Mem_27__4), .A1 (nx17697), .B0 (Mem_2__4)
          , .B1 (nx17389)) ;
    dff reg_Mem_27__4 (.Q (Mem_27__4), .QB (\$dummy [95]), .D (nx14284), .CLK (
        CLK)) ;
    mux21_ni ix14285 (.Y (nx14284), .A0 (Din[4]), .A1 (Mem_27__4), .S0 (nx17603)
             ) ;
    oai22 ix3439 (.Y (nx3438), .A0 (nx15482), .A1 (nx16000), .B0 (nx15469), .B1 (
          nx17607)) ;
    oai22 ix3433 (.Y (nx3432), .A0 (nx15461), .A1 (nx16006), .B0 (nx15474), .B1 (
          nx16008)) ;
    oai221 ix3427 (.Y (nx3426), .A0 (nx15477), .A1 (nx17611), .B0 (nx16438), .B1 (
           nx17613), .C0 (nx16442)) ;
    dff reg_Mem_21__4 (.Q (Mem_21__4), .QB (nx16438), .D (nx14254), .CLK (CLK)
        ) ;
    aoi22 ix16443 (.Y (nx16442), .A0 (Mem_20__4), .A1 (nx1674), .B0 (Mem_22__4)
          , .B1 (nx1626)) ;
    dff reg_Mem_20__4 (.Q (Mem_20__4), .QB (nx16446), .D (nx14274), .CLK (CLK)
        ) ;
    dff reg_Mem_22__4 (.Q (Mem_22__4), .QB (\$dummy [96]), .D (nx14264), .CLK (
        CLK)) ;
    mux21_ni ix14265 (.Y (nx14264), .A0 (Mem_22__4), .A1 (Din[4]), .S0 (nx17381)
             ) ;
    nand04 ix3907 (.Y (Dout[21]), .A0 (nx16451), .A1 (nx16462), .A2 (nx16479), .A3 (
           nx16510)) ;
    aoi222 ix16452 (.Y (nx16451), .A0 (Mem_28__5), .A1 (nx17441), .B0 (Mem_24__5
           ), .B1 (nx17835), .C0 (Mem_17__5), .C1 (nx17837)) ;
    dff reg_Mem_28__5 (.Q (Mem_28__5), .QB (nx16455), .D (nx14684), .CLK (CLK)
        ) ;
    dff reg_Mem_24__5 (.Q (Mem_24__5), .QB (\$dummy [97]), .D (nx14694), .CLK (
        CLK)) ;
    mux21_ni ix14695 (.Y (nx14694), .A0 (Din[5]), .A1 (Mem_24__5), .S0 (nx17569)
             ) ;
    dff reg_Mem_17__5 (.Q (Mem_17__5), .QB (nx16461), .D (nx14704), .CLK (CLK)
        ) ;
    aoi221 ix16463 (.Y (nx16462), .A0 (Mem_16__5), .A1 (nx17737), .B0 (Mem_23__5
           ), .B1 (nx17733), .C0 (nx3852)) ;
    dff reg_Mem_16__5 (.Q (Mem_16__5), .QB (nx16466), .D (nx14674), .CLK (CLK)
        ) ;
    dff reg_Mem_23__5 (.Q (Mem_23__5), .QB (\$dummy [98]), .D (nx14664), .CLK (
        CLK)) ;
    mux21_ni ix14665 (.Y (nx14664), .A0 (Mem_23__5), .A1 (Din[5]), .S0 (nx17433)
             ) ;
    oai22 ix3853 (.Y (nx3852), .A0 (nx16471), .A1 (nx15821), .B0 (nx16475), .B1 (
          nx17583)) ;
    dff reg_Mem_14__5 (.Q (Mem_14__5), .QB (nx16471), .D (nx14654), .CLK (CLK)
        ) ;
    dff reg_Mem_12__5 (.Q (Mem_12__5), .QB (nx16475), .D (nx14644), .CLK (CLK)
        ) ;
    and04 ix16480 (.Y (nx16479), .A0 (nx16481), .A1 (nx16489), .A2 (nx16497), .A3 (
          nx16502)) ;
    aoi22 ix16482 (.Y (nx16481), .A0 (Mem_19__5), .A1 (nx17729), .B0 (Mem_13__5)
          , .B1 (nx2336)) ;
    dff reg_Mem_19__5 (.Q (Mem_19__5), .QB (nx16485), .D (nx14624), .CLK (CLK)
        ) ;
    dff reg_Mem_13__5 (.Q (Mem_13__5), .QB (\$dummy [99]), .D (nx14634), .CLK (
        CLK)) ;
    mux21_ni ix14635 (.Y (nx14634), .A0 (Mem_13__5), .A1 (Din[5]), .S0 (nx17429)
             ) ;
    aoi22 ix16490 (.Y (nx16489), .A0 (Mem_10__5), .A1 (nx17725), .B0 (Mem_15__5)
          , .B1 (nx2220)) ;
    dff reg_Mem_10__5 (.Q (Mem_10__5), .QB (\$dummy [100]), .D (nx14614), .CLK (
        CLK)) ;
    mux21_ni ix14615 (.Y (nx14614), .A0 (Din[5]), .A1 (Mem_10__5), .S0 (nx17587)
             ) ;
    dff reg_Mem_15__5 (.Q (Mem_15__5), .QB (\$dummy [101]), .D (nx14604), .CLK (
        CLK)) ;
    mux21_ni ix14605 (.Y (nx14604), .A0 (Mem_15__5), .A1 (Din[5]), .S0 (nx17421)
             ) ;
    aoi22 ix16498 (.Y (nx16497), .A0 (Mem_9__5), .A1 (nx17721), .B0 (Mem_8__5), 
          .B1 (nx17717)) ;
    dff reg_Mem_9__5 (.Q (Mem_9__5), .QB (\$dummy [102]), .D (nx14594), .CLK (
        CLK)) ;
    mux21_ni ix14595 (.Y (nx14594), .A0 (Mem_9__5), .A1 (Din[5]), .S0 (nx17417)
             ) ;
    aoi22 ix16503 (.Y (nx16502), .A0 (Mem_29__5), .A1 (nx17709), .B0 (Mem_18__5)
          , .B1 (nx17713)) ;
    dff reg_Mem_29__5 (.Q (Mem_29__5), .QB (nx16506), .D (nx14574), .CLK (CLK)
        ) ;
    dff reg_Mem_18__5 (.Q (Mem_18__5), .QB (\$dummy [103]), .D (nx14584), .CLK (
        CLK)) ;
    mux21_ni ix14585 (.Y (nx14584), .A0 (Mem_18__5), .A1 (Din[5]), .S0 (nx17413)
             ) ;
    nor04 ix16511 (.Y (nx16510), .A0 (nx3760), .A1 (nx3694), .A2 (nx3688), .A3 (
          nx3682)) ;
    nand03 ix3761 (.Y (nx3760), .A0 (nx16513), .A1 (nx16524), .A2 (nx16532)) ;
    aoi222 ix16514 (.Y (nx16513), .A0 (Mem_31__5), .A1 (nx17405), .B0 (Mem_30__5
           ), .B1 (nx17833), .C0 (Mem_11__5), .C1 (nx17831)) ;
    dff reg_Mem_31__5 (.Q (Mem_31__5), .QB (nx16517), .D (nx14564), .CLK (CLK)
        ) ;
    dff reg_Mem_30__5 (.Q (Mem_30__5), .QB (\$dummy [104]), .D (nx14554), .CLK (
        CLK)) ;
    mux21_ni ix14555 (.Y (nx14554), .A0 (Din[5]), .A1 (Mem_30__5), .S0 (nx17595)
             ) ;
    dff reg_Mem_11__5 (.Q (Mem_11__5), .QB (\$dummy [105]), .D (nx14544), .CLK (
        CLK)) ;
    mux21_ni ix14545 (.Y (nx14544), .A0 (Mem_11__5), .A1 (Din[5]), .S0 (nx17397)
             ) ;
    aoi22 ix16525 (.Y (nx16524), .A0 (Mem_26__5), .A1 (nx17705), .B0 (Mem_25__5)
          , .B1 (nx17701)) ;
    dff reg_Mem_26__5 (.Q (Mem_26__5), .QB (\$dummy [106]), .D (nx14534), .CLK (
        CLK)) ;
    mux21_ni ix14535 (.Y (nx14534), .A0 (Din[5]), .A1 (Mem_26__5), .S0 (nx17599)
             ) ;
    dff reg_Mem_25__5 (.Q (Mem_25__5), .QB (\$dummy [107]), .D (nx14524), .CLK (
        CLK)) ;
    mux21_ni ix14525 (.Y (nx14524), .A0 (Mem_25__5), .A1 (Din[5]), .S0 (nx17393)
             ) ;
    aoi22 ix16533 (.Y (nx16532), .A0 (Mem_27__5), .A1 (nx17697), .B0 (Mem_2__5)
          , .B1 (nx17389)) ;
    dff reg_Mem_27__5 (.Q (Mem_27__5), .QB (\$dummy [108]), .D (nx14514), .CLK (
        CLK)) ;
    mux21_ni ix14515 (.Y (nx14514), .A0 (Din[5]), .A1 (Mem_27__5), .S0 (nx17603)
             ) ;
    oai22 ix3695 (.Y (nx3694), .A0 (nx15515), .A1 (nx16000), .B0 (nx15502), .B1 (
          nx17607)) ;
    oai22 ix3689 (.Y (nx3688), .A0 (nx15494), .A1 (nx16006), .B0 (nx15507), .B1 (
          nx16008)) ;
    oai221 ix3683 (.Y (nx3682), .A0 (nx15510), .A1 (nx16011), .B0 (nx16540), .B1 (
           nx16022), .C0 (nx16544)) ;
    dff reg_Mem_21__5 (.Q (Mem_21__5), .QB (nx16540), .D (nx14484), .CLK (CLK)
        ) ;
    aoi22 ix16545 (.Y (nx16544), .A0 (Mem_20__5), .A1 (nx1674), .B0 (Mem_22__5)
          , .B1 (nx1626)) ;
    dff reg_Mem_20__5 (.Q (Mem_20__5), .QB (nx16548), .D (nx14504), .CLK (CLK)
        ) ;
    dff reg_Mem_22__5 (.Q (Mem_22__5), .QB (\$dummy [109]), .D (nx14494), .CLK (
        CLK)) ;
    mux21_ni ix14495 (.Y (nx14494), .A0 (Mem_22__5), .A1 (Din[5]), .S0 (nx17381)
             ) ;
    nand04 ix4163 (.Y (Dout[22]), .A0 (nx16553), .A1 (nx16564), .A2 (nx16581), .A3 (
           nx16612)) ;
    aoi222 ix16554 (.Y (nx16553), .A0 (Mem_28__6), .A1 (nx17441), .B0 (Mem_24__6
           ), .B1 (nx2576), .C0 (Mem_17__6), .C1 (nx2614)) ;
    dff reg_Mem_28__6 (.Q (Mem_28__6), .QB (nx16557), .D (nx14914), .CLK (CLK)
        ) ;
    dff reg_Mem_24__6 (.Q (Mem_24__6), .QB (\$dummy [110]), .D (nx14924), .CLK (
        CLK)) ;
    mux21_ni ix14925 (.Y (nx14924), .A0 (Din[6]), .A1 (Mem_24__6), .S0 (nx17569)
             ) ;
    dff reg_Mem_17__6 (.Q (Mem_17__6), .QB (nx16563), .D (nx14934), .CLK (CLK)
        ) ;
    aoi221 ix16565 (.Y (nx16564), .A0 (Mem_16__6), .A1 (nx17737), .B0 (Mem_23__6
           ), .B1 (nx17733), .C0 (nx4108)) ;
    dff reg_Mem_16__6 (.Q (Mem_16__6), .QB (nx16568), .D (nx14904), .CLK (CLK)
        ) ;
    dff reg_Mem_23__6 (.Q (Mem_23__6), .QB (\$dummy [111]), .D (nx14894), .CLK (
        CLK)) ;
    mux21_ni ix14895 (.Y (nx14894), .A0 (Mem_23__6), .A1 (Din[6]), .S0 (nx17433)
             ) ;
    oai22 ix4109 (.Y (nx4108), .A0 (nx16573), .A1 (nx15821), .B0 (nx16577), .B1 (
          nx17583)) ;
    dff reg_Mem_14__6 (.Q (Mem_14__6), .QB (nx16573), .D (nx14884), .CLK (CLK)
        ) ;
    dff reg_Mem_12__6 (.Q (Mem_12__6), .QB (nx16577), .D (nx14874), .CLK (CLK)
        ) ;
    and04 ix16582 (.Y (nx16581), .A0 (nx16583), .A1 (nx16591), .A2 (nx16599), .A3 (
          nx16604)) ;
    aoi22 ix16584 (.Y (nx16583), .A0 (Mem_19__6), .A1 (nx17729), .B0 (Mem_13__6)
          , .B1 (nx2336)) ;
    dff reg_Mem_19__6 (.Q (Mem_19__6), .QB (nx16587), .D (nx14854), .CLK (CLK)
        ) ;
    dff reg_Mem_13__6 (.Q (Mem_13__6), .QB (\$dummy [112]), .D (nx14864), .CLK (
        CLK)) ;
    mux21_ni ix14865 (.Y (nx14864), .A0 (Mem_13__6), .A1 (Din[6]), .S0 (nx17429)
             ) ;
    aoi22 ix16592 (.Y (nx16591), .A0 (Mem_10__6), .A1 (nx17725), .B0 (Mem_15__6)
          , .B1 (nx2220)) ;
    dff reg_Mem_10__6 (.Q (Mem_10__6), .QB (\$dummy [113]), .D (nx14844), .CLK (
        CLK)) ;
    mux21_ni ix14845 (.Y (nx14844), .A0 (Din[6]), .A1 (Mem_10__6), .S0 (nx17587)
             ) ;
    dff reg_Mem_15__6 (.Q (Mem_15__6), .QB (\$dummy [114]), .D (nx14834), .CLK (
        CLK)) ;
    mux21_ni ix14835 (.Y (nx14834), .A0 (Mem_15__6), .A1 (Din[6]), .S0 (nx17421)
             ) ;
    aoi22 ix16600 (.Y (nx16599), .A0 (Mem_9__6), .A1 (nx17721), .B0 (Mem_8__6), 
          .B1 (nx17717)) ;
    dff reg_Mem_9__6 (.Q (Mem_9__6), .QB (\$dummy [115]), .D (nx14824), .CLK (
        CLK)) ;
    mux21_ni ix14825 (.Y (nx14824), .A0 (Mem_9__6), .A1 (Din[6]), .S0 (nx17417)
             ) ;
    aoi22 ix16605 (.Y (nx16604), .A0 (Mem_29__6), .A1 (nx17709), .B0 (Mem_18__6)
          , .B1 (nx17713)) ;
    dff reg_Mem_29__6 (.Q (Mem_29__6), .QB (nx16608), .D (nx14804), .CLK (CLK)
        ) ;
    dff reg_Mem_18__6 (.Q (Mem_18__6), .QB (\$dummy [116]), .D (nx14814), .CLK (
        CLK)) ;
    mux21_ni ix14815 (.Y (nx14814), .A0 (Mem_18__6), .A1 (Din[6]), .S0 (nx17413)
             ) ;
    nor04 ix16613 (.Y (nx16612), .A0 (nx4016), .A1 (nx3950), .A2 (nx3944), .A3 (
          nx3938)) ;
    nand03 ix4017 (.Y (nx4016), .A0 (nx16615), .A1 (nx16626), .A2 (nx16634)) ;
    aoi222 ix16616 (.Y (nx16615), .A0 (Mem_31__6), .A1 (nx17405), .B0 (Mem_30__6
           ), .B1 (nx1972), .C0 (Mem_11__6), .C1 (nx1916)) ;
    dff reg_Mem_31__6 (.Q (Mem_31__6), .QB (nx16619), .D (nx14794), .CLK (CLK)
        ) ;
    dff reg_Mem_30__6 (.Q (Mem_30__6), .QB (\$dummy [117]), .D (nx14784), .CLK (
        CLK)) ;
    mux21_ni ix14785 (.Y (nx14784), .A0 (Din[6]), .A1 (Mem_30__6), .S0 (nx17595)
             ) ;
    dff reg_Mem_11__6 (.Q (Mem_11__6), .QB (\$dummy [118]), .D (nx14774), .CLK (
        CLK)) ;
    mux21_ni ix14775 (.Y (nx14774), .A0 (Mem_11__6), .A1 (Din[6]), .S0 (nx17397)
             ) ;
    aoi22 ix16627 (.Y (nx16626), .A0 (Mem_26__6), .A1 (nx17705), .B0 (Mem_25__6)
          , .B1 (nx17701)) ;
    dff reg_Mem_26__6 (.Q (Mem_26__6), .QB (\$dummy [119]), .D (nx14764), .CLK (
        CLK)) ;
    mux21_ni ix14765 (.Y (nx14764), .A0 (Din[6]), .A1 (Mem_26__6), .S0 (nx17599)
             ) ;
    dff reg_Mem_25__6 (.Q (Mem_25__6), .QB (\$dummy [120]), .D (nx14754), .CLK (
        CLK)) ;
    mux21_ni ix14755 (.Y (nx14754), .A0 (Mem_25__6), .A1 (Din[6]), .S0 (nx17393)
             ) ;
    aoi22 ix16635 (.Y (nx16634), .A0 (Mem_27__6), .A1 (nx17697), .B0 (Mem_2__6)
          , .B1 (nx17389)) ;
    dff reg_Mem_27__6 (.Q (Mem_27__6), .QB (\$dummy [121]), .D (nx14744), .CLK (
        CLK)) ;
    mux21_ni ix14745 (.Y (nx14744), .A0 (Din[6]), .A1 (Mem_27__6), .S0 (nx17603)
             ) ;
    oai22 ix3951 (.Y (nx3950), .A0 (nx15548), .A1 (nx16000), .B0 (nx15535), .B1 (
          nx17607)) ;
    oai22 ix3945 (.Y (nx3944), .A0 (nx15527), .A1 (nx16006), .B0 (nx15540), .B1 (
          nx16008)) ;
    oai221 ix3939 (.Y (nx3938), .A0 (nx15543), .A1 (nx16011), .B0 (nx16642), .B1 (
           nx16022), .C0 (nx16646)) ;
    dff reg_Mem_21__6 (.Q (Mem_21__6), .QB (nx16642), .D (nx14714), .CLK (CLK)
        ) ;
    aoi22 ix16647 (.Y (nx16646), .A0 (Mem_20__6), .A1 (nx1674), .B0 (Mem_22__6)
          , .B1 (nx1626)) ;
    dff reg_Mem_20__6 (.Q (Mem_20__6), .QB (nx16650), .D (nx14734), .CLK (CLK)
        ) ;
    dff reg_Mem_22__6 (.Q (Mem_22__6), .QB (\$dummy [122]), .D (nx14724), .CLK (
        CLK)) ;
    mux21_ni ix14725 (.Y (nx14724), .A0 (Mem_22__6), .A1 (Din[6]), .S0 (nx17381)
             ) ;
    nand04 ix4419 (.Y (Dout[23]), .A0 (nx16655), .A1 (nx16666), .A2 (nx16683), .A3 (
           nx16714)) ;
    aoi222 ix16656 (.Y (nx16655), .A0 (Mem_28__7), .A1 (nx17443), .B0 (Mem_24__7
           ), .B1 (nx2576), .C0 (Mem_17__7), .C1 (nx2614)) ;
    dff reg_Mem_28__7 (.Q (Mem_28__7), .QB (nx16659), .D (nx15144), .CLK (CLK)
        ) ;
    dff reg_Mem_24__7 (.Q (Mem_24__7), .QB (\$dummy [123]), .D (nx15154), .CLK (
        CLK)) ;
    mux21_ni ix15155 (.Y (nx15154), .A0 (Din[7]), .A1 (Mem_24__7), .S0 (nx17571)
             ) ;
    dff reg_Mem_17__7 (.Q (Mem_17__7), .QB (nx16665), .D (nx15164), .CLK (CLK)
        ) ;
    aoi221 ix16667 (.Y (nx16666), .A0 (Mem_16__7), .A1 (nx17739), .B0 (Mem_23__7
           ), .B1 (nx17735), .C0 (nx4364)) ;
    dff reg_Mem_16__7 (.Q (Mem_16__7), .QB (nx16670), .D (nx15134), .CLK (CLK)
        ) ;
    dff reg_Mem_23__7 (.Q (Mem_23__7), .QB (\$dummy [124]), .D (nx15124), .CLK (
        CLK)) ;
    mux21_ni ix15125 (.Y (nx15124), .A0 (Mem_23__7), .A1 (Din[7]), .S0 (nx17435)
             ) ;
    oai22 ix4365 (.Y (nx4364), .A0 (nx16675), .A1 (nx15821), .B0 (nx16679), .B1 (
          nx17585)) ;
    dff reg_Mem_14__7 (.Q (Mem_14__7), .QB (nx16675), .D (nx15114), .CLK (CLK)
        ) ;
    dff reg_Mem_12__7 (.Q (Mem_12__7), .QB (nx16679), .D (nx15104), .CLK (CLK)
        ) ;
    and04 ix16684 (.Y (nx16683), .A0 (nx16685), .A1 (nx16693), .A2 (nx16701), .A3 (
          nx16706)) ;
    aoi22 ix16686 (.Y (nx16685), .A0 (Mem_19__7), .A1 (nx17731), .B0 (Mem_13__7)
          , .B1 (nx2336)) ;
    dff reg_Mem_19__7 (.Q (Mem_19__7), .QB (nx16689), .D (nx15084), .CLK (CLK)
        ) ;
    dff reg_Mem_13__7 (.Q (Mem_13__7), .QB (\$dummy [125]), .D (nx15094), .CLK (
        CLK)) ;
    mux21_ni ix15095 (.Y (nx15094), .A0 (Mem_13__7), .A1 (Din[7]), .S0 (nx17431)
             ) ;
    aoi22 ix16694 (.Y (nx16693), .A0 (Mem_10__7), .A1 (nx17727), .B0 (Mem_15__7)
          , .B1 (nx2220)) ;
    dff reg_Mem_10__7 (.Q (Mem_10__7), .QB (\$dummy [126]), .D (nx15074), .CLK (
        CLK)) ;
    mux21_ni ix15075 (.Y (nx15074), .A0 (Din[7]), .A1 (Mem_10__7), .S0 (nx17589)
             ) ;
    dff reg_Mem_15__7 (.Q (Mem_15__7), .QB (\$dummy [127]), .D (nx15064), .CLK (
        CLK)) ;
    mux21_ni ix15065 (.Y (nx15064), .A0 (Mem_15__7), .A1 (Din[7]), .S0 (nx17423)
             ) ;
    aoi22 ix16702 (.Y (nx16701), .A0 (Mem_9__7), .A1 (nx17723), .B0 (Mem_8__7), 
          .B1 (nx17719)) ;
    dff reg_Mem_9__7 (.Q (Mem_9__7), .QB (\$dummy [128]), .D (nx15054), .CLK (
        CLK)) ;
    mux21_ni ix15055 (.Y (nx15054), .A0 (Mem_9__7), .A1 (Din[7]), .S0 (nx17419)
             ) ;
    aoi22 ix16707 (.Y (nx16706), .A0 (Mem_29__7), .A1 (nx17711), .B0 (Mem_18__7)
          , .B1 (nx17715)) ;
    dff reg_Mem_29__7 (.Q (Mem_29__7), .QB (nx16710), .D (nx15034), .CLK (CLK)
        ) ;
    dff reg_Mem_18__7 (.Q (Mem_18__7), .QB (\$dummy [129]), .D (nx15044), .CLK (
        CLK)) ;
    mux21_ni ix15045 (.Y (nx15044), .A0 (Mem_18__7), .A1 (Din[7]), .S0 (nx17415)
             ) ;
    nor04 ix16715 (.Y (nx16714), .A0 (nx4272), .A1 (nx4206), .A2 (nx4200), .A3 (
          nx4194)) ;
    nand03 ix4273 (.Y (nx4272), .A0 (nx16717), .A1 (nx16728), .A2 (nx16736)) ;
    aoi222 ix16718 (.Y (nx16717), .A0 (Mem_31__7), .A1 (nx17407), .B0 (Mem_30__7
           ), .B1 (nx1972), .C0 (Mem_11__7), .C1 (nx1916)) ;
    dff reg_Mem_31__7 (.Q (Mem_31__7), .QB (nx16721), .D (nx15024), .CLK (CLK)
        ) ;
    dff reg_Mem_30__7 (.Q (Mem_30__7), .QB (\$dummy [130]), .D (nx15014), .CLK (
        CLK)) ;
    mux21_ni ix15015 (.Y (nx15014), .A0 (Din[7]), .A1 (Mem_30__7), .S0 (nx17597)
             ) ;
    dff reg_Mem_11__7 (.Q (Mem_11__7), .QB (\$dummy [131]), .D (nx15004), .CLK (
        CLK)) ;
    mux21_ni ix15005 (.Y (nx15004), .A0 (Mem_11__7), .A1 (Din[7]), .S0 (nx17399)
             ) ;
    aoi22 ix16729 (.Y (nx16728), .A0 (Mem_26__7), .A1 (nx17707), .B0 (Mem_25__7)
          , .B1 (nx17703)) ;
    dff reg_Mem_26__7 (.Q (Mem_26__7), .QB (\$dummy [132]), .D (nx14994), .CLK (
        CLK)) ;
    mux21_ni ix14995 (.Y (nx14994), .A0 (Din[7]), .A1 (Mem_26__7), .S0 (nx17601)
             ) ;
    dff reg_Mem_25__7 (.Q (Mem_25__7), .QB (\$dummy [133]), .D (nx14984), .CLK (
        CLK)) ;
    mux21_ni ix14985 (.Y (nx14984), .A0 (Mem_25__7), .A1 (Din[7]), .S0 (nx17395)
             ) ;
    aoi22 ix16737 (.Y (nx16736), .A0 (Mem_27__7), .A1 (nx17699), .B0 (Mem_2__7)
          , .B1 (nx17391)) ;
    dff reg_Mem_27__7 (.Q (Mem_27__7), .QB (\$dummy [134]), .D (nx14974), .CLK (
        CLK)) ;
    mux21_ni ix14975 (.Y (nx14974), .A0 (Din[7]), .A1 (Mem_27__7), .S0 (nx17605)
             ) ;
    oai22 ix4207 (.Y (nx4206), .A0 (nx15581), .A1 (nx16000), .B0 (nx15568), .B1 (
          nx17609)) ;
    oai22 ix4201 (.Y (nx4200), .A0 (nx15560), .A1 (nx16006), .B0 (nx15573), .B1 (
          nx16008)) ;
    oai221 ix4195 (.Y (nx4194), .A0 (nx15576), .A1 (nx16011), .B0 (nx16744), .B1 (
           nx16022), .C0 (nx16748)) ;
    dff reg_Mem_21__7 (.Q (Mem_21__7), .QB (nx16744), .D (nx14944), .CLK (CLK)
        ) ;
    aoi22 ix16749 (.Y (nx16748), .A0 (Mem_20__7), .A1 (nx1674), .B0 (Mem_22__7)
          , .B1 (nx1626)) ;
    dff reg_Mem_20__7 (.Q (Mem_20__7), .QB (nx16752), .D (nx14964), .CLK (CLK)
        ) ;
    dff reg_Mem_22__7 (.Q (Mem_22__7), .QB (\$dummy [135]), .D (nx14954), .CLK (
        CLK)) ;
    mux21_ni ix14955 (.Y (nx14954), .A0 (Mem_22__7), .A1 (Din[7]), .S0 (nx17383)
             ) ;
    nand04 ix4689 (.Y (Dout[24]), .A0 (nx16757), .A1 (nx16786), .A2 (nx16800), .A3 (
           nx16823)) ;
    aoi222 ix16758 (.Y (nx16757), .A0 (Mem_13__0), .A1 (nx17477), .B0 (Mem_8__0)
           , .B1 (nx17845), .C0 (Mem_28__0), .C1 (nx17473)) ;
    nor02_2x ix4677 (.Y (nx4676), .A0 (nx16760), .A1 (nx16762)) ;
    nand02 ix16761 (.Y (nx16760), .A0 (nx15208), .A1 (Address[6])) ;
    nand03 ix16763 (.Y (nx16762), .A0 (nx16764), .A1 (nx4428), .A2 (nx4436)) ;
    xnor2 ix16765 (.Y (nx16764), .A0 (nx4430), .A1 (Address[9])) ;
    oai21 ix16768 (.Y (nx16767), .A0 (Address[5]), .A1 (Address[6]), .B0 (
          Address[7])) ;
    nor02_2x ix16771 (.Y (nx16770), .A0 (Address[5]), .A1 (Address[6])) ;
    xnor2_2x ix4437 (.Y (nx4436), .A0 (Address[8]), .A1 (nx17615)) ;
    nand03 ix16777 (.Y (nx16776), .A0 (nx16764), .A1 (nx17617), .A2 (nx4436)) ;
    oai21 ix16779 (.Y (nx16778), .A0 (nx4420), .A1 (Address[7]), .B0 (nx17615)
          ) ;
    and02 ix4673 (.Y (nx4672), .A0 (nx17743), .A1 (nx4514)) ;
    nor03_2x ix4515 (.Y (nx4514), .A0 (nx16764), .A1 (nx17617), .A2 (nx16784)) ;
    aoi221 ix16787 (.Y (nx16786), .A0 (Mem_12__0), .A1 (nx17767), .B0 (Mem_21__0
           ), .B1 (nx17771), .C0 (nx4664)) ;
    oai22 ix4665 (.Y (nx4664), .A0 (nx15916), .A1 (nx16794), .B0 (nx16033), .B1 (
          nx17619)) ;
    nand02 ix16795 (.Y (nx16794), .A0 (nx4482), .A1 (nx4514)) ;
    nand02 ix16798 (.Y (nx16797), .A0 (nx17743), .A1 (nx4584)) ;
    nor03_2x ix4585 (.Y (nx4584), .A0 (nx16764), .A1 (nx17617), .A2 (nx4436)) ;
    and03 ix16801 (.Y (nx16800), .A0 (nx16802), .A1 (nx16811), .A2 (nx16817)) ;
    aoi222 ix16803 (.Y (nx16802), .A0 (Mem_14__0), .A1 (nx17465), .B0 (Mem_18__0
           ), .B1 (nx17843), .C0 (Mem_22__0), .C1 (nx17841)) ;
    nor02_2x ix4633 (.Y (nx4632), .A0 (nx17623), .A1 (nx16762)) ;
    nand02 ix16806 (.Y (nx16805), .A0 (Address[5]), .A1 (Address[6])) ;
    aoi22 ix16812 (.Y (nx16811), .A0 (Mem_9__0), .A1 (nx4620), .B0 (Mem_7__0), .B1 (
          nx4616)) ;
    nor02_2x ix4621 (.Y (nx4620), .A0 (nx16760), .A1 (nx16776)) ;
    and02 ix4617 (.Y (nx4616), .A0 (nx17741), .A1 (nx4498)) ;
    nor02_2x ix4455 (.Y (nx4454), .A0 (Address[5]), .A1 (Address[6])) ;
    nor03_2x ix4499 (.Y (nx4498), .A0 (nx4444), .A1 (nx17617), .A2 (nx4436)) ;
    aoi22 ix16818 (.Y (nx16817), .A0 (Mem_10__0), .A1 (nx4610), .B0 (Mem_11__0)
          , .B1 (nx17763)) ;
    nor02_2x ix4611 (.Y (nx4610), .A0 (nx17623), .A1 (nx16776)) ;
    nor04 ix16824 (.Y (nx16823), .A0 (nx4594), .A1 (nx4540), .A2 (nx4504), .A3 (
          nx4476)) ;
    nand03 ix4595 (.Y (nx4594), .A0 (nx16826), .A1 (nx16833), .A2 (nx16839)) ;
    aoi222 ix16827 (.Y (nx16826), .A0 (Mem_15__0), .A1 (nx17455), .B0 (Mem_23__0
           ), .B1 (nx17459), .C0 (Mem_6__0), .C1 (nx17839)) ;
    and02 ix4587 (.Y (nx4586), .A0 (nx17741), .A1 (nx4584)) ;
    aoi22 ix16834 (.Y (nx16833), .A0 (Mem_25__0), .A1 (nx4558), .B0 (Mem_24__0)
          , .B1 (nx17759)) ;
    nor02_2x ix4559 (.Y (nx4558), .A0 (nx16760), .A1 (nx16836)) ;
    nand03 ix16837 (.Y (nx16836), .A0 (nx4444), .A1 (nx17617), .A2 (nx4436)) ;
    aoi22 ix16840 (.Y (nx16839), .A0 (Mem_30__0), .A1 (nx17755), .B0 (Mem_27__0)
          , .B1 (nx17751)) ;
    oai221 ix4541 (.Y (nx4540), .A0 (nx15946), .A1 (nx17625), .B0 (nx15786), .B1 (
           nx17627), .C0 (nx16851)) ;
    nand02 ix16847 (.Y (nx16846), .A0 (nx17741), .A1 (nx4514)) ;
    nand02 ix16849 (.Y (nx16848), .A0 (nx17743), .A1 (nx4470)) ;
    nor03_2x ix4471 (.Y (nx4470), .A0 (nx16764), .A1 (nx4428), .A2 (nx4436)) ;
    aoi22 ix16852 (.Y (nx16851), .A0 (Mem_26__0), .A1 (nx4530), .B0 (Mem_5__0), 
          .B1 (nx17747)) ;
    nor02_2x ix4531 (.Y (nx4530), .A0 (nx16805), .A1 (nx16836)) ;
    oai22 ix4505 (.Y (nx4504), .A0 (nx15244), .A1 (nx16856), .B0 (nx15767), .B1 (
          nx17629)) ;
    nand02 ix16857 (.Y (nx16856), .A0 (nx17743), .A1 (nx4498)) ;
    nand02 ix16859 (.Y (nx16858), .A0 (nx4482), .A1 (nx4470)) ;
    oai22 ix4477 (.Y (nx4476), .A0 (nx15291), .A1 (nx16861), .B0 (nx15848), .B1 (
          nx17633)) ;
    nand04 ix16862 (.Y (nx16861), .A0 (nx17617), .A1 (nx16784), .A2 (nx16764), .A3 (
           nx17741)) ;
    nand02 ix16864 (.Y (nx16863), .A0 (nx17741), .A1 (nx4470)) ;
    nand04 ix4803 (.Y (Dout[25]), .A0 (nx16866), .A1 (nx16868), .A2 (nx16871), .A3 (
           nx16879)) ;
    aoi222 ix16867 (.Y (nx16866), .A0 (Mem_13__1), .A1 (nx17477), .B0 (Mem_8__1)
           , .B1 (nx17845), .C0 (Mem_28__1), .C1 (nx17473)) ;
    aoi221 ix16869 (.Y (nx16868), .A0 (Mem_12__1), .A1 (nx17767), .B0 (Mem_21__1
           ), .B1 (nx17771), .C0 (nx4784)) ;
    oai22 ix4785 (.Y (nx4784), .A0 (nx16098), .A1 (nx16794), .B0 (nx16140), .B1 (
          nx17619)) ;
    and03 ix16872 (.Y (nx16871), .A0 (nx16873), .A1 (nx16875), .A2 (nx16877)) ;
    aoi222 ix16874 (.Y (nx16873), .A0 (Mem_14__1), .A1 (nx17465), .B0 (Mem_18__1
           ), .B1 (nx17843), .C0 (Mem_22__1), .C1 (nx17841)) ;
    aoi22 ix16876 (.Y (nx16875), .A0 (Mem_9__1), .A1 (nx4620), .B0 (Mem_7__1), .B1 (
          nx4616)) ;
    aoi22 ix16878 (.Y (nx16877), .A0 (Mem_10__1), .A1 (nx4610), .B0 (Mem_11__1)
          , .B1 (nx17763)) ;
    nor04 ix16880 (.Y (nx16879), .A0 (nx4744), .A1 (nx4716), .A2 (nx4700), .A3 (
          nx4694)) ;
    nand03 ix4745 (.Y (nx4744), .A0 (nx16882), .A1 (nx16884), .A2 (nx16886)) ;
    aoi222 ix16883 (.Y (nx16882), .A0 (Mem_15__1), .A1 (nx17455), .B0 (Mem_23__1
           ), .B1 (nx17459), .C0 (Mem_6__1), .C1 (nx17839)) ;
    aoi22 ix16885 (.Y (nx16884), .A0 (Mem_25__1), .A1 (nx4558), .B0 (Mem_24__1)
          , .B1 (nx17759)) ;
    aoi22 ix16887 (.Y (nx16886), .A0 (Mem_30__1), .A1 (nx17755), .B0 (Mem_27__1)
          , .B1 (nx17751)) ;
    oai221 ix4717 (.Y (nx4716), .A0 (nx16109), .A1 (nx17625), .B0 (nx16058), .B1 (
           nx17627), .C0 (nx16889)) ;
    aoi22 ix16890 (.Y (nx16889), .A0 (Mem_26__1), .A1 (nx4530), .B0 (Mem_5__1), 
          .B1 (nx17747)) ;
    oai22 ix4701 (.Y (nx4700), .A0 (nx15362), .A1 (nx16856), .B0 (nx16053), .B1 (
          nx17629)) ;
    oai22 ix4695 (.Y (nx4694), .A0 (nx15375), .A1 (nx16861), .B0 (nx16077), .B1 (
          nx17633)) ;
    nand04 ix4917 (.Y (Dout[26]), .A0 (nx16894), .A1 (nx16896), .A2 (nx16899), .A3 (
           nx16907)) ;
    aoi222 ix16895 (.Y (nx16894), .A0 (Mem_13__2), .A1 (nx17477), .B0 (Mem_8__2)
           , .B1 (nx17845), .C0 (Mem_28__2), .C1 (nx17473)) ;
    aoi221 ix16897 (.Y (nx16896), .A0 (Mem_12__2), .A1 (nx17767), .B0 (Mem_21__2
           ), .B1 (nx17771), .C0 (nx4898)) ;
    oai22 ix4899 (.Y (nx4898), .A0 (nx16200), .A1 (nx16794), .B0 (nx16242), .B1 (
          nx17619)) ;
    and03 ix16900 (.Y (nx16899), .A0 (nx16901), .A1 (nx16903), .A2 (nx16905)) ;
    aoi222 ix16902 (.Y (nx16901), .A0 (Mem_14__2), .A1 (nx17465), .B0 (Mem_18__2
           ), .B1 (nx17843), .C0 (Mem_22__2), .C1 (nx17841)) ;
    aoi22 ix16904 (.Y (nx16903), .A0 (Mem_9__2), .A1 (nx4620), .B0 (Mem_7__2), .B1 (
          nx4616)) ;
    aoi22 ix16906 (.Y (nx16905), .A0 (Mem_10__2), .A1 (nx4610), .B0 (Mem_11__2)
          , .B1 (nx17763)) ;
    nor04 ix16908 (.Y (nx16907), .A0 (nx4858), .A1 (nx4830), .A2 (nx4814), .A3 (
          nx4808)) ;
    nand03 ix4859 (.Y (nx4858), .A0 (nx16910), .A1 (nx16912), .A2 (nx16914)) ;
    aoi222 ix16911 (.Y (nx16910), .A0 (Mem_15__2), .A1 (nx17455), .B0 (Mem_23__2
           ), .B1 (nx17459), .C0 (Mem_6__2), .C1 (nx17839)) ;
    aoi22 ix16913 (.Y (nx16912), .A0 (Mem_25__2), .A1 (nx4558), .B0 (Mem_24__2)
          , .B1 (nx17759)) ;
    aoi22 ix16915 (.Y (nx16914), .A0 (Mem_30__2), .A1 (nx17755), .B0 (Mem_27__2)
          , .B1 (nx17751)) ;
    oai221 ix4831 (.Y (nx4830), .A0 (nx16211), .A1 (nx17625), .B0 (nx16160), .B1 (
           nx17627), .C0 (nx16917)) ;
    aoi22 ix16918 (.Y (nx16917), .A0 (Mem_26__2), .A1 (nx4530), .B0 (Mem_5__2), 
          .B1 (nx17747)) ;
    oai22 ix4815 (.Y (nx4814), .A0 (nx15395), .A1 (nx16856), .B0 (nx16155), .B1 (
          nx17629)) ;
    oai22 ix4809 (.Y (nx4808), .A0 (nx15408), .A1 (nx16861), .B0 (nx16179), .B1 (
          nx17633)) ;
    nand04 ix5031 (.Y (Dout[27]), .A0 (nx16922), .A1 (nx16924), .A2 (nx16927), .A3 (
           nx16935)) ;
    aoi222 ix16923 (.Y (nx16922), .A0 (Mem_13__3), .A1 (nx17477), .B0 (Mem_8__3)
           , .B1 (nx17845), .C0 (Mem_28__3), .C1 (nx17473)) ;
    aoi221 ix16925 (.Y (nx16924), .A0 (Mem_12__3), .A1 (nx17767), .B0 (Mem_21__3
           ), .B1 (nx17771), .C0 (nx5012)) ;
    oai22 ix5013 (.Y (nx5012), .A0 (nx16302), .A1 (nx16794), .B0 (nx16344), .B1 (
          nx17619)) ;
    and03 ix16928 (.Y (nx16927), .A0 (nx16929), .A1 (nx16931), .A2 (nx16933)) ;
    aoi222 ix16930 (.Y (nx16929), .A0 (Mem_14__3), .A1 (nx17465), .B0 (Mem_18__3
           ), .B1 (nx17843), .C0 (Mem_22__3), .C1 (nx17841)) ;
    aoi22 ix16932 (.Y (nx16931), .A0 (Mem_9__3), .A1 (nx4620), .B0 (Mem_7__3), .B1 (
          nx4616)) ;
    aoi22 ix16934 (.Y (nx16933), .A0 (Mem_10__3), .A1 (nx4610), .B0 (Mem_11__3)
          , .B1 (nx17763)) ;
    nor04 ix16936 (.Y (nx16935), .A0 (nx4972), .A1 (nx4944), .A2 (nx4928), .A3 (
          nx4922)) ;
    nand03 ix4973 (.Y (nx4972), .A0 (nx16938), .A1 (nx16940), .A2 (nx16942)) ;
    aoi222 ix16939 (.Y (nx16938), .A0 (Mem_15__3), .A1 (nx17455), .B0 (Mem_23__3
           ), .B1 (nx17459), .C0 (Mem_6__3), .C1 (nx17839)) ;
    aoi22 ix16941 (.Y (nx16940), .A0 (Mem_25__3), .A1 (nx4558), .B0 (Mem_24__3)
          , .B1 (nx17759)) ;
    aoi22 ix16943 (.Y (nx16942), .A0 (Mem_30__3), .A1 (nx17755), .B0 (Mem_27__3)
          , .B1 (nx17751)) ;
    oai221 ix4945 (.Y (nx4944), .A0 (nx16313), .A1 (nx17625), .B0 (nx16262), .B1 (
           nx17627), .C0 (nx16945)) ;
    aoi22 ix16946 (.Y (nx16945), .A0 (Mem_26__3), .A1 (nx4530), .B0 (Mem_5__3), 
          .B1 (nx17747)) ;
    oai22 ix4929 (.Y (nx4928), .A0 (nx15428), .A1 (nx16856), .B0 (nx16257), .B1 (
          nx17629)) ;
    oai22 ix4923 (.Y (nx4922), .A0 (nx15441), .A1 (nx16861), .B0 (nx16281), .B1 (
          nx17633)) ;
    nand04 ix5145 (.Y (Dout[28]), .A0 (nx16950), .A1 (nx16952), .A2 (nx16955), .A3 (
           nx16963)) ;
    aoi222 ix16951 (.Y (nx16950), .A0 (Mem_13__4), .A1 (nx17477), .B0 (Mem_8__4)
           , .B1 (nx17845), .C0 (Mem_28__4), .C1 (nx17473)) ;
    aoi221 ix16953 (.Y (nx16952), .A0 (Mem_12__4), .A1 (nx17767), .B0 (Mem_21__4
           ), .B1 (nx17771), .C0 (nx5126)) ;
    oai22 ix5127 (.Y (nx5126), .A0 (nx16404), .A1 (nx16794), .B0 (nx16446), .B1 (
          nx17619)) ;
    and03 ix16956 (.Y (nx16955), .A0 (nx16957), .A1 (nx16959), .A2 (nx16961)) ;
    aoi222 ix16958 (.Y (nx16957), .A0 (Mem_14__4), .A1 (nx17465), .B0 (Mem_18__4
           ), .B1 (nx17843), .C0 (Mem_22__4), .C1 (nx17841)) ;
    aoi22 ix16960 (.Y (nx16959), .A0 (Mem_9__4), .A1 (nx4620), .B0 (Mem_7__4), .B1 (
          nx4616)) ;
    aoi22 ix16962 (.Y (nx16961), .A0 (Mem_10__4), .A1 (nx4610), .B0 (Mem_11__4)
          , .B1 (nx17763)) ;
    nor04 ix16964 (.Y (nx16963), .A0 (nx5086), .A1 (nx5058), .A2 (nx5042), .A3 (
          nx5036)) ;
    nand03 ix5087 (.Y (nx5086), .A0 (nx16966), .A1 (nx16968), .A2 (nx16970)) ;
    aoi222 ix16967 (.Y (nx16966), .A0 (Mem_15__4), .A1 (nx17455), .B0 (Mem_23__4
           ), .B1 (nx17459), .C0 (Mem_6__4), .C1 (nx17839)) ;
    aoi22 ix16969 (.Y (nx16968), .A0 (Mem_25__4), .A1 (nx4558), .B0 (Mem_24__4)
          , .B1 (nx17759)) ;
    aoi22 ix16971 (.Y (nx16970), .A0 (Mem_30__4), .A1 (nx17755), .B0 (Mem_27__4)
          , .B1 (nx17751)) ;
    oai221 ix5059 (.Y (nx5058), .A0 (nx16415), .A1 (nx17625), .B0 (nx16364), .B1 (
           nx17627), .C0 (nx16973)) ;
    aoi22 ix16974 (.Y (nx16973), .A0 (Mem_26__4), .A1 (nx4530), .B0 (Mem_5__4), 
          .B1 (nx17747)) ;
    oai22 ix5043 (.Y (nx5042), .A0 (nx15461), .A1 (nx16856), .B0 (nx16359), .B1 (
          nx17629)) ;
    oai22 ix5037 (.Y (nx5036), .A0 (nx15474), .A1 (nx16861), .B0 (nx16383), .B1 (
          nx17633)) ;
    nand04 ix5259 (.Y (Dout[29]), .A0 (nx16978), .A1 (nx16980), .A2 (nx16983), .A3 (
           nx16991)) ;
    aoi222 ix16979 (.Y (nx16978), .A0 (Mem_13__5), .A1 (nx17477), .B0 (Mem_8__5)
           , .B1 (nx17845), .C0 (Mem_28__5), .C1 (nx17473)) ;
    aoi221 ix16981 (.Y (nx16980), .A0 (Mem_12__5), .A1 (nx17767), .B0 (Mem_21__5
           ), .B1 (nx17771), .C0 (nx5240)) ;
    oai22 ix5241 (.Y (nx5240), .A0 (nx16506), .A1 (nx16794), .B0 (nx16548), .B1 (
          nx17619)) ;
    and03 ix16984 (.Y (nx16983), .A0 (nx16985), .A1 (nx16987), .A2 (nx16989)) ;
    aoi222 ix16986 (.Y (nx16985), .A0 (Mem_14__5), .A1 (nx17465), .B0 (Mem_18__5
           ), .B1 (nx17843), .C0 (Mem_22__5), .C1 (nx17841)) ;
    aoi22 ix16988 (.Y (nx16987), .A0 (Mem_9__5), .A1 (nx4620), .B0 (Mem_7__5), .B1 (
          nx4616)) ;
    aoi22 ix16990 (.Y (nx16989), .A0 (Mem_10__5), .A1 (nx4610), .B0 (Mem_11__5)
          , .B1 (nx17763)) ;
    nor04 ix16992 (.Y (nx16991), .A0 (nx5200), .A1 (nx5172), .A2 (nx5156), .A3 (
          nx5150)) ;
    nand03 ix5201 (.Y (nx5200), .A0 (nx16994), .A1 (nx16996), .A2 (nx16998)) ;
    aoi222 ix16995 (.Y (nx16994), .A0 (Mem_15__5), .A1 (nx17455), .B0 (Mem_23__5
           ), .B1 (nx17459), .C0 (Mem_6__5), .C1 (nx17839)) ;
    aoi22 ix16997 (.Y (nx16996), .A0 (Mem_25__5), .A1 (nx4558), .B0 (Mem_24__5)
          , .B1 (nx17759)) ;
    aoi22 ix16999 (.Y (nx16998), .A0 (Mem_30__5), .A1 (nx17755), .B0 (Mem_27__5)
          , .B1 (nx17751)) ;
    oai221 ix5173 (.Y (nx5172), .A0 (nx16517), .A1 (nx16846), .B0 (nx16466), .B1 (
           nx16848), .C0 (nx17001)) ;
    aoi22 ix17002 (.Y (nx17001), .A0 (Mem_26__5), .A1 (nx4530), .B0 (Mem_5__5), 
          .B1 (nx17747)) ;
    oai22 ix5157 (.Y (nx5156), .A0 (nx15494), .A1 (nx16856), .B0 (nx16461), .B1 (
          nx17629)) ;
    oai22 ix5151 (.Y (nx5150), .A0 (nx15507), .A1 (nx16861), .B0 (nx16485), .B1 (
          nx17633)) ;
    nand04 ix5373 (.Y (Dout[30]), .A0 (nx17006), .A1 (nx17008), .A2 (nx17011), .A3 (
           nx17019)) ;
    aoi222 ix17007 (.Y (nx17006), .A0 (Mem_13__6), .A1 (nx17477), .B0 (Mem_8__6)
           , .B1 (nx4668), .C0 (Mem_28__6), .C1 (nx17473)) ;
    aoi221 ix17009 (.Y (nx17008), .A0 (Mem_12__6), .A1 (nx17767), .B0 (Mem_21__6
           ), .B1 (nx17771), .C0 (nx5354)) ;
    oai22 ix5355 (.Y (nx5354), .A0 (nx16608), .A1 (nx16794), .B0 (nx16650), .B1 (
          nx17619)) ;
    and03 ix17012 (.Y (nx17011), .A0 (nx17013), .A1 (nx17015), .A2 (nx17017)) ;
    aoi222 ix17014 (.Y (nx17013), .A0 (Mem_14__6), .A1 (nx17465), .B0 (Mem_18__6
           ), .B1 (nx4636), .C0 (Mem_22__6), .C1 (nx4628)) ;
    aoi22 ix17016 (.Y (nx17015), .A0 (Mem_9__6), .A1 (nx4620), .B0 (Mem_7__6), .B1 (
          nx4616)) ;
    aoi22 ix17018 (.Y (nx17017), .A0 (Mem_10__6), .A1 (nx4610), .B0 (Mem_11__6)
          , .B1 (nx17763)) ;
    nor04 ix17020 (.Y (nx17019), .A0 (nx5314), .A1 (nx5286), .A2 (nx5270), .A3 (
          nx5264)) ;
    nand03 ix5315 (.Y (nx5314), .A0 (nx17022), .A1 (nx17024), .A2 (nx17026)) ;
    aoi222 ix17023 (.Y (nx17022), .A0 (Mem_15__6), .A1 (nx17455), .B0 (Mem_23__6
           ), .B1 (nx17459), .C0 (Mem_6__6), .C1 (nx4566)) ;
    aoi22 ix17025 (.Y (nx17024), .A0 (Mem_25__6), .A1 (nx4558), .B0 (Mem_24__6)
          , .B1 (nx17759)) ;
    aoi22 ix17027 (.Y (nx17026), .A0 (Mem_30__6), .A1 (nx17755), .B0 (Mem_27__6)
          , .B1 (nx17751)) ;
    oai221 ix5287 (.Y (nx5286), .A0 (nx16619), .A1 (nx16846), .B0 (nx16568), .B1 (
           nx16848), .C0 (nx17029)) ;
    aoi22 ix17030 (.Y (nx17029), .A0 (Mem_26__6), .A1 (nx4530), .B0 (Mem_5__6), 
          .B1 (nx17747)) ;
    oai22 ix5271 (.Y (nx5270), .A0 (nx15527), .A1 (nx16856), .B0 (nx16563), .B1 (
          nx17629)) ;
    oai22 ix5265 (.Y (nx5264), .A0 (nx15540), .A1 (nx16861), .B0 (nx16587), .B1 (
          nx17633)) ;
    nand04 ix5487 (.Y (Dout[31]), .A0 (nx17034), .A1 (nx17036), .A2 (nx17039), .A3 (
           nx17047)) ;
    aoi222 ix17035 (.Y (nx17034), .A0 (Mem_13__7), .A1 (nx17479), .B0 (Mem_8__7)
           , .B1 (nx4668), .C0 (Mem_28__7), .C1 (nx17475)) ;
    aoi221 ix17037 (.Y (nx17036), .A0 (Mem_12__7), .A1 (nx17769), .B0 (Mem_21__7
           ), .B1 (nx17773), .C0 (nx5468)) ;
    oai22 ix5469 (.Y (nx5468), .A0 (nx16710), .A1 (nx16794), .B0 (nx16752), .B1 (
          nx17621)) ;
    and03 ix17040 (.Y (nx17039), .A0 (nx17041), .A1 (nx17043), .A2 (nx17045)) ;
    aoi222 ix17042 (.Y (nx17041), .A0 (Mem_14__7), .A1 (nx17467), .B0 (Mem_18__7
           ), .B1 (nx4636), .C0 (Mem_22__7), .C1 (nx4628)) ;
    aoi22 ix17044 (.Y (nx17043), .A0 (Mem_9__7), .A1 (nx4620), .B0 (Mem_7__7), .B1 (
          nx4616)) ;
    aoi22 ix17046 (.Y (nx17045), .A0 (Mem_10__7), .A1 (nx4610), .B0 (Mem_11__7)
          , .B1 (nx17765)) ;
    nor04 ix17048 (.Y (nx17047), .A0 (nx5428), .A1 (nx5400), .A2 (nx5384), .A3 (
          nx5378)) ;
    nand03 ix5429 (.Y (nx5428), .A0 (nx17050), .A1 (nx17052), .A2 (nx17054)) ;
    aoi222 ix17051 (.Y (nx17050), .A0 (Mem_15__7), .A1 (nx17457), .B0 (Mem_23__7
           ), .B1 (nx17461), .C0 (Mem_6__7), .C1 (nx4566)) ;
    aoi22 ix17053 (.Y (nx17052), .A0 (Mem_25__7), .A1 (nx4558), .B0 (Mem_24__7)
          , .B1 (nx17761)) ;
    aoi22 ix17055 (.Y (nx17054), .A0 (Mem_30__7), .A1 (nx17757), .B0 (Mem_27__7)
          , .B1 (nx17753)) ;
    oai221 ix5401 (.Y (nx5400), .A0 (nx16721), .A1 (nx16846), .B0 (nx16670), .B1 (
           nx16848), .C0 (nx17057)) ;
    aoi22 ix17058 (.Y (nx17057), .A0 (Mem_26__7), .A1 (nx4530), .B0 (Mem_5__7), 
          .B1 (nx17749)) ;
    oai22 ix5385 (.Y (nx5384), .A0 (nx15560), .A1 (nx16856), .B0 (nx16665), .B1 (
          nx17631)) ;
    oai22 ix5379 (.Y (nx5378), .A0 (nx15573), .A1 (nx16861), .B0 (nx16689), .B1 (
          nx17635)) ;
    nand04 ix5725 (.Y (Dout[32]), .A0 (nx17062), .A1 (nx17118), .A2 (nx17134), .A3 (
           nx17143)) ;
    and04 ix17063 (.Y (nx17062), .A0 (nx17064), .A1 (nx17078), .A2 (nx17096), .A3 (
          nx17103)) ;
    aoi222 ix17065 (.Y (nx17064), .A0 (Mem_11__0), .A1 (nx17529), .B0 (Mem_15__0
           ), .B1 (nx17853), .C0 (Mem_8__0), .C1 (nx17525)) ;
    oai21 ix17070 (.Y (nx17069), .A0 (Address[2]), .A1 (Address[3]), .B0 (
          nx15798)) ;
    xnor2 ix5495 (.Y (nx5494), .A0 (Address[4]), .A1 (nx15798)) ;
    nand03 ix17073 (.Y (nx17072), .A0 (Address[0]), .A1 (Address[1]), .A2 (
           Address[2])) ;
    nand03 ix17076 (.Y (nx17075), .A0 (nx17533), .A1 (Address[1]), .A2 (
           Address[0])) ;
    nor04 ix5709 (.Y (nx5708), .A0 (nx18123), .A1 (Address[0]), .A2 (Address[1])
          , .A3 (nx17533)) ;
    aoi221 ix17079 (.Y (nx17078), .A0 (Mem_19__0), .A1 (nx17809), .B0 (Mem_22__0
           ), .B1 (nx17805), .C0 (nx5690)) ;
    nand02 ix17082 (.Y (nx17081), .A0 (nx17069), .A1 (nx5494)) ;
    oai22 ix5691 (.Y (nx5690), .A0 (nx15244), .A1 (nx17087), .B0 (nx15824), .B1 (
          nx17641)) ;
    nand02 ix17088 (.Y (nx17087), .A0 (nx5532), .A1 (nx5522)) ;
    nor03_2x ix5533 (.Y (nx5532), .A0 (Address[0]), .A1 (Address[1]), .A2 (
             Address[2])) ;
    nand02 ix17094 (.Y (nx17093), .A0 (nx17783), .A1 (nx5532)) ;
    nor02_2x ix5511 (.Y (nx5510), .A0 (nx17069), .A1 (nx5494)) ;
    aoi222 ix17097 (.Y (nx17096), .A0 (Mem_31__0), .A1 (nx17519), .B0 (Mem_23__0
           ), .B1 (nx17851), .C0 (Mem_24__0), .C1 (nx17513)) ;
    nor04 ix5665 (.Y (nx5664), .A0 (nx18135), .A1 (Address[0]), .A2 (Address[1])
          , .A3 (nx17533)) ;
    aoi221 ix17104 (.Y (nx17103), .A0 (Mem_13__0), .A1 (nx17801), .B0 (Mem_9__0)
           , .B1 (nx17797), .C0 (nx5650)) ;
    nand03 ix17107 (.Y (nx17106), .A0 (nx17535), .A1 (nx17545), .A2 (Address[0])
           ) ;
    nand03 ix17110 (.Y (nx17109), .A0 (Address[0]), .A1 (nx17545), .A2 (
           Address[2])) ;
    oai22 ix5651 (.Y (nx5650), .A0 (nx15337), .A1 (nx17112), .B0 (nx16033), .B1 (
          nx17649)) ;
    nand02 ix17113 (.Y (nx17112), .A0 (nx5640), .A1 (nx5522)) ;
    nand02 ix17116 (.Y (nx17115), .A0 (nx17787), .A1 (nx5532)) ;
    and03 ix17119 (.Y (nx17118), .A0 (nx17120), .A1 (nx17126), .A2 (nx17130)) ;
    aoi222 ix17121 (.Y (nx17120), .A0 (Mem_29__0), .A1 (nx17509), .B0 (Mem_10__0
           ), .B1 (nx17505), .C0 (Mem_25__0), .C1 (nx17849)) ;
    aoi22 ix17127 (.Y (nx17126), .A0 (Mem_18__0), .A1 (nx17495), .B0 (Mem_26__0)
          , .B1 (nx17499)) ;
    aoi22 ix17131 (.Y (nx17130), .A0 (Mem_17__0), .A1 (nx17789), .B0 (Mem_27__0)
          , .B1 (nx17793)) ;
    aoi222 ix17135 (.Y (nx17134), .A0 (Mem_21__0), .A1 (nx17489), .B0 (Mem_16__0
           ), .B1 (nx17485), .C0 (Mem_5__0), .C1 (nx17847)) ;
    nor04 ix5553 (.Y (nx5552), .A0 (nx17637), .A1 (Address[0]), .A2 (Address[1])
          , .A3 (nx17535)) ;
    aoi221 ix17144 (.Y (nx17143), .A0 (Mem_30__0), .A1 (nx17779), .B0 (Mem_14__0
           ), .B1 (nx17481), .C0 (nx5538)) ;
    nor03_2x ix5503 (.Y (nx5502), .A0 (Address[2]), .A1 (nx17547), .A2 (
             Address[0])) ;
    oai22 ix5539 (.Y (nx5538), .A0 (nx15717), .A1 (nx17149), .B0 (nx15326), .B1 (
          nx17653)) ;
    nand02 ix17150 (.Y (nx17149), .A0 (nx17775), .A1 (nx5532)) ;
    nand02 ix17153 (.Y (nx17152), .A0 (nx5522), .A1 (nx5502)) ;
    nand04 ix5835 (.Y (Dout[33]), .A0 (nx17155), .A1 (nx17167), .A2 (nx17175), .A3 (
           nx17177)) ;
    and04 ix17156 (.Y (nx17155), .A0 (nx17157), .A1 (nx17159), .A2 (nx17162), .A3 (
          nx17164)) ;
    aoi222 ix17158 (.Y (nx17157), .A0 (Mem_11__1), .A1 (nx17529), .B0 (Mem_15__1
           ), .B1 (nx17853), .C0 (Mem_8__1), .C1 (nx17525)) ;
    aoi221 ix17160 (.Y (nx17159), .A0 (Mem_19__1), .A1 (nx17809), .B0 (Mem_22__1
           ), .B1 (nx17805), .C0 (nx5810)) ;
    oai22 ix5811 (.Y (nx5810), .A0 (nx15362), .A1 (nx17087), .B0 (nx16067), .B1 (
          nx17641)) ;
    aoi222 ix17163 (.Y (nx17162), .A0 (Mem_31__1), .A1 (nx17519), .B0 (Mem_23__1
           ), .B1 (nx17851), .C0 (Mem_24__1), .C1 (nx17513)) ;
    aoi221 ix17165 (.Y (nx17164), .A0 (Mem_13__1), .A1 (nx17801), .B0 (Mem_9__1)
           , .B1 (nx17797), .C0 (nx5784)) ;
    oai22 ix5785 (.Y (nx5784), .A0 (nx15383), .A1 (nx17112), .B0 (nx16140), .B1 (
          nx17649)) ;
    and03 ix17168 (.Y (nx17167), .A0 (nx17169), .A1 (nx17171), .A2 (nx17173)) ;
    aoi222 ix17170 (.Y (nx17169), .A0 (Mem_29__1), .A1 (nx17509), .B0 (Mem_10__1
           ), .B1 (nx17505), .C0 (Mem_25__1), .C1 (nx17849)) ;
    aoi22 ix17172 (.Y (nx17171), .A0 (Mem_18__1), .A1 (nx17495), .B0 (Mem_26__1)
          , .B1 (nx17499)) ;
    aoi22 ix17174 (.Y (nx17173), .A0 (Mem_17__1), .A1 (nx17789), .B0 (Mem_27__1)
          , .B1 (nx17793)) ;
    aoi222 ix17176 (.Y (nx17175), .A0 (Mem_21__1), .A1 (nx17489), .B0 (Mem_16__1
           ), .B1 (nx17485), .C0 (Mem_5__1), .C1 (nx17847)) ;
    aoi221 ix17178 (.Y (nx17177), .A0 (Mem_30__1), .A1 (nx17779), .B0 (Mem_14__1
           ), .B1 (nx17481), .C0 (nx5736)) ;
    oai22 ix5737 (.Y (nx5736), .A0 (nx16047), .A1 (nx17149), .B0 (nx15378), .B1 (
          nx17653)) ;
    nand04 ix5945 (.Y (Dout[34]), .A0 (nx17181), .A1 (nx17193), .A2 (nx17201), .A3 (
           nx17203)) ;
    and04 ix17182 (.Y (nx17181), .A0 (nx17183), .A1 (nx17185), .A2 (nx17188), .A3 (
          nx17190)) ;
    aoi222 ix17184 (.Y (nx17183), .A0 (Mem_11__2), .A1 (nx17529), .B0 (Mem_15__2
           ), .B1 (nx17853), .C0 (Mem_8__2), .C1 (nx17525)) ;
    aoi221 ix17186 (.Y (nx17185), .A0 (Mem_19__2), .A1 (nx17809), .B0 (Mem_22__2
           ), .B1 (nx17805), .C0 (nx5920)) ;
    oai22 ix5921 (.Y (nx5920), .A0 (nx15395), .A1 (nx17087), .B0 (nx16169), .B1 (
          nx17641)) ;
    aoi222 ix17189 (.Y (nx17188), .A0 (Mem_31__2), .A1 (nx17519), .B0 (Mem_23__2
           ), .B1 (nx17851), .C0 (Mem_24__2), .C1 (nx17513)) ;
    aoi221 ix17191 (.Y (nx17190), .A0 (Mem_13__2), .A1 (nx17801), .B0 (Mem_9__2)
           , .B1 (nx17797), .C0 (nx5894)) ;
    oai22 ix5895 (.Y (nx5894), .A0 (nx15416), .A1 (nx17112), .B0 (nx16242), .B1 (
          nx17649)) ;
    and03 ix17194 (.Y (nx17193), .A0 (nx17195), .A1 (nx17197), .A2 (nx17199)) ;
    aoi222 ix17196 (.Y (nx17195), .A0 (Mem_29__2), .A1 (nx17509), .B0 (Mem_10__2
           ), .B1 (nx17505), .C0 (Mem_25__2), .C1 (nx17849)) ;
    aoi22 ix17198 (.Y (nx17197), .A0 (Mem_18__2), .A1 (nx17495), .B0 (Mem_26__2)
          , .B1 (nx17499)) ;
    aoi22 ix17200 (.Y (nx17199), .A0 (Mem_17__2), .A1 (nx17789), .B0 (Mem_27__2)
          , .B1 (nx17793)) ;
    aoi222 ix17202 (.Y (nx17201), .A0 (Mem_21__2), .A1 (nx17489), .B0 (Mem_16__2
           ), .B1 (nx17485), .C0 (Mem_5__2), .C1 (nx17847)) ;
    aoi221 ix17204 (.Y (nx17203), .A0 (Mem_30__2), .A1 (nx17779), .B0 (Mem_14__2
           ), .B1 (nx17481), .C0 (nx5846)) ;
    oai22 ix5847 (.Y (nx5846), .A0 (nx16149), .A1 (nx17149), .B0 (nx15411), .B1 (
          nx17653)) ;
    nand04 ix6055 (.Y (Dout[35]), .A0 (nx17207), .A1 (nx17219), .A2 (nx17227), .A3 (
           nx17229)) ;
    and04 ix17208 (.Y (nx17207), .A0 (nx17209), .A1 (nx17211), .A2 (nx17214), .A3 (
          nx17216)) ;
    aoi222 ix17210 (.Y (nx17209), .A0 (Mem_11__3), .A1 (nx17529), .B0 (Mem_15__3
           ), .B1 (nx17853), .C0 (Mem_8__3), .C1 (nx17525)) ;
    aoi221 ix17212 (.Y (nx17211), .A0 (Mem_19__3), .A1 (nx17809), .B0 (Mem_22__3
           ), .B1 (nx17805), .C0 (nx6030)) ;
    oai22 ix6031 (.Y (nx6030), .A0 (nx15428), .A1 (nx17087), .B0 (nx16271), .B1 (
          nx17641)) ;
    aoi222 ix17215 (.Y (nx17214), .A0 (Mem_31__3), .A1 (nx17519), .B0 (Mem_23__3
           ), .B1 (nx17851), .C0 (Mem_24__3), .C1 (nx17513)) ;
    aoi221 ix17217 (.Y (nx17216), .A0 (Mem_13__3), .A1 (nx17801), .B0 (Mem_9__3)
           , .B1 (nx17797), .C0 (nx6004)) ;
    oai22 ix6005 (.Y (nx6004), .A0 (nx15449), .A1 (nx17112), .B0 (nx16344), .B1 (
          nx17649)) ;
    and03 ix17220 (.Y (nx17219), .A0 (nx17221), .A1 (nx17223), .A2 (nx17225)) ;
    aoi222 ix17222 (.Y (nx17221), .A0 (Mem_29__3), .A1 (nx17509), .B0 (Mem_10__3
           ), .B1 (nx17505), .C0 (Mem_25__3), .C1 (nx17849)) ;
    aoi22 ix17224 (.Y (nx17223), .A0 (Mem_18__3), .A1 (nx17495), .B0 (Mem_26__3)
          , .B1 (nx17499)) ;
    aoi22 ix17226 (.Y (nx17225), .A0 (Mem_17__3), .A1 (nx17789), .B0 (Mem_27__3)
          , .B1 (nx17793)) ;
    aoi222 ix17228 (.Y (nx17227), .A0 (Mem_21__3), .A1 (nx17489), .B0 (Mem_16__3
           ), .B1 (nx17485), .C0 (Mem_5__3), .C1 (nx17847)) ;
    aoi221 ix17230 (.Y (nx17229), .A0 (Mem_30__3), .A1 (nx17779), .B0 (Mem_14__3
           ), .B1 (nx17481), .C0 (nx5956)) ;
    oai22 ix5957 (.Y (nx5956), .A0 (nx16251), .A1 (nx17149), .B0 (nx15444), .B1 (
          nx17653)) ;
    nand04 ix6165 (.Y (Dout[36]), .A0 (nx17233), .A1 (nx17245), .A2 (nx17253), .A3 (
           nx17255)) ;
    and04 ix17234 (.Y (nx17233), .A0 (nx17235), .A1 (nx17237), .A2 (nx17240), .A3 (
          nx17242)) ;
    aoi222 ix17236 (.Y (nx17235), .A0 (Mem_11__4), .A1 (nx17529), .B0 (Mem_15__4
           ), .B1 (nx17853), .C0 (Mem_8__4), .C1 (nx17525)) ;
    aoi221 ix17238 (.Y (nx17237), .A0 (Mem_19__4), .A1 (nx17809), .B0 (Mem_22__4
           ), .B1 (nx17805), .C0 (nx6140)) ;
    oai22 ix6141 (.Y (nx6140), .A0 (nx15461), .A1 (nx17087), .B0 (nx16373), .B1 (
          nx17641)) ;
    aoi222 ix17241 (.Y (nx17240), .A0 (Mem_31__4), .A1 (nx17519), .B0 (Mem_23__4
           ), .B1 (nx17851), .C0 (Mem_24__4), .C1 (nx17513)) ;
    aoi221 ix17243 (.Y (nx17242), .A0 (Mem_13__4), .A1 (nx17801), .B0 (Mem_9__4)
           , .B1 (nx17797), .C0 (nx6114)) ;
    oai22 ix6115 (.Y (nx6114), .A0 (nx15482), .A1 (nx17112), .B0 (nx16446), .B1 (
          nx17649)) ;
    and03 ix17246 (.Y (nx17245), .A0 (nx17247), .A1 (nx17249), .A2 (nx17251)) ;
    aoi222 ix17248 (.Y (nx17247), .A0 (Mem_29__4), .A1 (nx17509), .B0 (Mem_10__4
           ), .B1 (nx17505), .C0 (Mem_25__4), .C1 (nx17849)) ;
    aoi22 ix17250 (.Y (nx17249), .A0 (Mem_18__4), .A1 (nx17495), .B0 (Mem_26__4)
          , .B1 (nx17499)) ;
    aoi22 ix17252 (.Y (nx17251), .A0 (Mem_17__4), .A1 (nx17789), .B0 (Mem_27__4)
          , .B1 (nx17793)) ;
    aoi222 ix17254 (.Y (nx17253), .A0 (Mem_21__4), .A1 (nx17489), .B0 (Mem_16__4
           ), .B1 (nx17485), .C0 (Mem_5__4), .C1 (nx17847)) ;
    aoi221 ix17256 (.Y (nx17255), .A0 (Mem_30__4), .A1 (nx17779), .B0 (Mem_14__4
           ), .B1 (nx17481), .C0 (nx6066)) ;
    oai22 ix6067 (.Y (nx6066), .A0 (nx16353), .A1 (nx17149), .B0 (nx15477), .B1 (
          nx17653)) ;
    nand04 ix6275 (.Y (Dout[37]), .A0 (nx17259), .A1 (nx17271), .A2 (nx17279), .A3 (
           nx17281)) ;
    and04 ix17260 (.Y (nx17259), .A0 (nx17261), .A1 (nx17263), .A2 (nx17266), .A3 (
          nx17268)) ;
    aoi222 ix17262 (.Y (nx17261), .A0 (Mem_11__5), .A1 (nx17529), .B0 (Mem_15__5
           ), .B1 (nx17853), .C0 (Mem_8__5), .C1 (nx17525)) ;
    aoi221 ix17264 (.Y (nx17263), .A0 (Mem_19__5), .A1 (nx17809), .B0 (Mem_22__5
           ), .B1 (nx17805), .C0 (nx6250)) ;
    oai22 ix6251 (.Y (nx6250), .A0 (nx15494), .A1 (nx17087), .B0 (nx16475), .B1 (
          nx17641)) ;
    aoi222 ix17267 (.Y (nx17266), .A0 (Mem_31__5), .A1 (nx17519), .B0 (Mem_23__5
           ), .B1 (nx17851), .C0 (Mem_24__5), .C1 (nx17513)) ;
    aoi221 ix17269 (.Y (nx17268), .A0 (Mem_13__5), .A1 (nx17801), .B0 (Mem_9__5)
           , .B1 (nx17797), .C0 (nx6224)) ;
    oai22 ix6225 (.Y (nx6224), .A0 (nx15515), .A1 (nx17112), .B0 (nx16548), .B1 (
          nx17649)) ;
    and03 ix17272 (.Y (nx17271), .A0 (nx17273), .A1 (nx17275), .A2 (nx17277)) ;
    aoi222 ix17274 (.Y (nx17273), .A0 (Mem_29__5), .A1 (nx17509), .B0 (Mem_10__5
           ), .B1 (nx17505), .C0 (Mem_25__5), .C1 (nx17849)) ;
    aoi22 ix17276 (.Y (nx17275), .A0 (Mem_18__5), .A1 (nx17495), .B0 (Mem_26__5)
          , .B1 (nx17499)) ;
    aoi22 ix17278 (.Y (nx17277), .A0 (Mem_17__5), .A1 (nx17789), .B0 (Mem_27__5)
          , .B1 (nx17793)) ;
    aoi222 ix17280 (.Y (nx17279), .A0 (Mem_21__5), .A1 (nx17489), .B0 (Mem_16__5
           ), .B1 (nx17485), .C0 (Mem_5__5), .C1 (nx17847)) ;
    aoi221 ix17282 (.Y (nx17281), .A0 (Mem_30__5), .A1 (nx17779), .B0 (Mem_14__5
           ), .B1 (nx17481), .C0 (nx6176)) ;
    oai22 ix6177 (.Y (nx6176), .A0 (nx16455), .A1 (nx17149), .B0 (nx15510), .B1 (
          nx17653)) ;
    nand04 ix6385 (.Y (Dout[38]), .A0 (nx17285), .A1 (nx17297), .A2 (nx17305), .A3 (
           nx17307)) ;
    and04 ix17286 (.Y (nx17285), .A0 (nx17287), .A1 (nx17289), .A2 (nx17292), .A3 (
          nx17294)) ;
    aoi222 ix17288 (.Y (nx17287), .A0 (Mem_11__6), .A1 (nx17529), .B0 (Mem_15__6
           ), .B1 (nx5704), .C0 (Mem_8__6), .C1 (nx17525)) ;
    aoi221 ix17290 (.Y (nx17289), .A0 (Mem_19__6), .A1 (nx17809), .B0 (Mem_22__6
           ), .B1 (nx17805), .C0 (nx6360)) ;
    oai22 ix6361 (.Y (nx6360), .A0 (nx15527), .A1 (nx17087), .B0 (nx16577), .B1 (
          nx17641)) ;
    aoi222 ix17293 (.Y (nx17292), .A0 (Mem_31__6), .A1 (nx17519), .B0 (Mem_23__6
           ), .B1 (nx5668), .C0 (Mem_24__6), .C1 (nx17513)) ;
    aoi221 ix17295 (.Y (nx17294), .A0 (Mem_13__6), .A1 (nx17801), .B0 (Mem_9__6)
           , .B1 (nx17797), .C0 (nx6334)) ;
    oai22 ix6335 (.Y (nx6334), .A0 (nx15548), .A1 (nx17112), .B0 (nx16650), .B1 (
          nx17649)) ;
    and03 ix17298 (.Y (nx17297), .A0 (nx17299), .A1 (nx17301), .A2 (nx17303)) ;
    aoi222 ix17300 (.Y (nx17299), .A0 (Mem_29__6), .A1 (nx17509), .B0 (Mem_10__6
           ), .B1 (nx17505), .C0 (Mem_25__6), .C1 (nx5616)) ;
    aoi22 ix17302 (.Y (nx17301), .A0 (Mem_18__6), .A1 (nx17495), .B0 (Mem_26__6)
          , .B1 (nx17499)) ;
    aoi22 ix17304 (.Y (nx17303), .A0 (Mem_17__6), .A1 (nx17789), .B0 (Mem_27__6)
          , .B1 (nx17793)) ;
    aoi222 ix17306 (.Y (nx17305), .A0 (Mem_21__6), .A1 (nx17489), .B0 (Mem_16__6
           ), .B1 (nx17485), .C0 (Mem_5__6), .C1 (nx5566)) ;
    aoi221 ix17308 (.Y (nx17307), .A0 (Mem_30__6), .A1 (nx17779), .B0 (Mem_14__6
           ), .B1 (nx17481), .C0 (nx6286)) ;
    oai22 ix6287 (.Y (nx6286), .A0 (nx16557), .A1 (nx17149), .B0 (nx15543), .B1 (
          nx17653)) ;
    nand04 ix6495 (.Y (Dout[39]), .A0 (nx17311), .A1 (nx17323), .A2 (nx17331), .A3 (
           nx17333)) ;
    and04 ix17312 (.Y (nx17311), .A0 (nx17313), .A1 (nx17315), .A2 (nx17318), .A3 (
          nx17320)) ;
    aoi222 ix17314 (.Y (nx17313), .A0 (Mem_11__7), .A1 (nx17531), .B0 (Mem_15__7
           ), .B1 (nx5704), .C0 (Mem_8__7), .C1 (nx17527)) ;
    aoi221 ix17316 (.Y (nx17315), .A0 (Mem_19__7), .A1 (nx17811), .B0 (Mem_22__7
           ), .B1 (nx17807), .C0 (nx6470)) ;
    oai22 ix6471 (.Y (nx6470), .A0 (nx15560), .A1 (nx17087), .B0 (nx16679), .B1 (
          nx17643)) ;
    aoi222 ix17319 (.Y (nx17318), .A0 (Mem_31__7), .A1 (nx17521), .B0 (Mem_23__7
           ), .B1 (nx5668), .C0 (Mem_24__7), .C1 (nx17515)) ;
    aoi221 ix17321 (.Y (nx17320), .A0 (Mem_13__7), .A1 (nx17803), .B0 (Mem_9__7)
           , .B1 (nx17799), .C0 (nx6444)) ;
    oai22 ix6445 (.Y (nx6444), .A0 (nx15581), .A1 (nx17112), .B0 (nx16752), .B1 (
          nx17651)) ;
    and03 ix17324 (.Y (nx17323), .A0 (nx17325), .A1 (nx17327), .A2 (nx17329)) ;
    aoi222 ix17326 (.Y (nx17325), .A0 (Mem_29__7), .A1 (nx17511), .B0 (Mem_10__7
           ), .B1 (nx17507), .C0 (Mem_25__7), .C1 (nx5616)) ;
    aoi22 ix17328 (.Y (nx17327), .A0 (Mem_18__7), .A1 (nx17497), .B0 (Mem_26__7)
          , .B1 (nx17501)) ;
    aoi22 ix17330 (.Y (nx17329), .A0 (Mem_17__7), .A1 (nx17791), .B0 (Mem_27__7)
          , .B1 (nx17795)) ;
    aoi222 ix17332 (.Y (nx17331), .A0 (Mem_21__7), .A1 (nx17491), .B0 (Mem_16__7
           ), .B1 (nx17487), .C0 (Mem_5__7), .C1 (nx5566)) ;
    aoi221 ix17334 (.Y (nx17333), .A0 (Mem_30__7), .A1 (nx17781), .B0 (Mem_14__7
           ), .B1 (nx17483), .C0 (nx6396)) ;
    oai22 ix6397 (.Y (nx6396), .A0 (nx16659), .A1 (nx17149), .B0 (nx15576), .B1 (
          nx17655)) ;
    inv01 ix5641 (.Y (nx5640), .A (nx17075)) ;
    inv02 ix17068 (.Y (nx17067), .A (nx5510)) ;
    inv01 ix4483 (.Y (nx4482), .A (nx16760)) ;
    inv01 ix4445 (.Y (nx4444), .A (nx16764)) ;
    inv01 ix16785 (.Y (nx16784), .A (nx4436)) ;
    inv01 ix4429 (.Y (nx4428), .A (nx16778)) ;
    inv01 ix4421 (.Y (nx4420), .A (nx16770)) ;
    inv01 ix15888 (.Y (nx15887), .A (nx2196)) ;
    inv01 ix15818 (.Y (nx15817), .A (nx2180)) ;
    inv01 ix2171 (.Y (nx2170), .A (nx15819)) ;
    inv01 ix15757 (.Y (nx15756), .A (nx2066)) ;
    inv01 ix15913 (.Y (nx15912), .A (nx1950)) ;
    inv01 ix15705 (.Y (nx15704), .A (nx1932)) ;
    inv01 ix15792 (.Y (nx15791), .A (nx1770)) ;
    inv01 ix15980 (.Y (nx15979), .A (nx1762)) ;
    inv01 ix1745 (.Y (nx1744), .A (nx15944)) ;
    inv01 ix15998 (.Y (nx15997), .A (nx1692)) ;
    inv01 ix1633 (.Y (nx1632), .A (nx15715)) ;
    inv01 ix15954 (.Y (nx15953), .A (nx1594)) ;
    inv01 ix1585 (.Y (nx1584), .A (nx15956)) ;
    inv01 ix15772 (.Y (nx15771), .A (nx1552)) ;
    inv01 ix1547 (.Y (nx1546), .A (nx15746)) ;
    inv01 ix16019 (.Y (nx16018), .A (nx1502)) ;
    inv01 ix15597 (.Y (nx15596), .A (nx1152)) ;
    inv01 ix15876 (.Y (nx15875), .A (nx1138)) ;
    inv01 ix15734 (.Y (nx15733), .A (nx1130)) ;
    inv01 ix1123 (.Y (nx1122), .A (nx15873)) ;
    inv01 ix15193 (.Y (nx15192), .A (nx458)) ;
    inv01 ix447 (.Y (nx446), .A (nx15230)) ;
    inv01 ix437 (.Y (nx436), .A (nx15210)) ;
    inv01 ix15834 (.Y (nx15833), .A (nx430)) ;
    inv02 ix423 (.Y (nx422), .A (nx15203)) ;
    inv01 ix15259 (.Y (nx15258), .A (nx346)) ;
    inv01 ix327 (.Y (nx326), .A (nx15260)) ;
    inv01 ix15227 (.Y (nx15226), .A (nx204)) ;
    inv01 ix15992 (.Y (nx15991), .A (nx198)) ;
    inv01 ix189 (.Y (nx188), .A (nx15316)) ;
    inv01 ix185 (.Y (nx184), .A (nx15318)) ;
    inv01 ix15307 (.Y (nx15306), .A (nx166)) ;
    inv01 ix15940 (.Y (nx15939), .A (nx158)) ;
    inv02 ix125 (.Y (nx124), .A (nx15286)) ;
    inv01 ix121 (.Y (nx120), .A (nx15242)) ;
    inv01 ix15878 (.Y (nx15877), .A (nx108)) ;
    inv01 ix81 (.Y (nx80), .A (nx15200)) ;
    inv01 ix75 (.Y (nx74), .A (nx15180)) ;
    inv01 ix65 (.Y (nx64), .A (nx15343)) ;
    inv02 ix15187 (.Y (nx15186), .A (nx44)) ;
    inv01 ix33 (.Y (nx32), .A (nx15348)) ;
    inv01 ix15814 (.Y (nx15813), .A (nx22)) ;
    inv01 ix15282 (.Y (nx15281), .A (nx14)) ;
    inv01 ix3 (.Y (nx2), .A (nx15301)) ;
    inv02 ix17340 (.Y (nx17341), .A (nx15186)) ;
    inv02 ix17342 (.Y (nx17343), .A (nx15308)) ;
    buf02 ix17346 (.Y (nx17347), .A (nx212)) ;
    buf02 ix17348 (.Y (nx17349), .A (nx212)) ;
    buf02 ix17350 (.Y (nx17351), .A (nx258)) ;
    buf02 ix17352 (.Y (nx17353), .A (nx258)) ;
    buf02 ix17354 (.Y (nx17355), .A (nx366)) ;
    buf02 ix17356 (.Y (nx17357), .A (nx366)) ;
    buf02 ix17358 (.Y (nx17359), .A (nx404)) ;
    buf02 ix17360 (.Y (nx17361), .A (nx404)) ;
    buf02 ix17362 (.Y (nx17363), .A (nx464)) ;
    buf02 ix17364 (.Y (nx17365), .A (nx464)) ;
    buf02 ix17366 (.Y (nx17367), .A (nx504)) ;
    buf02 ix17368 (.Y (nx17369), .A (nx504)) ;
    buf02 ix17370 (.Y (nx17371), .A (nx1162)) ;
    buf02 ix17372 (.Y (nx17373), .A (nx1162)) ;
    buf02 ix17374 (.Y (nx17375), .A (nx1522)) ;
    buf02 ix17376 (.Y (nx17377), .A (nx1522)) ;
    inv02 ix17378 (.Y (nx17379), .A (nx17829)) ;
    buf02 ix17380 (.Y (nx17381), .A (nx1616)) ;
    buf02 ix17382 (.Y (nx17383), .A (nx1616)) ;
    buf02 ix17384 (.Y (nx17385), .A (nx1664)) ;
    buf02 ix17386 (.Y (nx17387), .A (nx1664)) ;
    buf02 ix17388 (.Y (nx17389), .A (nx1730)) ;
    buf02 ix17390 (.Y (nx17391), .A (nx1730)) ;
    buf02 ix17392 (.Y (nx17393), .A (nx1824)) ;
    buf02 ix17394 (.Y (nx17395), .A (nx1824)) ;
    buf02 ix17396 (.Y (nx17397), .A (nx1904)) ;
    buf02 ix17398 (.Y (nx17399), .A (nx1904)) ;
    buf02 ix17404 (.Y (nx17405), .A (nx2010)) ;
    buf02 ix17406 (.Y (nx17407), .A (nx2010)) ;
    buf02 ix17408 (.Y (nx17409), .A (nx2046)) ;
    buf02 ix17410 (.Y (nx17411), .A (nx2046)) ;
    buf02 ix17412 (.Y (nx17413), .A (nx2096)) ;
    buf02 ix17414 (.Y (nx17415), .A (nx2096)) ;
    buf02 ix17416 (.Y (nx17417), .A (nx2150)) ;
    buf02 ix17418 (.Y (nx17419), .A (nx2150)) ;
    buf02 ix17420 (.Y (nx17421), .A (nx2204)) ;
    buf02 ix17422 (.Y (nx17423), .A (nx2204)) ;
    buf02 ix17424 (.Y (nx17425), .A (nx2288)) ;
    buf02 ix17426 (.Y (nx17427), .A (nx2288)) ;
    buf02 ix17428 (.Y (nx17429), .A (nx2326)) ;
    buf02 ix17430 (.Y (nx17431), .A (nx2326)) ;
    buf02 ix17432 (.Y (nx17433), .A (nx2448)) ;
    buf02 ix17434 (.Y (nx17435), .A (nx2448)) ;
    buf02 ix17436 (.Y (nx17437), .A (nx2486)) ;
    buf02 ix17438 (.Y (nx17439), .A (nx2486)) ;
    buf02 ix17440 (.Y (nx17441), .A (nx2538)) ;
    buf02 ix17442 (.Y (nx17443), .A (nx2538)) ;
    buf02 ix17446 (.Y (nx17447), .A (nx2604)) ;
    buf02 ix17448 (.Y (nx17449), .A (nx2604)) ;
    buf02 ix17454 (.Y (nx17455), .A (nx4576)) ;
    buf02 ix17456 (.Y (nx17457), .A (nx4576)) ;
    buf02 ix17458 (.Y (nx17459), .A (nx4586)) ;
    buf02 ix17460 (.Y (nx17461), .A (nx4586)) ;
    buf02 ix17464 (.Y (nx17465), .A (nx4632)) ;
    buf02 ix17466 (.Y (nx17467), .A (nx4632)) ;
    buf02 ix17472 (.Y (nx17473), .A (nx4672)) ;
    buf02 ix17474 (.Y (nx17475), .A (nx4672)) ;
    buf02 ix17476 (.Y (nx17477), .A (nx4676)) ;
    buf02 ix17478 (.Y (nx17479), .A (nx4676)) ;
    buf02 ix17480 (.Y (nx17481), .A (nx5512)) ;
    buf02 ix17482 (.Y (nx17483), .A (nx5512)) ;
    buf02 ix17484 (.Y (nx17485), .A (nx5552)) ;
    buf02 ix17486 (.Y (nx17487), .A (nx5552)) ;
    buf02 ix17488 (.Y (nx17489), .A (nx5562)) ;
    buf02 ix17490 (.Y (nx17491), .A (nx5562)) ;
    buf02 ix17494 (.Y (nx17495), .A (nx5604)) ;
    buf02 ix17496 (.Y (nx17497), .A (nx5604)) ;
    buf02 ix17498 (.Y (nx17499), .A (nx5608)) ;
    buf02 ix17500 (.Y (nx17501), .A (nx5608)) ;
    buf02 ix17504 (.Y (nx17505), .A (nx5620)) ;
    buf02 ix17506 (.Y (nx17507), .A (nx5620)) ;
    buf02 ix17508 (.Y (nx17509), .A (nx5624)) ;
    buf02 ix17510 (.Y (nx17511), .A (nx5624)) ;
    buf02 ix17512 (.Y (nx17513), .A (nx5664)) ;
    buf02 ix17514 (.Y (nx17515), .A (nx5664)) ;
    buf02 ix17518 (.Y (nx17519), .A (nx5672)) ;
    buf02 ix17520 (.Y (nx17521), .A (nx5672)) ;
    buf02 ix17524 (.Y (nx17525), .A (nx5708)) ;
    buf02 ix17526 (.Y (nx17527), .A (nx5708)) ;
    buf02 ix17528 (.Y (nx17529), .A (nx5712)) ;
    buf02 ix17530 (.Y (nx17531), .A (nx5712)) ;
    inv02 ix17532 (.Y (nx17533), .A (Address[2])) ;
    inv02 ix17534 (.Y (nx17535), .A (Address[2])) ;
    inv02 ix17536 (.Y (nx17537), .A (Address[4])) ;
    inv02 ix17538 (.Y (nx17539), .A (Address[4])) ;
    inv02 ix17542 (.Y (nx17543), .A (nx17675)) ;
    inv02 ix17544 (.Y (nx17545), .A (Address[1])) ;
    inv02 ix17546 (.Y (nx17547), .A (Address[1])) ;
    inv02 ix17548 (.Y (nx17549), .A (Address[14])) ;
    inv02 ix17550 (.Y (nx17551), .A (Address[14])) ;
    inv02 ix17552 (.Y (nx17553), .A (nx17673)) ;
    buf02 ix17554 (.Y (nx17555), .A (nx15296)) ;
    buf02 ix17556 (.Y (nx17557), .A (nx15296)) ;
    buf02 ix17560 (.Y (nx17561), .A (nx15341)) ;
    buf02 ix17562 (.Y (nx17563), .A (nx15341)) ;
    buf02 ix17564 (.Y (nx17565), .A (nx15702)) ;
    buf02 ix17566 (.Y (nx17567), .A (nx15702)) ;
    buf02 ix17568 (.Y (nx17569), .A (nx15731)) ;
    buf02 ix17570 (.Y (nx17571), .A (nx15731)) ;
    inv02 ix17572 (.Y (nx17573), .A (nx1546)) ;
    buf02 ix17574 (.Y (nx17575), .A (nx15811)) ;
    buf02 ix17576 (.Y (nx17577), .A (nx15811)) ;
    buf02 ix17578 (.Y (nx17579), .A (nx15828)) ;
    buf02 ix17580 (.Y (nx17581), .A (nx15828)) ;
    buf02 ix17582 (.Y (nx17583), .A (nx15836)) ;
    buf02 ix17584 (.Y (nx17585), .A (nx15836)) ;
    buf02 ix17586 (.Y (nx17587), .A (nx15869)) ;
    buf02 ix17588 (.Y (nx17589), .A (nx15869)) ;
    buf02 ix17590 (.Y (nx17591), .A (nx15936)) ;
    buf02 ix17592 (.Y (nx17593), .A (nx15936)) ;
    buf02 ix17594 (.Y (nx17595), .A (nx15950)) ;
    buf02 ix17596 (.Y (nx17597), .A (nx15950)) ;
    buf02 ix17598 (.Y (nx17599), .A (nx15971)) ;
    buf02 ix17600 (.Y (nx17601), .A (nx15971)) ;
    buf02 ix17602 (.Y (nx17603), .A (nx15989)) ;
    buf02 ix17604 (.Y (nx17605), .A (nx15989)) ;
    buf02 ix17606 (.Y (nx17607), .A (nx16003)) ;
    buf02 ix17608 (.Y (nx17609), .A (nx16003)) ;
    nand02 ix17610 (.Y (nx17611), .A0 (nx17823), .A1 (nx1572)) ;
    nand02 ix17612 (.Y (nx17613), .A0 (nx17829), .A1 (nx1558)) ;
    buf02 ix17614 (.Y (nx17615), .A (nx16767)) ;
    inv02 ix17616 (.Y (nx17617), .A (nx4428)) ;
    buf02 ix17618 (.Y (nx17619), .A (nx16797)) ;
    buf02 ix17620 (.Y (nx17621), .A (nx16797)) ;
    nand02 ix17622 (.Y (nx17623), .A0 (Address[5]), .A1 (Address[6])) ;
    nand02 ix17624 (.Y (nx17625), .A0 (nx17741), .A1 (nx4514)) ;
    nand02 ix17626 (.Y (nx17627), .A0 (nx17743), .A1 (nx4470)) ;
    buf02 ix17628 (.Y (nx17629), .A (nx16858)) ;
    buf02 ix17630 (.Y (nx17631), .A (nx16858)) ;
    buf02 ix17632 (.Y (nx17633), .A (nx16863)) ;
    buf02 ix17634 (.Y (nx17635), .A (nx16863)) ;
    inv02 ix17636 (.Y (nx17637), .A (nx17787)) ;
    buf02 ix17640 (.Y (nx17641), .A (nx17093)) ;
    buf02 ix17642 (.Y (nx17643), .A (nx17093)) ;
    inv02 ix17644 (.Y (nx17645), .A (nx5496)) ;
    buf02 ix17648 (.Y (nx17649), .A (nx17115)) ;
    buf02 ix17650 (.Y (nx17651), .A (nx17115)) ;
    buf02 ix17652 (.Y (nx17653), .A (nx17152)) ;
    buf02 ix17654 (.Y (nx17655), .A (nx17152)) ;
    nor02ii ix431 (.Y (nx430), .A0 (Address[6]), .A1 (nx44)) ;
    nor02ii ix163 (.Y (nx15308), .A0 (Address[11]), .A1 (Address[10])) ;
    nor02ii ix15243 (.Y (nx15242), .A0 (Address[5]), .A1 (Address[4])) ;
    nor02ii ix15261 (.Y (nx15260), .A0 (Address[9]), .A1 (Address[8])) ;
    nor02ii ix417 (.Y (nx416), .A0 (Address[17]), .A1 (nx15318)) ;
    and02 ix377 (.Y (nx376), .A0 (Address[17]), .A1 (nx15318)) ;
    nor02ii ix15302 (.Y (nx15301), .A0 (Address[1]), .A1 (Address[2])) ;
    nor02ii ix29 (.Y (nx28), .A0 (Address[12]), .A1 (WR)) ;
    nor02ii ix15319 (.Y (nx15318), .A0 (Address[16]), .A1 (Address[15])) ;
    nor02ii ix15325 (.Y (nx15324), .A0 (Address[0]), .A1 (Address[1])) ;
    nor02ii ix309 (.Y (nx308), .A0 (nx108), .A1 (Address[17])) ;
    nor02ii ix229 (.Y (nx228), .A0 (nx224), .A1 (Address[17])) ;
    nor02ii ix15344 (.Y (nx15343), .A0 (Address[13]), .A1 (Address[14])) ;
    nor02ii ix15601 (.Y (nx15600), .A0 (Address[10]), .A1 (Address[11])) ;
    nor02ii ix2539 (.Y (nx2538), .A0 (nx15720), .A1 (nx17825)) ;
    nor02ii ix2577 (.Y (nx2576), .A0 (nx15744), .A1 (nx17827)) ;
    nor02ii ix1481 (.Y (nx1480), .A0 (nx354), .A1 (Address[4])) ;
    nor02ii ix2497 (.Y (nx2496), .A0 (nx15769), .A1 (nx17827)) ;
    nor02ii ix2259 (.Y (nx2258), .A0 (nx15881), .A1 (nx17823)) ;
    nor02ii ix1693 (.Y (nx1692), .A0 (nx1540), .A1 (nx15746)) ;
    nor02ii ix2123 (.Y (nx2122), .A0 (nx15881), .A1 (nx17827)) ;
    nor02ii ix2115 (.Y (nx2114), .A0 (nx15769), .A1 (nx15350)) ;
    nor02ii ix1973 (.Y (nx1972), .A0 (nx15720), .A1 (nx15350)) ;
    nor02ii ix1873 (.Y (nx1872), .A0 (nx15744), .A1 (nx15350)) ;
    nor02ii ix4431 (.Y (nx4430), .A0 (nx17615), .A1 (Address[8])) ;
    nor02ii ix4669 (.Y (nx4668), .A0 (nx16776), .A1 (nx17743)) ;
    nor02ii ix4491 (.Y (nx4490), .A0 (Address[6]), .A1 (Address[5])) ;
    nor02ii ix4647 (.Y (nx4646), .A0 (nx16762), .A1 (nx17743)) ;
    nor02ii ix4651 (.Y (nx4650), .A0 (nx16760), .A1 (nx4584)) ;
    nor02ii ix4637 (.Y (nx4636), .A0 (nx17623), .A1 (nx4470)) ;
    nor02ii ix4629 (.Y (nx4628), .A0 (nx17623), .A1 (nx4584)) ;
    nor02ii ix4607 (.Y (nx4606), .A0 (nx16776), .A1 (nx17741)) ;
    nor02ii ix4577 (.Y (nx4576), .A0 (nx16762), .A1 (nx4454)) ;
    nor02ii ix4567 (.Y (nx4566), .A0 (nx17623), .A1 (nx4498)) ;
    nor02ii ix4555 (.Y (nx4554), .A0 (nx16836), .A1 (nx17745)) ;
    nor02ii ix4549 (.Y (nx4548), .A0 (nx16805), .A1 (nx4514)) ;
    nor02ii ix4545 (.Y (nx4544), .A0 (nx16836), .A1 (nx4454)) ;
    nor02ii ix4535 (.Y (nx4534), .A0 (nx16760), .A1 (nx4498)) ;
    nor02ii ix5523 (.Y (nx5522), .A0 (nx5494), .A1 (nx17069)) ;
    nor02ii ix17100 (.Y (nx5496), .A0 (nx17069), .A1 (nx5494)) ;
    inv01 ix17668 (.Y (nx17669), .A (Address[0])) ;
    nor02ii ix5567 (.Y (nx5566), .A0 (nx17106), .A1 (nx5522)) ;
    nor02ii ix17402 (.Y (nx17403), .A0 (nx15720), .A1 (nx15350)) ;
    nor02ii ix17444 (.Y (nx17445), .A0 (nx15744), .A1 (nx17827)) ;
    nor02ii ix17452 (.Y (nx17453), .A0 (nx16805), .A1 (nx4498)) ;
    nor02ii ix17462 (.Y (nx17463), .A0 (nx16805), .A1 (nx4584)) ;
    nor02ii ix17468 (.Y (nx17469), .A0 (nx16805), .A1 (nx4470)) ;
    nor02ii ix17470 (.Y (nx17471), .A0 (nx16776), .A1 (nx17745)) ;
    nor02ii ix17492 (.Y (nx17493), .A0 (nx17106), .A1 (nx5522)) ;
    inv02 ix17670 (.Y (nx17671), .A (nx17559)) ;
    inv02 ix17672 (.Y (nx17673), .A (nx15286)) ;
    inv02 ix17674 (.Y (nx17675), .A (nx17541)) ;
    buf02 ix17678 (.Y (nx17679), .A (nx228)) ;
    buf02 ix17680 (.Y (nx17681), .A (nx228)) ;
    buf02 ix17682 (.Y (nx17683), .A (nx308)) ;
    buf02 ix17684 (.Y (nx17685), .A (nx308)) ;
    buf02 ix17686 (.Y (nx17687), .A (nx416)) ;
    buf02 ix17688 (.Y (nx17689), .A (nx416)) ;
    inv01 ix17690 (.Y (nx17691), .A (nx15833)) ;
    buf02 ix17692 (.Y (nx17693), .A (nx1480)) ;
    buf02 ix17694 (.Y (nx17695), .A (nx1488)) ;
    buf02 ix17696 (.Y (nx17697), .A (nx1794)) ;
    buf02 ix17698 (.Y (nx17699), .A (nx1794)) ;
    buf02 ix17700 (.Y (nx17701), .A (nx1834)) ;
    buf02 ix17702 (.Y (nx17703), .A (nx1834)) ;
    buf02 ix17704 (.Y (nx17705), .A (nx1872)) ;
    buf02 ix17706 (.Y (nx17707), .A (nx1872)) ;
    buf02 ix17708 (.Y (nx17709), .A (nx2056)) ;
    buf02 ix17710 (.Y (nx17711), .A (nx2056)) ;
    buf02 ix17712 (.Y (nx17713), .A (nx2114)) ;
    buf02 ix17714 (.Y (nx17715), .A (nx2114)) ;
    buf02 ix17716 (.Y (nx17717), .A (nx2122)) ;
    buf02 ix17718 (.Y (nx17719), .A (nx2122)) ;
    buf02 ix17720 (.Y (nx17721), .A (nx2160)) ;
    buf02 ix17722 (.Y (nx17723), .A (nx2160)) ;
    buf02 ix17724 (.Y (nx17725), .A (nx2258)) ;
    buf02 ix17726 (.Y (nx17727), .A (nx2258)) ;
    buf02 ix17728 (.Y (nx17729), .A (nx2298)) ;
    buf02 ix17730 (.Y (nx17731), .A (nx2298)) ;
    buf02 ix17732 (.Y (nx17733), .A (nx2458)) ;
    buf02 ix17734 (.Y (nx17735), .A (nx2458)) ;
    buf02 ix17736 (.Y (nx17737), .A (nx2496)) ;
    buf02 ix17738 (.Y (nx17739), .A (nx2496)) ;
    nor02_2x ix17740 (.Y (nx17741), .A0 (Address[5]), .A1 (Address[6])) ;
    buf02 ix17742 (.Y (nx17743), .A (nx4490)) ;
    buf02 ix17744 (.Y (nx17745), .A (nx4490)) ;
    buf02 ix17746 (.Y (nx17747), .A (nx4534)) ;
    buf02 ix17748 (.Y (nx17749), .A (nx4534)) ;
    buf02 ix17750 (.Y (nx17751), .A (nx4544)) ;
    buf02 ix17752 (.Y (nx17753), .A (nx4544)) ;
    buf02 ix17754 (.Y (nx17755), .A (nx4548)) ;
    buf02 ix17756 (.Y (nx17757), .A (nx4548)) ;
    buf02 ix17758 (.Y (nx17759), .A (nx4554)) ;
    buf02 ix17760 (.Y (nx17761), .A (nx4554)) ;
    buf02 ix17762 (.Y (nx17763), .A (nx4606)) ;
    buf02 ix17764 (.Y (nx17765), .A (nx4606)) ;
    buf02 ix17766 (.Y (nx17767), .A (nx4646)) ;
    buf02 ix17768 (.Y (nx17769), .A (nx4646)) ;
    buf02 ix17770 (.Y (nx17771), .A (nx4650)) ;
    buf02 ix17772 (.Y (nx17773), .A (nx4650)) ;
    inv01 ix17774 (.Y (nx17775), .A (nx18135)) ;
    buf02 ix17778 (.Y (nx17779), .A (nx5504)) ;
    buf02 ix17780 (.Y (nx17781), .A (nx5504)) ;
    inv01 ix17782 (.Y (nx17783), .A (nx18123)) ;
    inv01 ix17786 (.Y (nx17787), .A (nx17081)) ;
    buf02 ix17788 (.Y (nx17789), .A (nx5582)) ;
    buf02 ix17790 (.Y (nx17791), .A (nx5582)) ;
    buf02 ix17792 (.Y (nx17793), .A (nx5592)) ;
    buf02 ix17794 (.Y (nx17795), .A (nx5592)) ;
    buf02 ix17796 (.Y (nx17797), .A (nx5652)) ;
    buf02 ix17798 (.Y (nx17799), .A (nx5652)) ;
    buf02 ix17800 (.Y (nx17801), .A (nx5656)) ;
    buf02 ix17802 (.Y (nx17803), .A (nx5656)) ;
    buf02 ix17804 (.Y (nx17805), .A (nx5692)) ;
    buf02 ix17806 (.Y (nx17807), .A (nx5692)) ;
    buf02 ix17808 (.Y (nx17809), .A (nx5696)) ;
    buf02 ix17810 (.Y (nx17811), .A (nx5696)) ;
    inv01 ix17812 (.Y (nx17813), .A (nx120)) ;
    inv02 ix17814 (.Y (nx17815), .A (nx326)) ;
    inv01 ix17816 (.Y (nx17817), .A (nx18129)) ;
    buf02 ix17820 (.Y (nx17821), .A (nx15324)) ;
    nor02_2x ix17822 (.Y (nx17823), .A0 (Address[11]), .A1 (Address[10])) ;
    buf02 ix17824 (.Y (nx17825), .A (nx15600)) ;
    buf02 ix17826 (.Y (nx17827), .A (nx15600)) ;
    inv01 ix17828 (.Y (nx17829), .A (nx1534)) ;
    buf02 ix17830 (.Y (nx17831), .A (nx17401)) ;
    buf02 ix17832 (.Y (nx17833), .A (nx17403)) ;
    buf02 ix17834 (.Y (nx17835), .A (nx17445)) ;
    buf02 ix17836 (.Y (nx17837), .A (nx17451)) ;
    buf02 ix17838 (.Y (nx17839), .A (nx17453)) ;
    buf02 ix17840 (.Y (nx17841), .A (nx17463)) ;
    buf02 ix17842 (.Y (nx17843), .A (nx17469)) ;
    buf02 ix17844 (.Y (nx17845), .A (nx17471)) ;
    buf02 ix17846 (.Y (nx17847), .A (nx17493)) ;
    buf02 ix17848 (.Y (nx17849), .A (nx17503)) ;
    buf02 ix17850 (.Y (nx17851), .A (nx17517)) ;
    buf02 ix17852 (.Y (nx17853), .A (nx17523)) ;
    mux21 ix12685 (.Y (nx12684), .A0 (nx18137), .A1 (nx15244), .S0 (nx18051)) ;
    inv01 ix18048 (.Y (nx18049), .A (Din[0])) ;
    inv02 ix18050 (.Y (nx18051), .A (nx17367)) ;
    oai222 ix15229 (.Y (nx17665), .A0 (nx446), .A1 (nx15316), .B0 (nx436), .B1 (
           nx15306), .C0 (nx120), .C1 (nx15833)) ;
    mux21 ix12655 (.Y (nx12654), .A0 (nx18137), .A1 (nx15272), .S0 (nx18053)) ;
    inv02 ix18052 (.Y (nx18053), .A (nx17355)) ;
    mux21 ix12635 (.Y (nx12634), .A0 (nx18137), .A1 (nx15291), .S0 (nx18055)) ;
    inv02 ix18054 (.Y (nx18055), .A (nx17351)) ;
    mux21 ix12645 (.Y (nx12644), .A0 (nx18137), .A1 (nx15326), .S0 (nx17555)) ;
    mux21 ix12625 (.Y (nx12624), .A0 (nx18137), .A1 (nx15337), .S0 (nx18057)) ;
    inv02 ix18056 (.Y (nx18057), .A (nx17347)) ;
    mux21 ix12765 (.Y (nx12764), .A0 (nx18141), .A1 (nx15362), .S0 (nx18051)) ;
    inv01 ix18058 (.Y (nx18059), .A (Din[1])) ;
    mux21 ix12735 (.Y (nx12734), .A0 (nx18141), .A1 (nx15370), .S0 (nx18053)) ;
    mux21 ix12715 (.Y (nx12714), .A0 (nx18141), .A1 (nx15375), .S0 (nx18055)) ;
    mux21 ix12725 (.Y (nx12724), .A0 (nx18141), .A1 (nx15378), .S0 (nx17555)) ;
    mux21 ix12705 (.Y (nx12704), .A0 (nx18141), .A1 (nx15383), .S0 (nx18057)) ;
    mux21 ix12845 (.Y (nx12844), .A0 (nx18145), .A1 (nx15395), .S0 (nx18051)) ;
    inv01 ix18060 (.Y (nx18061), .A (Din[2])) ;
    mux21 ix12815 (.Y (nx12814), .A0 (nx18145), .A1 (nx15403), .S0 (nx18053)) ;
    mux21 ix12795 (.Y (nx12794), .A0 (nx18145), .A1 (nx15408), .S0 (nx18055)) ;
    mux21 ix12805 (.Y (nx12804), .A0 (nx18145), .A1 (nx15411), .S0 (nx17555)) ;
    mux21 ix12785 (.Y (nx12784), .A0 (nx18145), .A1 (nx15416), .S0 (nx18057)) ;
    mux21 ix12925 (.Y (nx12924), .A0 (nx18149), .A1 (nx15428), .S0 (nx18051)) ;
    inv01 ix18062 (.Y (nx18063), .A (Din[3])) ;
    mux21 ix12895 (.Y (nx12894), .A0 (nx18149), .A1 (nx15436), .S0 (nx18053)) ;
    mux21 ix12875 (.Y (nx12874), .A0 (nx18149), .A1 (nx15441), .S0 (nx18055)) ;
    mux21 ix12885 (.Y (nx12884), .A0 (nx18149), .A1 (nx15444), .S0 (nx17555)) ;
    mux21 ix12865 (.Y (nx12864), .A0 (nx18149), .A1 (nx15449), .S0 (nx18057)) ;
    mux21 ix13005 (.Y (nx13004), .A0 (nx18153), .A1 (nx15461), .S0 (nx18051)) ;
    inv01 ix18064 (.Y (nx18065), .A (Din[4])) ;
    mux21 ix12975 (.Y (nx12974), .A0 (nx18153), .A1 (nx15469), .S0 (nx18053)) ;
    mux21 ix12955 (.Y (nx12954), .A0 (nx18153), .A1 (nx15474), .S0 (nx18055)) ;
    mux21 ix12965 (.Y (nx12964), .A0 (nx18153), .A1 (nx15477), .S0 (nx17555)) ;
    mux21 ix12945 (.Y (nx12944), .A0 (nx18153), .A1 (nx15482), .S0 (nx18057)) ;
    mux21 ix13085 (.Y (nx13084), .A0 (nx18157), .A1 (nx15494), .S0 (nx18051)) ;
    inv01 ix18066 (.Y (nx18067), .A (Din[5])) ;
    mux21 ix13055 (.Y (nx13054), .A0 (nx18157), .A1 (nx15502), .S0 (nx18053)) ;
    mux21 ix13035 (.Y (nx13034), .A0 (nx18157), .A1 (nx15507), .S0 (nx18055)) ;
    mux21 ix13045 (.Y (nx13044), .A0 (nx18157), .A1 (nx15510), .S0 (nx17555)) ;
    mux21 ix13025 (.Y (nx13024), .A0 (nx18157), .A1 (nx15515), .S0 (nx18057)) ;
    mux21 ix13165 (.Y (nx13164), .A0 (nx18161), .A1 (nx15527), .S0 (nx18051)) ;
    inv01 ix18068 (.Y (nx18069), .A (Din[6])) ;
    mux21 ix13135 (.Y (nx13134), .A0 (nx18161), .A1 (nx15535), .S0 (nx18053)) ;
    mux21 ix13115 (.Y (nx13114), .A0 (nx18161), .A1 (nx15540), .S0 (nx18055)) ;
    mux21 ix13125 (.Y (nx13124), .A0 (nx18161), .A1 (nx15543), .S0 (nx17555)) ;
    mux21 ix13105 (.Y (nx13104), .A0 (nx18161), .A1 (nx15548), .S0 (nx18057)) ;
    mux21 ix13245 (.Y (nx13244), .A0 (nx18165), .A1 (nx15560), .S0 (nx18073)) ;
    inv01 ix18070 (.Y (nx18071), .A (Din[7])) ;
    inv01 ix18072 (.Y (nx18073), .A (nx17369)) ;
    mux21 ix13215 (.Y (nx13214), .A0 (nx18165), .A1 (nx15568), .S0 (nx18075)) ;
    inv01 ix18074 (.Y (nx18075), .A (nx17357)) ;
    mux21 ix13195 (.Y (nx13194), .A0 (nx18165), .A1 (nx15573), .S0 (nx18077)) ;
    inv01 ix18076 (.Y (nx18077), .A (nx17353)) ;
    mux21 ix13205 (.Y (nx13204), .A0 (nx18165), .A1 (nx15576), .S0 (nx17557)) ;
    mux21 ix13185 (.Y (nx13184), .A0 (nx18165), .A1 (nx15581), .S0 (nx18079)) ;
    inv01 ix18078 (.Y (nx18079), .A (nx17349)) ;
    mux21 ix13535 (.Y (nx13534), .A0 (nx18139), .A1 (nx15717), .S0 (nx17565)) ;
    mux21 ix13555 (.Y (nx13554), .A0 (nx18139), .A1 (nx15767), .S0 (nx18081)) ;
    inv02 ix18080 (.Y (nx18081), .A (nx17447)) ;
    mux21 ix13525 (.Y (nx13524), .A0 (nx18139), .A1 (nx15786), .S0 (nx18083)) ;
    inv02 ix18082 (.Y (nx18083), .A (nx17437)) ;
    mux21 ix13505 (.Y (nx13504), .A0 (nx18139), .A1 (nx15807), .S0 (nx17575)) ;
    mux21 ix13495 (.Y (nx13494), .A0 (nx18139), .A1 (nx15824), .S0 (nx17579)) ;
    mux21 ix13475 (.Y (nx13474), .A0 (nx18049), .A1 (nx15848), .S0 (nx18085)) ;
    inv02 ix18084 (.Y (nx18085), .A (nx17425)) ;
    mux21 ix13425 (.Y (nx13424), .A0 (nx18049), .A1 (nx15916), .S0 (nx18087)) ;
    inv02 ix18086 (.Y (nx18087), .A (nx17409)) ;
    mux21 ix13415 (.Y (nx13414), .A0 (nx18049), .A1 (nx15946), .S0 (nx17591)) ;
    mux21 ix13335 (.Y (nx13334), .A0 (nx18049), .A1 (nx16013), .S0 (nx18089)) ;
    inv02 ix18088 (.Y (nx18089), .A (nx17375)) ;
    mux21 ix13355 (.Y (nx13354), .A0 (nx18049), .A1 (nx16033), .S0 (nx18091)) ;
    inv02 ix18090 (.Y (nx18091), .A (nx17385)) ;
    mux21 ix13765 (.Y (nx13764), .A0 (nx18143), .A1 (nx16047), .S0 (nx17565)) ;
    mux21 ix13785 (.Y (nx13784), .A0 (nx18143), .A1 (nx16053), .S0 (nx18081)) ;
    mux21 ix13755 (.Y (nx13754), .A0 (nx18143), .A1 (nx16058), .S0 (nx18083)) ;
    mux21 ix13735 (.Y (nx13734), .A0 (nx18143), .A1 (nx16063), .S0 (nx17575)) ;
    mux21 ix13725 (.Y (nx13724), .A0 (nx18143), .A1 (nx16067), .S0 (nx17579)) ;
    mux21 ix13705 (.Y (nx13704), .A0 (nx18059), .A1 (nx16077), .S0 (nx18085)) ;
    mux21 ix13655 (.Y (nx13654), .A0 (nx18059), .A1 (nx16098), .S0 (nx18087)) ;
    mux21 ix13645 (.Y (nx13644), .A0 (nx18059), .A1 (nx16109), .S0 (nx17591)) ;
    mux21 ix13565 (.Y (nx13564), .A0 (nx18059), .A1 (nx16132), .S0 (nx18089)) ;
    mux21 ix13585 (.Y (nx13584), .A0 (nx18059), .A1 (nx16140), .S0 (nx18091)) ;
    mux21 ix13995 (.Y (nx13994), .A0 (nx18147), .A1 (nx16149), .S0 (nx17565)) ;
    mux21 ix14015 (.Y (nx14014), .A0 (nx18147), .A1 (nx16155), .S0 (nx18081)) ;
    mux21 ix13985 (.Y (nx13984), .A0 (nx18147), .A1 (nx16160), .S0 (nx18083)) ;
    mux21 ix13965 (.Y (nx13964), .A0 (nx18147), .A1 (nx16165), .S0 (nx17575)) ;
    mux21 ix13955 (.Y (nx13954), .A0 (nx18147), .A1 (nx16169), .S0 (nx17579)) ;
    mux21 ix13935 (.Y (nx13934), .A0 (nx18061), .A1 (nx16179), .S0 (nx18085)) ;
    mux21 ix13885 (.Y (nx13884), .A0 (nx18061), .A1 (nx16200), .S0 (nx18087)) ;
    mux21 ix13875 (.Y (nx13874), .A0 (nx18061), .A1 (nx16211), .S0 (nx17591)) ;
    mux21 ix13795 (.Y (nx13794), .A0 (nx18061), .A1 (nx16234), .S0 (nx18089)) ;
    mux21 ix13815 (.Y (nx13814), .A0 (nx18061), .A1 (nx16242), .S0 (nx18091)) ;
    mux21 ix14225 (.Y (nx14224), .A0 (nx18151), .A1 (nx16251), .S0 (nx17565)) ;
    mux21 ix14245 (.Y (nx14244), .A0 (nx18151), .A1 (nx16257), .S0 (nx18081)) ;
    mux21 ix14215 (.Y (nx14214), .A0 (nx18151), .A1 (nx16262), .S0 (nx18083)) ;
    mux21 ix14195 (.Y (nx14194), .A0 (nx18151), .A1 (nx16267), .S0 (nx17575)) ;
    mux21 ix14185 (.Y (nx14184), .A0 (nx18151), .A1 (nx16271), .S0 (nx17579)) ;
    mux21 ix14165 (.Y (nx14164), .A0 (nx18063), .A1 (nx16281), .S0 (nx18085)) ;
    mux21 ix14115 (.Y (nx14114), .A0 (nx18063), .A1 (nx16302), .S0 (nx18087)) ;
    mux21 ix14105 (.Y (nx14104), .A0 (nx18063), .A1 (nx16313), .S0 (nx17591)) ;
    mux21 ix14025 (.Y (nx14024), .A0 (nx18063), .A1 (nx16336), .S0 (nx18089)) ;
    mux21 ix14045 (.Y (nx14044), .A0 (nx18063), .A1 (nx16344), .S0 (nx18091)) ;
    mux21 ix14455 (.Y (nx14454), .A0 (nx18155), .A1 (nx16353), .S0 (nx17565)) ;
    mux21 ix14475 (.Y (nx14474), .A0 (nx18155), .A1 (nx16359), .S0 (nx18081)) ;
    mux21 ix14445 (.Y (nx14444), .A0 (nx18155), .A1 (nx16364), .S0 (nx18083)) ;
    mux21 ix14425 (.Y (nx14424), .A0 (nx18155), .A1 (nx16369), .S0 (nx17575)) ;
    mux21 ix14415 (.Y (nx14414), .A0 (nx18155), .A1 (nx16373), .S0 (nx17579)) ;
    mux21 ix14395 (.Y (nx14394), .A0 (nx18065), .A1 (nx16383), .S0 (nx18085)) ;
    mux21 ix14345 (.Y (nx14344), .A0 (nx18065), .A1 (nx16404), .S0 (nx18087)) ;
    mux21 ix14335 (.Y (nx14334), .A0 (nx18065), .A1 (nx16415), .S0 (nx17591)) ;
    mux21 ix14255 (.Y (nx14254), .A0 (nx18065), .A1 (nx16438), .S0 (nx18089)) ;
    mux21 ix14275 (.Y (nx14274), .A0 (nx18065), .A1 (nx16446), .S0 (nx18091)) ;
    mux21 ix14685 (.Y (nx14684), .A0 (nx18159), .A1 (nx16455), .S0 (nx17565)) ;
    mux21 ix14705 (.Y (nx14704), .A0 (nx18159), .A1 (nx16461), .S0 (nx18081)) ;
    mux21 ix14675 (.Y (nx14674), .A0 (nx18159), .A1 (nx16466), .S0 (nx18083)) ;
    mux21 ix14655 (.Y (nx14654), .A0 (nx18159), .A1 (nx16471), .S0 (nx17575)) ;
    mux21 ix14645 (.Y (nx14644), .A0 (nx18159), .A1 (nx16475), .S0 (nx17579)) ;
    mux21 ix14625 (.Y (nx14624), .A0 (nx18067), .A1 (nx16485), .S0 (nx18085)) ;
    mux21 ix14575 (.Y (nx14574), .A0 (nx18067), .A1 (nx16506), .S0 (nx18087)) ;
    mux21 ix14565 (.Y (nx14564), .A0 (nx18067), .A1 (nx16517), .S0 (nx17591)) ;
    mux21 ix14485 (.Y (nx14484), .A0 (nx18067), .A1 (nx16540), .S0 (nx18089)) ;
    mux21 ix14505 (.Y (nx14504), .A0 (nx18067), .A1 (nx16548), .S0 (nx18091)) ;
    mux21 ix14915 (.Y (nx14914), .A0 (nx18163), .A1 (nx16557), .S0 (nx17565)) ;
    mux21 ix14935 (.Y (nx14934), .A0 (nx18163), .A1 (nx16563), .S0 (nx18081)) ;
    mux21 ix14905 (.Y (nx14904), .A0 (nx18163), .A1 (nx16568), .S0 (nx18083)) ;
    mux21 ix14885 (.Y (nx14884), .A0 (nx18163), .A1 (nx16573), .S0 (nx17575)) ;
    mux21 ix14875 (.Y (nx14874), .A0 (nx18163), .A1 (nx16577), .S0 (nx17579)) ;
    mux21 ix14855 (.Y (nx14854), .A0 (nx18069), .A1 (nx16587), .S0 (nx18085)) ;
    mux21 ix14805 (.Y (nx14804), .A0 (nx18069), .A1 (nx16608), .S0 (nx18087)) ;
    mux21 ix14795 (.Y (nx14794), .A0 (nx18069), .A1 (nx16619), .S0 (nx17591)) ;
    mux21 ix14715 (.Y (nx14714), .A0 (nx18069), .A1 (nx16642), .S0 (nx18089)) ;
    mux21 ix14735 (.Y (nx14734), .A0 (nx18069), .A1 (nx16650), .S0 (nx18091)) ;
    mux21 ix15145 (.Y (nx15144), .A0 (nx18167), .A1 (nx16659), .S0 (nx17567)) ;
    mux21 ix15165 (.Y (nx15164), .A0 (nx18167), .A1 (nx16665), .S0 (nx18093)) ;
    inv01 ix18092 (.Y (nx18093), .A (nx17449)) ;
    mux21 ix15135 (.Y (nx15134), .A0 (nx18167), .A1 (nx16670), .S0 (nx18095)) ;
    inv01 ix18094 (.Y (nx18095), .A (nx17439)) ;
    mux21 ix15115 (.Y (nx15114), .A0 (nx18167), .A1 (nx16675), .S0 (nx17577)) ;
    mux21 ix15105 (.Y (nx15104), .A0 (nx18167), .A1 (nx16679), .S0 (nx17581)) ;
    mux21 ix15085 (.Y (nx15084), .A0 (nx18071), .A1 (nx16689), .S0 (nx18097)) ;
    inv01 ix18096 (.Y (nx18097), .A (nx17427)) ;
    mux21 ix15035 (.Y (nx15034), .A0 (nx18071), .A1 (nx16710), .S0 (nx18099)) ;
    inv01 ix18098 (.Y (nx18099), .A (nx17411)) ;
    mux21 ix15025 (.Y (nx15024), .A0 (nx18071), .A1 (nx16721), .S0 (nx17593)) ;
    mux21 ix14945 (.Y (nx14944), .A0 (nx18071), .A1 (nx16744), .S0 (nx18101)) ;
    inv01 ix18100 (.Y (nx18101), .A (nx17377)) ;
    mux21 ix14965 (.Y (nx14964), .A0 (nx18071), .A1 (nx16752), .S0 (nx18103)) ;
    inv01 ix18102 (.Y (nx18103), .A (nx17387)) ;
    nor02_2x ix5621 (.Y (nx5620), .A0 (nx18123), .A1 (nx18105)) ;
    nand03 ix5603 (.Y (nx18105), .A0 (nx17669), .A1 (Address[1]), .A2 (
           Address[2])) ;
    nor02_2x ix5513 (.Y (nx5512), .A0 (nx18123), .A1 (nx18107)) ;
    inv01 ix18106 (.Y (nx18107), .A (nx5502)) ;
    oai221 ix505 (.Y (nx504), .A0 (nx18131), .A1 (nx15192), .B0 (nx422), .B1 (
           nx15226), .C0 (nx18109)) ;
    inv01 ix18108 (.Y (nx18109), .A (nx17665)) ;
    nand03 ix15222 (.Y (nx17541), .A0 (WR), .A1 (nx15188), .A2 (Address[2])) ;
    nor02_2x ix335 (.Y (nx334), .A0 (Address[6]), .A1 (nx18131)) ;
    nor02_2x ix129 (.Y (nx128), .A0 (Address[6]), .A1 (nx15286)) ;
    nor02_2x ix91 (.Y (nx90), .A0 (Address[6]), .A1 (nx18133)) ;
    nand03 ix15300 (.Y (nx17559), .A0 (WR), .A1 (Address[3]), .A2 (nx17533)) ;
    oai221 ix1163 (.Y (nx1162), .A0 (nx422), .A1 (nx15596), .B0 (nx18133), .B1 (
           nx15192), .C0 (nx15598)) ;
    nor02_2x ix1951 (.Y (nx1950), .A0 (nx15708), .A1 (nx18119)) ;
    nor02_2x ix1473 (.Y (nx1472), .A0 (nx18111), .A1 (nx18131)) ;
    inv01 ix18110 (.Y (nx18111), .A (Address[6])) ;
    nor02_2x ix2615 (.Y (nx2614), .A0 (nx15769), .A1 (nx18119)) ;
    nor02_2x ix1489 (.Y (nx1488), .A0 (nx15708), .A1 (nx18129)) ;
    nor02_2x ix2459 (.Y (nx2458), .A0 (nx18129), .A1 (nx18113)) ;
    inv01 ix18112 (.Y (nx18113), .A (nx1558)) ;
    nor02_2x ix2299 (.Y (nx2298), .A0 (nx15769), .A1 (nx18129)) ;
    nor02_2x ix2337 (.Y (nx2336), .A0 (nx18119), .A1 (nx18115)) ;
    inv01 ix18114 (.Y (nx18115), .A (nx2216)) ;
    nor02_2x ix2221 (.Y (nx2220), .A0 (nx18129), .A1 (nx18115)) ;
    nor02_2x ix2161 (.Y (nx2160), .A0 (nx15881), .A1 (nx18119)) ;
    nor02_2x ix2057 (.Y (nx2056), .A0 (nx15720), .A1 (nx18121)) ;
    nor02_2x ix1595 (.Y (nx1594), .A0 (nx18111), .A1 (nx18133)) ;
    nor02_2x ix2011 (.Y (nx2010), .A0 (nx15720), .A1 (nx18129)) ;
    nor02_2x ix1917 (.Y (nx1916), .A0 (nx15881), .A1 (nx17343)) ;
    nor02_2x ix1835 (.Y (nx1834), .A0 (nx15744), .A1 (nx18121)) ;
    nor02_2x ix1795 (.Y (nx1794), .A0 (nx15744), .A1 (nx17343)) ;
    nor03_2x ix1559 (.Y (nx1558), .A0 (nx18117), .A1 (nx15746), .A2 (nx1552)) ;
    inv01 ix18116 (.Y (nx18117), .A (nx1540)) ;
    nor02_2x ix5713 (.Y (nx5712), .A0 (nx17072), .A1 (nx18123)) ;
    nor02_2x ix5705 (.Y (nx5704), .A0 (nx17075), .A1 (nx18123)) ;
    nor02_2x ix5697 (.Y (nx5696), .A0 (nx17072), .A1 (nx18125)) ;
    nor02_2x ix5693 (.Y (nx5692), .A0 (nx18125), .A1 (nx18107)) ;
    nor02_2x ix5673 (.Y (nx5672), .A0 (nx17075), .A1 (nx18135)) ;
    nor02_2x ix5669 (.Y (nx5668), .A0 (nx17075), .A1 (nx18125)) ;
    nor02_2x ix5657 (.Y (nx5656), .A0 (nx17106), .A1 (nx18123)) ;
    nor02_2x ix5653 (.Y (nx5652), .A0 (nx17109), .A1 (nx17067)) ;
    nor02_2x ix5625 (.Y (nx5624), .A0 (nx17106), .A1 (nx18135)) ;
    nor02_2x ix5617 (.Y (nx5616), .A0 (nx17109), .A1 (nx18135)) ;
    nor04 ix5605 (.Y (nx5604), .A0 (nx18125), .A1 (Address[0]), .A2 (nx17545), .A3 (
          nx17533)) ;
    nor04 ix5609 (.Y (nx5608), .A0 (nx18135), .A1 (Address[0]), .A2 (nx17545), .A3 (
          nx17533)) ;
    nor02_2x ix5583 (.Y (nx5582), .A0 (nx17109), .A1 (nx18127)) ;
    nor02_2x ix5593 (.Y (nx5592), .A0 (nx17072), .A1 (nx18135)) ;
    nor02_2x ix5563 (.Y (nx5562), .A0 (nx17106), .A1 (nx18127)) ;
    nor02_2x ix5505 (.Y (nx5504), .A0 (nx17645), .A1 (nx18107)) ;
    nor02_2x ix17400 (.Y (nx17401), .A0 (nx15881), .A1 (nx17343)) ;
    nor02_2x ix17450 (.Y (nx17451), .A0 (nx15769), .A1 (nx18121)) ;
    nor02_2x ix17502 (.Y (nx17503), .A0 (nx17109), .A1 (nx17645)) ;
    nor02_2x ix17516 (.Y (nx17517), .A0 (nx17075), .A1 (nx18127)) ;
    nor02_2x ix17522 (.Y (nx17523), .A0 (nx17075), .A1 (nx17067)) ;
    inv01 ix18118 (.Y (nx18119), .A (nx17829)) ;
    inv01 ix18120 (.Y (nx18121), .A (nx17829)) ;
    inv02 ix18122 (.Y (nx18123), .A (nx5510)) ;
    inv01 ix18124 (.Y (nx18125), .A (nx17787)) ;
    inv01 ix18126 (.Y (nx18127), .A (nx17787)) ;
    inv02 ix18128 (.Y (nx18129), .A (nx15308)) ;
    inv02 ix18130 (.Y (nx18131), .A (nx17675)) ;
    inv02 ix18132 (.Y (nx18133), .A (nx17671)) ;
    inv02 ix18134 (.Y (nx18135), .A (nx5496)) ;
    inv01 ix18136 (.Y (nx18137), .A (Din[0])) ;
    inv01 ix18138 (.Y (nx18139), .A (Din[0])) ;
    inv01 ix18140 (.Y (nx18141), .A (Din[1])) ;
    inv01 ix18142 (.Y (nx18143), .A (Din[1])) ;
    inv01 ix18144 (.Y (nx18145), .A (Din[2])) ;
    inv01 ix18146 (.Y (nx18147), .A (Din[2])) ;
    inv01 ix18148 (.Y (nx18149), .A (Din[3])) ;
    inv01 ix18150 (.Y (nx18151), .A (Din[3])) ;
    inv01 ix18152 (.Y (nx18153), .A (Din[4])) ;
    inv01 ix18154 (.Y (nx18155), .A (Din[4])) ;
    inv01 ix18156 (.Y (nx18157), .A (Din[5])) ;
    inv01 ix18158 (.Y (nx18159), .A (Din[5])) ;
    inv01 ix18160 (.Y (nx18161), .A (Din[6])) ;
    inv01 ix18162 (.Y (nx18163), .A (Din[6])) ;
    inv01 ix18164 (.Y (nx18165), .A (Din[7])) ;
    inv01 ix18166 (.Y (nx18167), .A (Din[7])) ;
endmodule

