LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

PACKAGE common IS

    TYPE matrix_byte IS
    ARRAY(NATURAL RANGE<>, NATURAL RANGE<>) OF STD_LOGIC_VECTOR(7 DOWNTO 0);

    TYPE matrix_bit IS
    ARRAY(NATURAL RANGE<>, NATURAL RANGE<>) OF STD_LOGIC;

    TYPE array_clen IS
    ARRAY(NATURAL RANGE<>) OF STD_LOGIC_VECTOR(18 DOWNTO 0);

    TYPE array_byte IS
    ARRAY(NATURAL RANGE<>) OF STD_LOGIC_VECTOR(7 DOWNTO 0);

END PACKAGE;