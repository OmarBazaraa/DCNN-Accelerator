//
// Verilog description for cell RAM, 
// Wed May  9 07:36:13 2018
//
// LeonardoSpectrum Level 3, 2017a.2 
//


module RAM ( CLK, WR, Address, Din, Dout ) ;

    input CLK ;
    input WR ;
    input [4:0]Address ;
    input [7:0]Din ;
    output [39:0]Dout ;

    wire Mem_24__0, nx14, Mem_25__0, nx32, nx42, Mem_26__0, nx54, Mem_27__0, 
         nx66, nx68, nx78, nx82, nx88, nx104, Mem_4__0, nx116, nx122, Mem_5__0, 
         nx136, nx146, Mem_6__0, nx154, Mem_7__0, nx166, nx176, nx180, nx190, 
         Mem_16__0, nx202, Mem_17__0, nx216, nx226, Mem_18__0, nx234, Mem_19__0, 
         nx246, nx256, nx260, nx266, Mem_12__0, nx274, Mem_13__0, nx298, 
         Mem_14__0, nx306, Mem_15__0, nx318, nx328, nx332, nx340, Mem_8__0, 
         nx352, nx358, Mem_9__0, nx372, nx382, Mem_10__0, nx390, Mem_11__0, 
         nx402, nx412, nx416, nx422, Mem_20__0, nx428, Mem_21__0, nx456, 
         Mem_22__0, Mem_23__0, nx486, nx490, nx498, Mem_28__0, nx502, Mem_29__0, 
         nx530, Mem_30__0, Mem_31__0, nx560, nx564, nx570, Mem_24__1, Mem_25__1, 
         nx598, Mem_26__1, Mem_27__1, nx622, nx626, Mem_4__1, Mem_5__1, nx648, 
         Mem_6__1, Mem_7__1, nx672, nx676, Mem_16__1, Mem_17__1, nx700, 
         Mem_18__1, Mem_19__1, nx724, nx728, Mem_12__1, Mem_13__1, nx750, 
         Mem_14__1, Mem_15__1, nx774, nx778, Mem_8__1, Mem_9__1, nx804, 
         Mem_10__1, Mem_11__1, nx828, nx832, Mem_20__1, Mem_21__1, nx854, 
         Mem_22__1, Mem_23__1, nx878, nx882, Mem_28__1, Mem_29__1, nx904, 
         Mem_30__1, Mem_31__1, nx928, nx932, Mem_24__2, Mem_25__2, nx960, 
         Mem_26__2, Mem_27__2, nx984, nx988, Mem_4__2, Mem_5__2, nx1010, 
         Mem_6__2, Mem_7__2, nx1034, nx1038, Mem_16__2, Mem_17__2, nx1062, 
         Mem_18__2, Mem_19__2, nx1086, nx1090, Mem_12__2, Mem_13__2, nx1112, 
         Mem_14__2, Mem_15__2, nx1136, nx1140, Mem_8__2, Mem_9__2, nx1166, 
         Mem_10__2, Mem_11__2, nx1190, nx1194, Mem_20__2, Mem_21__2, nx1216, 
         Mem_22__2, Mem_23__2, nx1240, nx1244, Mem_28__2, Mem_29__2, nx1266, 
         Mem_30__2, Mem_31__2, nx1290, nx1294, Mem_24__3, Mem_25__3, nx1322, 
         Mem_26__3, Mem_27__3, nx1346, nx1350, Mem_4__3, Mem_5__3, nx1372, 
         Mem_6__3, Mem_7__3, nx1396, nx1400, Mem_16__3, Mem_17__3, nx1424, 
         Mem_18__3, Mem_19__3, nx1448, nx1452, Mem_12__3, Mem_13__3, nx1474, 
         Mem_14__3, Mem_15__3, nx1498, nx1502, Mem_8__3, Mem_9__3, nx1528, 
         Mem_10__3, Mem_11__3, nx1552, nx1556, Mem_20__3, Mem_21__3, nx1578, 
         Mem_22__3, Mem_23__3, nx1602, nx1606, Mem_28__3, Mem_29__3, nx1628, 
         Mem_30__3, Mem_31__3, nx1652, nx1656, Mem_24__4, Mem_25__4, nx1684, 
         Mem_26__4, Mem_27__4, nx1708, nx1712, Mem_4__4, Mem_5__4, nx1734, 
         Mem_6__4, Mem_7__4, nx1758, nx1762, Mem_16__4, Mem_17__4, nx1786, 
         Mem_18__4, Mem_19__4, nx1810, nx1814, Mem_12__4, Mem_13__4, nx1836, 
         Mem_14__4, Mem_15__4, nx1860, nx1864, Mem_8__4, Mem_9__4, nx1890, 
         Mem_10__4, Mem_11__4, nx1914, nx1918, Mem_20__4, Mem_21__4, nx1940, 
         Mem_22__4, Mem_23__4, nx1964, nx1968, Mem_28__4, Mem_29__4, nx1990, 
         Mem_30__4, Mem_31__4, nx2014, nx2018, Mem_24__5, Mem_25__5, nx2046, 
         Mem_26__5, Mem_27__5, nx2070, nx2074, Mem_4__5, Mem_5__5, nx2096, 
         Mem_6__5, Mem_7__5, nx2120, nx2124, Mem_16__5, Mem_17__5, nx2148, 
         Mem_18__5, Mem_19__5, nx2172, nx2176, Mem_12__5, Mem_13__5, nx2198, 
         Mem_14__5, Mem_15__5, nx2222, nx2226, Mem_8__5, Mem_9__5, nx2252, 
         Mem_10__5, Mem_11__5, nx2276, nx2280, Mem_20__5, Mem_21__5, nx2302, 
         Mem_22__5, Mem_23__5, nx2326, nx2330, Mem_28__5, Mem_29__5, nx2352, 
         Mem_30__5, Mem_31__5, nx2376, nx2380, Mem_24__6, Mem_25__6, nx2408, 
         Mem_26__6, Mem_27__6, nx2432, nx2436, Mem_4__6, Mem_5__6, nx2458, 
         Mem_6__6, Mem_7__6, nx2482, nx2486, Mem_16__6, Mem_17__6, nx2510, 
         Mem_18__6, Mem_19__6, nx2534, nx2538, Mem_12__6, Mem_13__6, nx2560, 
         Mem_14__6, Mem_15__6, nx2584, nx2588, Mem_8__6, Mem_9__6, nx2614, 
         Mem_10__6, Mem_11__6, nx2638, nx2642, Mem_20__6, Mem_21__6, nx2664, 
         Mem_22__6, Mem_23__6, nx2688, nx2692, Mem_28__6, Mem_29__6, nx2714, 
         Mem_30__6, Mem_31__6, nx2738, nx2742, Mem_24__7, Mem_25__7, nx2770, 
         Mem_26__7, Mem_27__7, nx2794, nx2798, Mem_4__7, Mem_5__7, nx2820, 
         Mem_6__7, Mem_7__7, nx2844, nx2848, Mem_16__7, Mem_17__7, nx2872, 
         Mem_18__7, Mem_19__7, nx2896, nx2900, Mem_12__7, Mem_13__7, nx2922, 
         Mem_14__7, Mem_15__7, nx2946, nx2950, Mem_8__7, Mem_9__7, nx2976, 
         Mem_10__7, Mem_11__7, nx3000, nx3004, Mem_20__7, Mem_21__7, nx3026, 
         Mem_22__7, Mem_23__7, nx3050, nx3054, Mem_28__7, Mem_29__7, nx3076, 
         Mem_30__7, Mem_31__7, nx3100, nx3104, nx3120, nx3122, nx3126, nx3136, 
         nx3148, nx3152, nx3162, nx3172, nx3184, nx3188, nx3194, nx3204, nx3210, 
         nx3224, nx3232, nx3242, nx3248, nx3260, nx3262, nx3272, nx3278, nx3294, 
         nx3300, Mem_3__0, nx3308, nx3330, nx3342, nx3344, nx3354, nx3362, 
         nx3376, nx3382, nx3392, nx3396, nx3406, nx3414, nx3432, nx3442, nx3454, 
         nx3464, nx3478, nx3488, nx3500, nx3510, nx3526, Mem_3__1, nx3546, 
         nx3556, nx3570, nx3580, nx3590, nx3608, nx3618, nx3630, nx3640, nx3654, 
         nx3664, nx3676, nx3686, nx3702, Mem_3__2, nx3722, nx3732, nx3746, 
         nx3756, nx3766, nx3784, nx3794, nx3806, nx3816, nx3830, nx3840, nx3852, 
         nx3862, nx3878, Mem_3__3, nx3898, nx3908, nx3922, nx3932, nx3942, 
         nx3960, nx3970, nx3982, nx3992, nx4006, nx4016, nx4028, nx4038, nx4054, 
         Mem_3__4, nx4074, nx4084, nx4098, nx4108, nx4118, nx4136, nx4146, 
         nx4158, nx4168, nx4182, nx4192, nx4204, nx4214, nx4230, Mem_3__5, 
         nx4250, nx4260, nx4274, nx4284, nx4294, nx4312, nx4322, nx4334, nx4344, 
         nx4358, nx4368, nx4380, nx4390, nx4406, Mem_3__6, nx4426, nx4436, 
         nx4450, nx4460, nx4470, nx4488, nx4498, nx4510, nx4520, nx4534, nx4544, 
         nx4556, nx4566, nx4582, Mem_3__7, nx4602, nx4612, nx4626, nx4636, 
         nx4646, Mem_2__0, nx4676, nx4708, nx4716, nx4724, nx4730, nx4742, 
         nx4752, nx4764, nx4768, nx4782, nx4792, nx4798, nx4806, nx4814, nx4822, 
         nx4830, Mem_2__1, nx4854, Mem_2__2, nx4926, Mem_2__3, nx4998, Mem_2__4, 
         nx5070, Mem_2__5, nx5142, Mem_2__6, nx5214, Mem_2__7, nx5286, nx5346, 
         nx5352, nx5364, nx5366, nx5372, nx5382, nx5390, nx5406, nx5412, nx5418, 
         nx5428, nx5434, nx5440, nx5450, nx5458, nx5466, nx5472, nx5478, 
         Mem_1__0, nx5486, nx5506, nx5512, nx5520, nx5526, nx5538, nx5542, 
         nx5550, nx5586, Mem_1__1, nx5622, nx5658, Mem_1__2, nx5694, nx5730, 
         Mem_1__3, nx5766, nx5802, Mem_1__4, nx5838, nx5874, Mem_1__5, nx5910, 
         nx5946, Mem_1__6, nx5982, nx6018, Mem_1__7, nx6054, nx6058, nx6064, 
         nx6070, nx6080, nx6084, Mem_0__0, nx6098, Mem_0__1, Mem_0__2, Mem_0__3, 
         Mem_0__4, Mem_0__5, Mem_0__6, Mem_0__7, nx4375, nx4385, nx4395, nx4405, 
         nx4415, nx4425, nx4435, nx4445, nx4455, nx4465, nx4475, nx4485, nx4495, 
         nx4505, nx4515, nx4525, nx4535, nx4545, nx4555, nx4565, nx4575, nx4585, 
         nx4595, nx4605, nx4615, nx4625, nx4635, nx4645, nx4655, nx4665, nx4675, 
         nx4685, nx4695, nx4705, nx4715, nx4725, nx4735, nx4745, nx4755, nx4765, 
         nx4775, nx4785, nx4795, nx4805, nx4815, nx4825, nx4835, nx4845, nx4855, 
         nx4865, nx4875, nx4885, nx4895, nx4905, nx4915, nx4925, nx4935, nx4945, 
         nx4955, nx4965, nx4975, nx4985, nx4995, nx5005, nx5015, nx5025, nx5035, 
         nx5045, nx5055, nx5065, nx5075, nx5085, nx5095, nx5105, nx5115, nx5125, 
         nx5135, nx5145, nx5155, nx5165, nx5175, nx5185, nx5195, nx5205, nx5215, 
         nx5225, nx5235, nx5245, nx5255, nx5265, nx5275, nx5285, nx5295, nx5305, 
         nx5315, nx5325, nx5335, nx5345, nx5355, nx5365, nx5375, nx5385, nx5395, 
         nx5405, nx5415, nx5425, nx5435, nx5445, nx5455, nx5465, nx5475, nx5485, 
         nx5495, nx5505, nx5515, nx5525, nx5535, nx5545, nx5555, nx5565, nx5575, 
         nx5585, nx5595, nx5605, nx5615, nx5625, nx5635, nx5645, nx5655, nx5665, 
         nx5675, nx5685, nx5695, nx5705, nx5715, nx5725, nx5735, nx5745, nx5755, 
         nx5765, nx5775, nx5785, nx5795, nx5805, nx5815, nx5825, nx5835, nx5845, 
         nx5855, nx5865, nx5875, nx5885, nx5895, nx5905, nx5915, nx5925, nx5935, 
         nx5945, nx5955, nx5965, nx5975, nx5985, nx5995, nx6005, nx6015, nx6025, 
         nx6035, nx6045, nx6055, nx6065, nx6075, nx6085, nx6095, nx6105, nx6115, 
         nx6125, nx6135, nx6145, nx6155, nx6165, nx6175, nx6185, nx6195, nx6205, 
         nx6215, nx6225, nx6235, nx6245, nx6255, nx6265, nx6275, nx6285, nx6295, 
         nx6305, nx6315, nx6325, nx6335, nx6345, nx6355, nx6365, nx6375, nx6385, 
         nx6395, nx6405, nx6415, nx6425, nx6435, nx6445, nx6455, nx6465, nx6475, 
         nx6485, nx6495, nx6505, nx6515, nx6525, nx6535, nx6545, nx6555, nx6565, 
         nx6575, nx6585, nx6595, nx6605, nx6615, nx6625, nx6635, nx6645, nx6655, 
         nx6665, nx6675, nx6685, nx6695, nx6705, nx6715, nx6725, nx6735, nx6745, 
         nx6755, nx6765, nx6775, nx6785, nx6795, nx6805, nx6815, nx6825, nx6835, 
         nx6845, nx6855, nx6865, nx6875, nx6885, nx6895, nx6905, nx6915, nx6925, 
         nx6936, nx6942, nx6944, nx6947, nx6949, nx6954, nx6956, nx6958, nx6964, 
         nx6966, nx6973, nx6986, nx6994, nx7000, nx7005, nx7015, nx7033, nx7037, 
         nx7044, nx7050, nx7068, nx7070, nx7087, nx7094, nx7117, nx7135, nx7182, 
         nx7214, nx7247, nx7294, nx7326, nx7359, nx7406, nx7438, nx7471, nx7518, 
         nx7550, nx7583, nx7630, nx7662, nx7695, nx7742, nx7774, nx7807, nx7854, 
         nx7886, nx7919, nx7926, nx7929, nx7934, nx7939, nx7941, nx7945, nx7947, 
         nx7951, nx7955, nx7957, nx7963, nx7968, nx7970, nx7972, nx7979, nx7985, 
         nx7991, nx7998, nx8003, nx8007, nx8013, nx8015, nx8019, nx8023, nx8027, 
         nx8032, nx8037, nx8041, nx8047, nx8049, nx8053, nx8057, nx8061, nx8066, 
         nx8071, nx8075, nx8081, nx8083, nx8087, nx8091, nx8095, nx8100, nx8105, 
         nx8109, nx8115, nx8117, nx8121, nx8125, nx8129, nx8134, nx8139, nx8143, 
         nx8149, nx8151, nx8155, nx8159, nx8163, nx8168, nx8173, nx8177, nx8183, 
         nx8185, nx8189, nx8193, nx8197, nx8202, nx8207, nx8211, nx8217, nx8219, 
         nx8223, nx8227, nx8231, nx8236, nx8241, nx8245, nx8249, nx8251, nx8255, 
         nx8259, nx8263, nx8269, nx8274, nx8276, nx8278, nx8280, nx8282, nx8284, 
         nx8286, nx8288, nx8295, nx8297, nx8299, nx8301, nx8303, nx8305, nx8307, 
         nx8309, nx8316, nx8318, nx8320, nx8322, nx8324, nx8326, nx8328, nx8330, 
         nx8337, nx8339, nx8341, nx8343, nx8345, nx8347, nx8349, nx8351, nx8358, 
         nx8360, nx8362, nx8364, nx8366, nx8368, nx8370, nx8372, nx8379, nx8381, 
         nx8383, nx8385, nx8387, nx8389, nx8391, nx8393, nx8400, nx8402, nx8404, 
         nx8406, nx8408, nx8410, nx8412, nx8414, nx8422, nx8427, nx8432, nx8435, 
         nx8437, nx8442, nx8445, nx8448, nx8450, nx8452, nx8456, nx8463, nx8466, 
         nx8471, nx8475, nx8478, nx8481, nx8485, nx8492, nx8494, nx8496, nx8501, 
         nx8504, nx8506, nx8508, nx8510, nx8514, nx8516, nx8518, nx8523, nx8526, 
         nx8528, nx8530, nx8532, nx8536, nx8538, nx8540, nx8545, nx8548, nx8550, 
         nx8552, nx8554, nx8558, nx8560, nx8562, nx8567, nx8570, nx8572, nx8574, 
         nx8576, nx8580, nx8582, nx8584, nx8589, nx8592, nx8594, nx8596, nx8598, 
         nx8602, nx8604, nx8606, nx8611, nx8614, nx8616, nx8618, nx8620, nx8624, 
         nx8626, nx8628, nx8633, nx8636, nx8638, nx8640, nx8642, nx8645, nx8647, 
         nx8651, nx8655, nx8659, nx8665, nx8667, nx8672, nx8674, nx8677, nx8679, 
         nx8684, nx8686, nx8689, nx8691, nx8696, nx8698, nx8701, nx8703, nx8708, 
         nx8710, nx8713, nx8715, nx8720, nx8722, nx8725, nx8727, nx8732, nx8734, 
         nx8737, nx8739, nx8744, nx8746, nx8753, nx8755, nx8757, nx8759, nx8761, 
         nx8763, nx8765, nx8767, nx8769, nx8771, nx8773, nx8775, nx8777, nx8779, 
         nx8781, nx8783, nx8785, nx8787, nx8789, nx8791, nx8793, nx8795, nx8797, 
         nx8799, nx8801, nx8803, nx8805, nx8807, nx8809, nx8811, nx8813, nx8815, 
         nx8817, nx8819, nx8821, nx8823, nx8825, nx8827, nx8829, nx8831, nx8833, 
         nx8835, nx8837, nx8839, nx8841, nx8843, nx8845, nx8847, nx8849, nx8851, 
         nx8853, nx8855, nx8857, nx8859, nx8861, nx8863, nx8865, nx8867, nx8869, 
         nx8871, nx8873, nx8875, nx8877, nx8879, nx8881, nx8883, nx8885, nx8887, 
         nx8889, nx8891, nx8893, nx8895, nx8897, nx8899, nx8901, nx8903, nx8905, 
         nx8907, nx8909, nx8911, nx8913, nx8915, nx8917, nx8919, nx8921, nx8923, 
         nx8925, nx8927, nx8929, nx8931, nx8933, nx8935, nx8937, nx8939, nx8941, 
         nx8943, nx8945, nx8947, nx8949, nx8951, nx8955, nx8957, nx8959, nx8961, 
         nx8963, nx8965, nx8967, nx8969, nx8971, nx8973, nx8975, nx8977, nx8979, 
         nx8981, nx8983, nx8985, nx8987, nx8989, nx8991, nx8993, nx8997, nx8999, 
         nx9001, nx9003, nx9005, nx9007, nx9009, nx9011, nx9013, nx9015, nx9017, 
         nx9019, nx9021, nx9023, nx9025, nx9027, nx9029, nx9031, nx9049, nx9051, 
         nx9053, nx9055, nx9057, nx9059, nx9061, nx9063, nx9065, nx9067, nx9069, 
         nx9071, nx9073, nx9075, nx9077, nx9079, nx9081, nx9083, nx9085, nx9087, 
         nx9089, nx9091, nx9093, nx9095, nx9097, nx9099, nx9101, nx9103, nx9105, 
         nx9107, nx9109, nx9111, nx9113, nx9115, nx9117, nx9119, nx9121, nx9123, 
         nx9125;
    wire [255:0] \$dummy ;




    nand03 ix579 (.Y (Dout[0]), .A0 (nx6936), .A1 (nx7037), .A2 (nx7087)) ;
    aoi222 ix6937 (.Y (nx6936), .A0 (nx564), .A1 (nx8809), .B0 (nx490), .B1 (
           nx8805), .C0 (nx416), .C1 (nx8801)) ;
    mux21_ni ix565 (.Y (nx564), .A0 (nx530), .A1 (nx560), .S0 (Address[1])) ;
    mux21_ni ix531 (.Y (nx530), .A0 (Mem_28__0), .A1 (Mem_29__0), .S0 (
             Address[0])) ;
    dff reg_Mem_28__0 (.Q (Mem_28__0), .QB (\$dummy [0]), .D (nx4615), .CLK (CLK
        )) ;
    mux21_ni ix4616 (.Y (nx4615), .A0 (Din[0]), .A1 (Mem_28__0), .S0 (nx8939)) ;
    nand02 ix6943 (.Y (nx6942), .A0 (nx9067), .A1 (nx502)) ;
    nor02_2x ix6945 (.Y (nx6944), .A0 (Address[1]), .A1 (Address[0])) ;
    nor02_2x ix503 (.Y (nx502), .A0 (nx6947), .A1 (nx6949)) ;
    nand02 ix6948 (.Y (nx6947), .A0 (Address[3]), .A1 (Address[2])) ;
    nand02 ix6950 (.Y (nx6949), .A0 (Address[4]), .A1 (WR)) ;
    dff reg_Mem_29__0 (.Q (Mem_29__0), .QB (\$dummy [1]), .D (nx4625), .CLK (CLK
        )) ;
    mux21_ni ix4626 (.Y (nx4625), .A0 (Din[0]), .A1 (Mem_29__0), .S0 (nx8943)) ;
    nand02 ix6955 (.Y (nx6954), .A0 (nx9071), .A1 (nx502)) ;
    inv01 ix6959 (.Y (nx6958), .A (Address[0])) ;
    mux21_ni ix561 (.Y (nx560), .A0 (Mem_30__0), .A1 (Mem_31__0), .S0 (
             Address[0])) ;
    dff reg_Mem_30__0 (.Q (Mem_30__0), .QB (\$dummy [2]), .D (nx4635), .CLK (CLK
        )) ;
    mux21_ni ix4636 (.Y (nx4635), .A0 (Din[0]), .A1 (Mem_30__0), .S0 (nx8947)) ;
    nand02 ix6965 (.Y (nx6964), .A0 (nx9075), .A1 (nx502)) ;
    dff reg_Mem_31__0 (.Q (Mem_31__0), .QB (\$dummy [3]), .D (nx4645), .CLK (CLK
        )) ;
    mux21_ni ix4646 (.Y (nx4645), .A0 (Din[0]), .A1 (Mem_31__0), .S0 (nx8955)) ;
    nand02 ix6974 (.Y (nx6973), .A0 (nx9049), .A1 (nx502)) ;
    nor03_2x ix571 (.Y (nx570), .A0 (nx8959), .A1 (nx8963), .A2 (Address[2])) ;
    mux21_ni ix491 (.Y (nx490), .A0 (nx456), .A1 (nx486), .S0 (Address[1])) ;
    mux21_ni ix457 (.Y (nx456), .A0 (Mem_20__0), .A1 (Mem_21__0), .S0 (
             Address[0])) ;
    dff reg_Mem_20__0 (.Q (Mem_20__0), .QB (\$dummy [4]), .D (nx4575), .CLK (CLK
        )) ;
    mux21_ni ix4576 (.Y (nx4575), .A0 (Din[0]), .A1 (Mem_20__0), .S0 (nx8967)) ;
    nand02 ix6987 (.Y (nx6986), .A0 (nx9067), .A1 (nx428)) ;
    nor03_2x ix429 (.Y (nx428), .A0 (nx8971), .A1 (Address[3]), .A2 (nx6949)) ;
    dff reg_Mem_21__0 (.Q (Mem_21__0), .QB (\$dummy [5]), .D (nx4585), .CLK (CLK
        )) ;
    mux21_ni ix4586 (.Y (nx4585), .A0 (Din[0]), .A1 (Mem_21__0), .S0 (nx8977)) ;
    nand02 ix6995 (.Y (nx6994), .A0 (nx9071), .A1 (nx428)) ;
    mux21_ni ix487 (.Y (nx486), .A0 (Mem_22__0), .A1 (Mem_23__0), .S0 (
             Address[0])) ;
    dff reg_Mem_22__0 (.Q (Mem_22__0), .QB (\$dummy [6]), .D (nx4595), .CLK (CLK
        )) ;
    mux21_ni ix4596 (.Y (nx4595), .A0 (Din[0]), .A1 (Mem_22__0), .S0 (nx8981)) ;
    nand02 ix7001 (.Y (nx7000), .A0 (nx9075), .A1 (nx428)) ;
    dff reg_Mem_23__0 (.Q (Mem_23__0), .QB (\$dummy [7]), .D (nx4605), .CLK (CLK
        )) ;
    mux21_ni ix4606 (.Y (nx4605), .A0 (Din[0]), .A1 (Mem_23__0), .S0 (nx8985)) ;
    nand02 ix7006 (.Y (nx7005), .A0 (nx9049), .A1 (nx428)) ;
    nor03_2x ix499 (.Y (nx498), .A0 (nx8959), .A1 (Address[3]), .A2 (Address[2])
             ) ;
    mux21_ni ix417 (.Y (nx416), .A0 (nx382), .A1 (nx412), .S0 (Address[1])) ;
    mux21_ni ix383 (.Y (nx382), .A0 (Mem_8__0), .A1 (Mem_9__0), .S0 (Address[0])
             ) ;
    dff reg_Mem_8__0 (.Q (Mem_8__0), .QB (\$dummy [8]), .D (nx4535), .CLK (CLK)
        ) ;
    mux21_ni ix4536 (.Y (nx4535), .A0 (Mem_8__0), .A1 (Din[0]), .S0 (nx9115)) ;
    nand02 ix7016 (.Y (nx7015), .A0 (WR), .A1 (nx8789)) ;
    nor03_2x ix353 (.Y (nx352), .A0 (Address[4]), .A1 (Address[2]), .A2 (nx8963)
             ) ;
    dff reg_Mem_9__0 (.Q (Mem_9__0), .QB (\$dummy [9]), .D (nx4545), .CLK (CLK)
        ) ;
    mux21_ni ix4546 (.Y (nx4545), .A0 (Mem_9__0), .A1 (Din[0]), .S0 (nx9117)) ;
    mux21_ni ix413 (.Y (nx412), .A0 (Mem_10__0), .A1 (Mem_11__0), .S0 (
             Address[0])) ;
    dff reg_Mem_10__0 (.Q (Mem_10__0), .QB (\$dummy [10]), .D (nx4555), .CLK (
        CLK)) ;
    mux21_ni ix4556 (.Y (nx4555), .A0 (Mem_10__0), .A1 (Din[0]), .S0 (nx9119)) ;
    dff reg_Mem_11__0 (.Q (Mem_11__0), .QB (\$dummy [11]), .D (nx4565), .CLK (
        CLK)) ;
    mux21_ni ix4566 (.Y (nx4565), .A0 (Mem_11__0), .A1 (Din[0]), .S0 (nx9121)) ;
    nand02 ix7034 (.Y (nx7033), .A0 (Address[0]), .A1 (Address[1])) ;
    nor03_2x ix423 (.Y (nx422), .A0 (Address[4]), .A1 (Address[3]), .A2 (nx8971)
             ) ;
    aoi22 ix7038 (.Y (nx7037), .A0 (nx332), .A1 (nx340), .B0 (nx260), .B1 (nx266
          )) ;
    mux21_ni ix333 (.Y (nx332), .A0 (nx298), .A1 (nx328), .S0 (Address[1])) ;
    mux21_ni ix299 (.Y (nx298), .A0 (Mem_12__0), .A1 (Mem_13__0), .S0 (
             Address[0])) ;
    dff reg_Mem_12__0 (.Q (Mem_12__0), .QB (\$dummy [12]), .D (nx4495), .CLK (
        CLK)) ;
    mux21_ni ix4496 (.Y (nx4495), .A0 (Mem_12__0), .A1 (Din[0]), .S0 (nx9109)) ;
    nand02_2x ix7045 (.Y (nx7044), .A0 (WR), .A1 (nx8761)) ;
    nor02_2x ix89 (.Y (nx88), .A0 (Address[4]), .A1 (nx6947)) ;
    dff reg_Mem_13__0 (.Q (Mem_13__0), .QB (\$dummy [13]), .D (nx4505), .CLK (
        CLK)) ;
    mux21_ni ix4506 (.Y (nx4505), .A0 (Din[0]), .A1 (Mem_13__0), .S0 (nx8997)) ;
    nand03 ix7051 (.Y (nx7050), .A0 (nx9071), .A1 (WR), .A2 (nx8761)) ;
    mux21_ni ix329 (.Y (nx328), .A0 (Mem_14__0), .A1 (Mem_15__0), .S0 (
             Address[0])) ;
    dff reg_Mem_14__0 (.Q (Mem_14__0), .QB (\$dummy [14]), .D (nx4515), .CLK (
        CLK)) ;
    mux21_ni ix4516 (.Y (nx4515), .A0 (Mem_14__0), .A1 (Din[0]), .S0 (nx9111)) ;
    dff reg_Mem_15__0 (.Q (Mem_15__0), .QB (\$dummy [15]), .D (nx4525), .CLK (
        CLK)) ;
    mux21_ni ix4526 (.Y (nx4525), .A0 (Mem_15__0), .A1 (Din[0]), .S0 (nx9113)) ;
    nor03_2x ix341 (.Y (nx340), .A0 (Address[4]), .A1 (nx8963), .A2 (Address[2])
             ) ;
    mux21_ni ix261 (.Y (nx260), .A0 (nx226), .A1 (nx256), .S0 (Address[1])) ;
    mux21_ni ix227 (.Y (nx226), .A0 (Mem_16__0), .A1 (Mem_17__0), .S0 (
             Address[0])) ;
    dff reg_Mem_16__0 (.Q (Mem_16__0), .QB (\$dummy [16]), .D (nx4455), .CLK (
        CLK)) ;
    mux21_ni ix4456 (.Y (nx4455), .A0 (Mem_16__0), .A1 (Din[0]), .S0 (nx9101)) ;
    nand03 ix7069 (.Y (nx7068), .A0 (nx7070), .A1 (Address[4]), .A2 (WR)) ;
    nor02_2x ix7071 (.Y (nx7070), .A0 (Address[2]), .A1 (Address[3])) ;
    dff reg_Mem_17__0 (.Q (Mem_17__0), .QB (\$dummy [17]), .D (nx4465), .CLK (
        CLK)) ;
    mux21_ni ix4466 (.Y (nx4465), .A0 (Mem_17__0), .A1 (Din[0]), .S0 (nx9103)) ;
    mux21_ni ix257 (.Y (nx256), .A0 (Mem_18__0), .A1 (Mem_19__0), .S0 (
             Address[0])) ;
    dff reg_Mem_18__0 (.Q (Mem_18__0), .QB (\$dummy [18]), .D (nx4475), .CLK (
        CLK)) ;
    mux21_ni ix4476 (.Y (nx4475), .A0 (Mem_18__0), .A1 (Din[0]), .S0 (nx9105)) ;
    dff reg_Mem_19__0 (.Q (Mem_19__0), .QB (\$dummy [19]), .D (nx4485), .CLK (
        CLK)) ;
    mux21_ni ix4486 (.Y (nx4485), .A0 (Mem_19__0), .A1 (Din[0]), .S0 (nx9107)) ;
    nor03_2x ix267 (.Y (nx266), .A0 (Address[4]), .A1 (nx8963), .A2 (nx8971)) ;
    aoi22 ix7088 (.Y (nx7087), .A0 (nx180), .A1 (nx190), .B0 (nx82), .B1 (nx104)
          ) ;
    mux21_ni ix181 (.Y (nx180), .A0 (nx146), .A1 (nx176), .S0 (Address[1])) ;
    mux21_ni ix147 (.Y (nx146), .A0 (Mem_4__0), .A1 (Mem_5__0), .S0 (Address[0])
             ) ;
    dff reg_Mem_4__0 (.Q (Mem_4__0), .QB (\$dummy [20]), .D (nx4415), .CLK (CLK)
        ) ;
    mux21_ni ix4416 (.Y (nx4415), .A0 (Mem_4__0), .A1 (Din[0]), .S0 (nx9093)) ;
    nand02 ix7095 (.Y (nx7094), .A0 (WR), .A1 (nx8763)) ;
    nor03_2x ix117 (.Y (nx116), .A0 (Address[4]), .A1 (nx8971), .A2 (Address[3])
             ) ;
    dff reg_Mem_5__0 (.Q (Mem_5__0), .QB (\$dummy [21]), .D (nx4425), .CLK (CLK)
        ) ;
    mux21_ni ix4426 (.Y (nx4425), .A0 (Mem_5__0), .A1 (Din[0]), .S0 (nx9095)) ;
    mux21_ni ix177 (.Y (nx176), .A0 (Mem_6__0), .A1 (Mem_7__0), .S0 (Address[0])
             ) ;
    dff reg_Mem_6__0 (.Q (Mem_6__0), .QB (\$dummy [22]), .D (nx4435), .CLK (CLK)
        ) ;
    mux21_ni ix4436 (.Y (nx4435), .A0 (Mem_6__0), .A1 (Din[0]), .S0 (nx9097)) ;
    dff reg_Mem_7__0 (.Q (Mem_7__0), .QB (\$dummy [23]), .D (nx4445), .CLK (CLK)
        ) ;
    mux21_ni ix4446 (.Y (nx4445), .A0 (Mem_7__0), .A1 (Din[0]), .S0 (nx9099)) ;
    nor03_2x ix191 (.Y (nx190), .A0 (Address[4]), .A1 (Address[3]), .A2 (
             Address[2])) ;
    mux21_ni ix83 (.Y (nx82), .A0 (nx42), .A1 (nx78), .S0 (Address[1])) ;
    mux21_ni ix43 (.Y (nx42), .A0 (Mem_24__0), .A1 (Mem_25__0), .S0 (Address[0])
             ) ;
    dff reg_Mem_24__0 (.Q (Mem_24__0), .QB (\$dummy [24]), .D (nx4375), .CLK (
        CLK)) ;
    mux21_ni ix4376 (.Y (nx4375), .A0 (Mem_24__0), .A1 (Din[0]), .S0 (nx9085)) ;
    nand04 ix7118 (.Y (nx7117), .A0 (nx8971), .A1 (Address[3]), .A2 (Address[4])
           , .A3 (WR)) ;
    dff reg_Mem_25__0 (.Q (Mem_25__0), .QB (\$dummy [25]), .D (nx4385), .CLK (
        CLK)) ;
    mux21_ni ix4386 (.Y (nx4385), .A0 (Mem_25__0), .A1 (Din[0]), .S0 (nx9087)) ;
    mux21_ni ix79 (.Y (nx78), .A0 (Mem_26__0), .A1 (Mem_27__0), .S0 (Address[0])
             ) ;
    dff reg_Mem_26__0 (.Q (Mem_26__0), .QB (\$dummy [26]), .D (nx4395), .CLK (
        CLK)) ;
    mux21_ni ix4396 (.Y (nx4395), .A0 (Mem_26__0), .A1 (Din[0]), .S0 (nx9089)) ;
    dff reg_Mem_27__0 (.Q (Mem_27__0), .QB (\$dummy [27]), .D (nx4405), .CLK (
        CLK)) ;
    mux21_ni ix4406 (.Y (nx4405), .A0 (Mem_27__0), .A1 (Din[0]), .S0 (nx9091)) ;
    nor03_2x ix105 (.Y (nx104), .A0 (nx8959), .A1 (Address[3]), .A2 (nx8971)) ;
    nand03 ix941 (.Y (Dout[1]), .A0 (nx7135), .A1 (nx7182), .A2 (nx7214)) ;
    aoi222 ix7136 (.Y (nx7135), .A0 (nx932), .A1 (nx8809), .B0 (nx882), .B1 (
           nx8805), .C0 (nx832), .C1 (nx8801)) ;
    mux21_ni ix933 (.Y (nx932), .A0 (nx904), .A1 (nx928), .S0 (Address[1])) ;
    mux21_ni ix905 (.Y (nx904), .A0 (Mem_28__1), .A1 (Mem_29__1), .S0 (
             Address[0])) ;
    dff reg_Mem_28__1 (.Q (Mem_28__1), .QB (\$dummy [28]), .D (nx4895), .CLK (
        CLK)) ;
    mux21_ni ix4896 (.Y (nx4895), .A0 (Din[1]), .A1 (Mem_28__1), .S0 (nx8939)) ;
    dff reg_Mem_29__1 (.Q (Mem_29__1), .QB (\$dummy [29]), .D (nx4905), .CLK (
        CLK)) ;
    mux21_ni ix4906 (.Y (nx4905), .A0 (Din[1]), .A1 (Mem_29__1), .S0 (nx8943)) ;
    mux21_ni ix929 (.Y (nx928), .A0 (Mem_30__1), .A1 (Mem_31__1), .S0 (
             Address[0])) ;
    dff reg_Mem_30__1 (.Q (Mem_30__1), .QB (\$dummy [30]), .D (nx4915), .CLK (
        CLK)) ;
    mux21_ni ix4916 (.Y (nx4915), .A0 (Din[1]), .A1 (Mem_30__1), .S0 (nx8947)) ;
    dff reg_Mem_31__1 (.Q (Mem_31__1), .QB (\$dummy [31]), .D (nx4925), .CLK (
        CLK)) ;
    mux21_ni ix4926 (.Y (nx4925), .A0 (Din[1]), .A1 (Mem_31__1), .S0 (nx8955)) ;
    mux21_ni ix883 (.Y (nx882), .A0 (nx854), .A1 (nx878), .S0 (Address[1])) ;
    mux21_ni ix855 (.Y (nx854), .A0 (Mem_20__1), .A1 (Mem_21__1), .S0 (
             Address[0])) ;
    dff reg_Mem_20__1 (.Q (Mem_20__1), .QB (\$dummy [32]), .D (nx4855), .CLK (
        CLK)) ;
    mux21_ni ix4856 (.Y (nx4855), .A0 (Din[1]), .A1 (Mem_20__1), .S0 (nx8967)) ;
    dff reg_Mem_21__1 (.Q (Mem_21__1), .QB (\$dummy [33]), .D (nx4865), .CLK (
        CLK)) ;
    mux21_ni ix4866 (.Y (nx4865), .A0 (Din[1]), .A1 (Mem_21__1), .S0 (nx8977)) ;
    mux21_ni ix879 (.Y (nx878), .A0 (Mem_22__1), .A1 (Mem_23__1), .S0 (
             Address[0])) ;
    dff reg_Mem_22__1 (.Q (Mem_22__1), .QB (\$dummy [34]), .D (nx4875), .CLK (
        CLK)) ;
    mux21_ni ix4876 (.Y (nx4875), .A0 (Din[1]), .A1 (Mem_22__1), .S0 (nx8981)) ;
    dff reg_Mem_23__1 (.Q (Mem_23__1), .QB (\$dummy [35]), .D (nx4885), .CLK (
        CLK)) ;
    mux21_ni ix4886 (.Y (nx4885), .A0 (Din[1]), .A1 (Mem_23__1), .S0 (nx8985)) ;
    mux21_ni ix833 (.Y (nx832), .A0 (nx804), .A1 (nx828), .S0 (Address[1])) ;
    mux21_ni ix805 (.Y (nx804), .A0 (Mem_8__1), .A1 (Mem_9__1), .S0 (Address[0])
             ) ;
    dff reg_Mem_8__1 (.Q (Mem_8__1), .QB (\$dummy [36]), .D (nx4815), .CLK (CLK)
        ) ;
    mux21_ni ix4816 (.Y (nx4815), .A0 (Mem_8__1), .A1 (Din[1]), .S0 (nx9115)) ;
    dff reg_Mem_9__1 (.Q (Mem_9__1), .QB (\$dummy [37]), .D (nx4825), .CLK (CLK)
        ) ;
    mux21_ni ix4826 (.Y (nx4825), .A0 (Mem_9__1), .A1 (Din[1]), .S0 (nx9117)) ;
    mux21_ni ix829 (.Y (nx828), .A0 (Mem_10__1), .A1 (Mem_11__1), .S0 (
             Address[0])) ;
    dff reg_Mem_10__1 (.Q (Mem_10__1), .QB (\$dummy [38]), .D (nx4835), .CLK (
        CLK)) ;
    mux21_ni ix4836 (.Y (nx4835), .A0 (Mem_10__1), .A1 (Din[1]), .S0 (nx9119)) ;
    dff reg_Mem_11__1 (.Q (Mem_11__1), .QB (\$dummy [39]), .D (nx4845), .CLK (
        CLK)) ;
    mux21_ni ix4846 (.Y (nx4845), .A0 (Mem_11__1), .A1 (Din[1]), .S0 (nx9121)) ;
    aoi22 ix7183 (.Y (nx7182), .A0 (nx778), .A1 (nx340), .B0 (nx728), .B1 (nx266
          )) ;
    mux21_ni ix779 (.Y (nx778), .A0 (nx750), .A1 (nx774), .S0 (Address[1])) ;
    mux21_ni ix751 (.Y (nx750), .A0 (Mem_12__1), .A1 (Mem_13__1), .S0 (
             Address[0])) ;
    dff reg_Mem_12__1 (.Q (Mem_12__1), .QB (\$dummy [40]), .D (nx4775), .CLK (
        CLK)) ;
    mux21_ni ix4776 (.Y (nx4775), .A0 (Mem_12__1), .A1 (Din[1]), .S0 (nx9109)) ;
    dff reg_Mem_13__1 (.Q (Mem_13__1), .QB (\$dummy [41]), .D (nx4785), .CLK (
        CLK)) ;
    mux21_ni ix4786 (.Y (nx4785), .A0 (Din[1]), .A1 (Mem_13__1), .S0 (nx8997)) ;
    mux21_ni ix775 (.Y (nx774), .A0 (Mem_14__1), .A1 (Mem_15__1), .S0 (
             Address[0])) ;
    dff reg_Mem_14__1 (.Q (Mem_14__1), .QB (\$dummy [42]), .D (nx4795), .CLK (
        CLK)) ;
    mux21_ni ix4796 (.Y (nx4795), .A0 (Mem_14__1), .A1 (Din[1]), .S0 (nx9111)) ;
    dff reg_Mem_15__1 (.Q (Mem_15__1), .QB (\$dummy [43]), .D (nx4805), .CLK (
        CLK)) ;
    mux21_ni ix4806 (.Y (nx4805), .A0 (Mem_15__1), .A1 (Din[1]), .S0 (nx9113)) ;
    mux21_ni ix729 (.Y (nx728), .A0 (nx700), .A1 (nx724), .S0 (Address[1])) ;
    mux21_ni ix701 (.Y (nx700), .A0 (Mem_16__1), .A1 (Mem_17__1), .S0 (
             Address[0])) ;
    dff reg_Mem_16__1 (.Q (Mem_16__1), .QB (\$dummy [44]), .D (nx4735), .CLK (
        CLK)) ;
    mux21_ni ix4736 (.Y (nx4735), .A0 (Mem_16__1), .A1 (Din[1]), .S0 (nx9101)) ;
    dff reg_Mem_17__1 (.Q (Mem_17__1), .QB (\$dummy [45]), .D (nx4745), .CLK (
        CLK)) ;
    mux21_ni ix4746 (.Y (nx4745), .A0 (Mem_17__1), .A1 (Din[1]), .S0 (nx9103)) ;
    mux21_ni ix725 (.Y (nx724), .A0 (Mem_18__1), .A1 (Mem_19__1), .S0 (
             Address[0])) ;
    dff reg_Mem_18__1 (.Q (Mem_18__1), .QB (\$dummy [46]), .D (nx4755), .CLK (
        CLK)) ;
    mux21_ni ix4756 (.Y (nx4755), .A0 (Mem_18__1), .A1 (Din[1]), .S0 (nx9105)) ;
    dff reg_Mem_19__1 (.Q (Mem_19__1), .QB (\$dummy [47]), .D (nx4765), .CLK (
        CLK)) ;
    mux21_ni ix4766 (.Y (nx4765), .A0 (Mem_19__1), .A1 (Din[1]), .S0 (nx9107)) ;
    aoi22 ix7215 (.Y (nx7214), .A0 (nx676), .A1 (nx190), .B0 (nx626), .B1 (nx104
          )) ;
    mux21_ni ix677 (.Y (nx676), .A0 (nx648), .A1 (nx672), .S0 (Address[1])) ;
    mux21_ni ix649 (.Y (nx648), .A0 (Mem_4__1), .A1 (Mem_5__1), .S0 (Address[0])
             ) ;
    dff reg_Mem_4__1 (.Q (Mem_4__1), .QB (\$dummy [48]), .D (nx4695), .CLK (CLK)
        ) ;
    mux21_ni ix4696 (.Y (nx4695), .A0 (Mem_4__1), .A1 (Din[1]), .S0 (nx9093)) ;
    dff reg_Mem_5__1 (.Q (Mem_5__1), .QB (\$dummy [49]), .D (nx4705), .CLK (CLK)
        ) ;
    mux21_ni ix4706 (.Y (nx4705), .A0 (Mem_5__1), .A1 (Din[1]), .S0 (nx9095)) ;
    mux21_ni ix673 (.Y (nx672), .A0 (Mem_6__1), .A1 (Mem_7__1), .S0 (Address[0])
             ) ;
    dff reg_Mem_6__1 (.Q (Mem_6__1), .QB (\$dummy [50]), .D (nx4715), .CLK (CLK)
        ) ;
    mux21_ni ix4716 (.Y (nx4715), .A0 (Mem_6__1), .A1 (Din[1]), .S0 (nx9097)) ;
    dff reg_Mem_7__1 (.Q (Mem_7__1), .QB (\$dummy [51]), .D (nx4725), .CLK (CLK)
        ) ;
    mux21_ni ix4726 (.Y (nx4725), .A0 (Mem_7__1), .A1 (Din[1]), .S0 (nx9099)) ;
    mux21_ni ix627 (.Y (nx626), .A0 (nx598), .A1 (nx622), .S0 (Address[1])) ;
    mux21_ni ix599 (.Y (nx598), .A0 (Mem_24__1), .A1 (Mem_25__1), .S0 (
             Address[0])) ;
    dff reg_Mem_24__1 (.Q (Mem_24__1), .QB (\$dummy [52]), .D (nx4655), .CLK (
        CLK)) ;
    mux21_ni ix4656 (.Y (nx4655), .A0 (Mem_24__1), .A1 (Din[1]), .S0 (nx9085)) ;
    dff reg_Mem_25__1 (.Q (Mem_25__1), .QB (\$dummy [53]), .D (nx4665), .CLK (
        CLK)) ;
    mux21_ni ix4666 (.Y (nx4665), .A0 (Mem_25__1), .A1 (Din[1]), .S0 (nx9087)) ;
    mux21_ni ix623 (.Y (nx622), .A0 (Mem_26__1), .A1 (Mem_27__1), .S0 (
             Address[0])) ;
    dff reg_Mem_26__1 (.Q (Mem_26__1), .QB (\$dummy [54]), .D (nx4675), .CLK (
        CLK)) ;
    mux21_ni ix4676 (.Y (nx4675), .A0 (Mem_26__1), .A1 (Din[1]), .S0 (nx9089)) ;
    dff reg_Mem_27__1 (.Q (Mem_27__1), .QB (\$dummy [55]), .D (nx4685), .CLK (
        CLK)) ;
    mux21_ni ix4686 (.Y (nx4685), .A0 (Mem_27__1), .A1 (Din[1]), .S0 (nx9091)) ;
    nand03 ix1303 (.Y (Dout[2]), .A0 (nx7247), .A1 (nx7294), .A2 (nx7326)) ;
    aoi222 ix7248 (.Y (nx7247), .A0 (nx1294), .A1 (nx8809), .B0 (nx1244), .B1 (
           nx8805), .C0 (nx1194), .C1 (nx8801)) ;
    mux21_ni ix1295 (.Y (nx1294), .A0 (nx1266), .A1 (nx1290), .S0 (Address[1])
             ) ;
    mux21_ni ix1267 (.Y (nx1266), .A0 (Mem_28__2), .A1 (Mem_29__2), .S0 (
             Address[0])) ;
    dff reg_Mem_28__2 (.Q (Mem_28__2), .QB (\$dummy [56]), .D (nx5175), .CLK (
        CLK)) ;
    mux21_ni ix5176 (.Y (nx5175), .A0 (Din[2]), .A1 (Mem_28__2), .S0 (nx8939)) ;
    dff reg_Mem_29__2 (.Q (Mem_29__2), .QB (\$dummy [57]), .D (nx5185), .CLK (
        CLK)) ;
    mux21_ni ix5186 (.Y (nx5185), .A0 (Din[2]), .A1 (Mem_29__2), .S0 (nx8943)) ;
    mux21_ni ix1291 (.Y (nx1290), .A0 (Mem_30__2), .A1 (Mem_31__2), .S0 (
             Address[0])) ;
    dff reg_Mem_30__2 (.Q (Mem_30__2), .QB (\$dummy [58]), .D (nx5195), .CLK (
        CLK)) ;
    mux21_ni ix5196 (.Y (nx5195), .A0 (Din[2]), .A1 (Mem_30__2), .S0 (nx8947)) ;
    dff reg_Mem_31__2 (.Q (Mem_31__2), .QB (\$dummy [59]), .D (nx5205), .CLK (
        CLK)) ;
    mux21_ni ix5206 (.Y (nx5205), .A0 (Din[2]), .A1 (Mem_31__2), .S0 (nx8955)) ;
    mux21_ni ix1245 (.Y (nx1244), .A0 (nx1216), .A1 (nx1240), .S0 (Address[1])
             ) ;
    mux21_ni ix1217 (.Y (nx1216), .A0 (Mem_20__2), .A1 (Mem_21__2), .S0 (
             Address[0])) ;
    dff reg_Mem_20__2 (.Q (Mem_20__2), .QB (\$dummy [60]), .D (nx5135), .CLK (
        CLK)) ;
    mux21_ni ix5136 (.Y (nx5135), .A0 (Din[2]), .A1 (Mem_20__2), .S0 (nx8967)) ;
    dff reg_Mem_21__2 (.Q (Mem_21__2), .QB (\$dummy [61]), .D (nx5145), .CLK (
        CLK)) ;
    mux21_ni ix5146 (.Y (nx5145), .A0 (Din[2]), .A1 (Mem_21__2), .S0 (nx8977)) ;
    mux21_ni ix1241 (.Y (nx1240), .A0 (Mem_22__2), .A1 (Mem_23__2), .S0 (
             Address[0])) ;
    dff reg_Mem_22__2 (.Q (Mem_22__2), .QB (\$dummy [62]), .D (nx5155), .CLK (
        CLK)) ;
    mux21_ni ix5156 (.Y (nx5155), .A0 (Din[2]), .A1 (Mem_22__2), .S0 (nx8981)) ;
    dff reg_Mem_23__2 (.Q (Mem_23__2), .QB (\$dummy [63]), .D (nx5165), .CLK (
        CLK)) ;
    mux21_ni ix5166 (.Y (nx5165), .A0 (Din[2]), .A1 (Mem_23__2), .S0 (nx8985)) ;
    mux21_ni ix1195 (.Y (nx1194), .A0 (nx1166), .A1 (nx1190), .S0 (Address[1])
             ) ;
    mux21_ni ix1167 (.Y (nx1166), .A0 (Mem_8__2), .A1 (Mem_9__2), .S0 (
             Address[0])) ;
    dff reg_Mem_8__2 (.Q (Mem_8__2), .QB (\$dummy [64]), .D (nx5095), .CLK (CLK)
        ) ;
    mux21_ni ix5096 (.Y (nx5095), .A0 (Mem_8__2), .A1 (Din[2]), .S0 (nx9115)) ;
    dff reg_Mem_9__2 (.Q (Mem_9__2), .QB (\$dummy [65]), .D (nx5105), .CLK (CLK)
        ) ;
    mux21_ni ix5106 (.Y (nx5105), .A0 (Mem_9__2), .A1 (Din[2]), .S0 (nx9117)) ;
    mux21_ni ix1191 (.Y (nx1190), .A0 (Mem_10__2), .A1 (Mem_11__2), .S0 (
             Address[0])) ;
    dff reg_Mem_10__2 (.Q (Mem_10__2), .QB (\$dummy [66]), .D (nx5115), .CLK (
        CLK)) ;
    mux21_ni ix5116 (.Y (nx5115), .A0 (Mem_10__2), .A1 (Din[2]), .S0 (nx9119)) ;
    dff reg_Mem_11__2 (.Q (Mem_11__2), .QB (\$dummy [67]), .D (nx5125), .CLK (
        CLK)) ;
    mux21_ni ix5126 (.Y (nx5125), .A0 (Mem_11__2), .A1 (Din[2]), .S0 (nx9121)) ;
    aoi22 ix7295 (.Y (nx7294), .A0 (nx1140), .A1 (nx340), .B0 (nx1090), .B1 (
          nx266)) ;
    mux21_ni ix1141 (.Y (nx1140), .A0 (nx1112), .A1 (nx1136), .S0 (Address[1])
             ) ;
    mux21_ni ix1113 (.Y (nx1112), .A0 (Mem_12__2), .A1 (Mem_13__2), .S0 (
             Address[0])) ;
    dff reg_Mem_12__2 (.Q (Mem_12__2), .QB (\$dummy [68]), .D (nx5055), .CLK (
        CLK)) ;
    mux21_ni ix5056 (.Y (nx5055), .A0 (Mem_12__2), .A1 (Din[2]), .S0 (nx9109)) ;
    dff reg_Mem_13__2 (.Q (Mem_13__2), .QB (\$dummy [69]), .D (nx5065), .CLK (
        CLK)) ;
    mux21_ni ix5066 (.Y (nx5065), .A0 (Din[2]), .A1 (Mem_13__2), .S0 (nx8997)) ;
    mux21_ni ix1137 (.Y (nx1136), .A0 (Mem_14__2), .A1 (Mem_15__2), .S0 (
             Address[0])) ;
    dff reg_Mem_14__2 (.Q (Mem_14__2), .QB (\$dummy [70]), .D (nx5075), .CLK (
        CLK)) ;
    mux21_ni ix5076 (.Y (nx5075), .A0 (Mem_14__2), .A1 (Din[2]), .S0 (nx9111)) ;
    dff reg_Mem_15__2 (.Q (Mem_15__2), .QB (\$dummy [71]), .D (nx5085), .CLK (
        CLK)) ;
    mux21_ni ix5086 (.Y (nx5085), .A0 (Mem_15__2), .A1 (Din[2]), .S0 (nx9113)) ;
    mux21_ni ix1091 (.Y (nx1090), .A0 (nx1062), .A1 (nx1086), .S0 (Address[1])
             ) ;
    mux21_ni ix1063 (.Y (nx1062), .A0 (Mem_16__2), .A1 (Mem_17__2), .S0 (
             Address[0])) ;
    dff reg_Mem_16__2 (.Q (Mem_16__2), .QB (\$dummy [72]), .D (nx5015), .CLK (
        CLK)) ;
    mux21_ni ix5016 (.Y (nx5015), .A0 (Mem_16__2), .A1 (Din[2]), .S0 (nx9101)) ;
    dff reg_Mem_17__2 (.Q (Mem_17__2), .QB (\$dummy [73]), .D (nx5025), .CLK (
        CLK)) ;
    mux21_ni ix5026 (.Y (nx5025), .A0 (Mem_17__2), .A1 (Din[2]), .S0 (nx9103)) ;
    mux21_ni ix1087 (.Y (nx1086), .A0 (Mem_18__2), .A1 (Mem_19__2), .S0 (
             Address[0])) ;
    dff reg_Mem_18__2 (.Q (Mem_18__2), .QB (\$dummy [74]), .D (nx5035), .CLK (
        CLK)) ;
    mux21_ni ix5036 (.Y (nx5035), .A0 (Mem_18__2), .A1 (Din[2]), .S0 (nx9105)) ;
    dff reg_Mem_19__2 (.Q (Mem_19__2), .QB (\$dummy [75]), .D (nx5045), .CLK (
        CLK)) ;
    mux21_ni ix5046 (.Y (nx5045), .A0 (Mem_19__2), .A1 (Din[2]), .S0 (nx9107)) ;
    aoi22 ix7327 (.Y (nx7326), .A0 (nx1038), .A1 (nx190), .B0 (nx988), .B1 (
          nx104)) ;
    mux21_ni ix1039 (.Y (nx1038), .A0 (nx1010), .A1 (nx1034), .S0 (Address[1])
             ) ;
    mux21_ni ix1011 (.Y (nx1010), .A0 (Mem_4__2), .A1 (Mem_5__2), .S0 (
             Address[0])) ;
    dff reg_Mem_4__2 (.Q (Mem_4__2), .QB (\$dummy [76]), .D (nx4975), .CLK (CLK)
        ) ;
    mux21_ni ix4976 (.Y (nx4975), .A0 (Mem_4__2), .A1 (Din[2]), .S0 (nx9093)) ;
    dff reg_Mem_5__2 (.Q (Mem_5__2), .QB (\$dummy [77]), .D (nx4985), .CLK (CLK)
        ) ;
    mux21_ni ix4986 (.Y (nx4985), .A0 (Mem_5__2), .A1 (Din[2]), .S0 (nx9095)) ;
    mux21_ni ix1035 (.Y (nx1034), .A0 (Mem_6__2), .A1 (Mem_7__2), .S0 (
             Address[0])) ;
    dff reg_Mem_6__2 (.Q (Mem_6__2), .QB (\$dummy [78]), .D (nx4995), .CLK (CLK)
        ) ;
    mux21_ni ix4996 (.Y (nx4995), .A0 (Mem_6__2), .A1 (Din[2]), .S0 (nx9097)) ;
    dff reg_Mem_7__2 (.Q (Mem_7__2), .QB (\$dummy [79]), .D (nx5005), .CLK (CLK)
        ) ;
    mux21_ni ix5006 (.Y (nx5005), .A0 (Mem_7__2), .A1 (Din[2]), .S0 (nx9099)) ;
    mux21_ni ix989 (.Y (nx988), .A0 (nx960), .A1 (nx984), .S0 (Address[1])) ;
    mux21_ni ix961 (.Y (nx960), .A0 (Mem_24__2), .A1 (Mem_25__2), .S0 (
             Address[0])) ;
    dff reg_Mem_24__2 (.Q (Mem_24__2), .QB (\$dummy [80]), .D (nx4935), .CLK (
        CLK)) ;
    mux21_ni ix4936 (.Y (nx4935), .A0 (Mem_24__2), .A1 (Din[2]), .S0 (nx9085)) ;
    dff reg_Mem_25__2 (.Q (Mem_25__2), .QB (\$dummy [81]), .D (nx4945), .CLK (
        CLK)) ;
    mux21_ni ix4946 (.Y (nx4945), .A0 (Mem_25__2), .A1 (Din[2]), .S0 (nx9087)) ;
    mux21_ni ix985 (.Y (nx984), .A0 (Mem_26__2), .A1 (Mem_27__2), .S0 (
             Address[0])) ;
    dff reg_Mem_26__2 (.Q (Mem_26__2), .QB (\$dummy [82]), .D (nx4955), .CLK (
        CLK)) ;
    mux21_ni ix4956 (.Y (nx4955), .A0 (Mem_26__2), .A1 (Din[2]), .S0 (nx9089)) ;
    dff reg_Mem_27__2 (.Q (Mem_27__2), .QB (\$dummy [83]), .D (nx4965), .CLK (
        CLK)) ;
    mux21_ni ix4966 (.Y (nx4965), .A0 (Mem_27__2), .A1 (Din[2]), .S0 (nx9091)) ;
    nand03 ix1665 (.Y (Dout[3]), .A0 (nx7359), .A1 (nx7406), .A2 (nx7438)) ;
    aoi222 ix7360 (.Y (nx7359), .A0 (nx1656), .A1 (nx8809), .B0 (nx1606), .B1 (
           nx8805), .C0 (nx1556), .C1 (nx8801)) ;
    mux21_ni ix1657 (.Y (nx1656), .A0 (nx1628), .A1 (nx1652), .S0 (Address[1])
             ) ;
    mux21_ni ix1629 (.Y (nx1628), .A0 (Mem_28__3), .A1 (Mem_29__3), .S0 (
             Address[0])) ;
    dff reg_Mem_28__3 (.Q (Mem_28__3), .QB (\$dummy [84]), .D (nx5455), .CLK (
        CLK)) ;
    mux21_ni ix5456 (.Y (nx5455), .A0 (Din[3]), .A1 (Mem_28__3), .S0 (nx8939)) ;
    dff reg_Mem_29__3 (.Q (Mem_29__3), .QB (\$dummy [85]), .D (nx5465), .CLK (
        CLK)) ;
    mux21_ni ix5466 (.Y (nx5465), .A0 (Din[3]), .A1 (Mem_29__3), .S0 (nx8943)) ;
    mux21_ni ix1653 (.Y (nx1652), .A0 (Mem_30__3), .A1 (Mem_31__3), .S0 (
             Address[0])) ;
    dff reg_Mem_30__3 (.Q (Mem_30__3), .QB (\$dummy [86]), .D (nx5475), .CLK (
        CLK)) ;
    mux21_ni ix5476 (.Y (nx5475), .A0 (Din[3]), .A1 (Mem_30__3), .S0 (nx8947)) ;
    dff reg_Mem_31__3 (.Q (Mem_31__3), .QB (\$dummy [87]), .D (nx5485), .CLK (
        CLK)) ;
    mux21_ni ix5486 (.Y (nx5485), .A0 (Din[3]), .A1 (Mem_31__3), .S0 (nx8955)) ;
    mux21_ni ix1607 (.Y (nx1606), .A0 (nx1578), .A1 (nx1602), .S0 (Address[1])
             ) ;
    mux21_ni ix1579 (.Y (nx1578), .A0 (Mem_20__3), .A1 (Mem_21__3), .S0 (
             Address[0])) ;
    dff reg_Mem_20__3 (.Q (Mem_20__3), .QB (\$dummy [88]), .D (nx5415), .CLK (
        CLK)) ;
    mux21_ni ix5416 (.Y (nx5415), .A0 (Din[3]), .A1 (Mem_20__3), .S0 (nx8967)) ;
    dff reg_Mem_21__3 (.Q (Mem_21__3), .QB (\$dummy [89]), .D (nx5425), .CLK (
        CLK)) ;
    mux21_ni ix5426 (.Y (nx5425), .A0 (Din[3]), .A1 (Mem_21__3), .S0 (nx8977)) ;
    mux21_ni ix1603 (.Y (nx1602), .A0 (Mem_22__3), .A1 (Mem_23__3), .S0 (
             Address[0])) ;
    dff reg_Mem_22__3 (.Q (Mem_22__3), .QB (\$dummy [90]), .D (nx5435), .CLK (
        CLK)) ;
    mux21_ni ix5436 (.Y (nx5435), .A0 (Din[3]), .A1 (Mem_22__3), .S0 (nx8981)) ;
    dff reg_Mem_23__3 (.Q (Mem_23__3), .QB (\$dummy [91]), .D (nx5445), .CLK (
        CLK)) ;
    mux21_ni ix5446 (.Y (nx5445), .A0 (Din[3]), .A1 (Mem_23__3), .S0 (nx8985)) ;
    mux21_ni ix1557 (.Y (nx1556), .A0 (nx1528), .A1 (nx1552), .S0 (Address[1])
             ) ;
    mux21_ni ix1529 (.Y (nx1528), .A0 (Mem_8__3), .A1 (Mem_9__3), .S0 (
             Address[0])) ;
    dff reg_Mem_8__3 (.Q (Mem_8__3), .QB (\$dummy [92]), .D (nx5375), .CLK (CLK)
        ) ;
    mux21_ni ix5376 (.Y (nx5375), .A0 (Mem_8__3), .A1 (Din[3]), .S0 (nx9115)) ;
    dff reg_Mem_9__3 (.Q (Mem_9__3), .QB (\$dummy [93]), .D (nx5385), .CLK (CLK)
        ) ;
    mux21_ni ix5386 (.Y (nx5385), .A0 (Mem_9__3), .A1 (Din[3]), .S0 (nx9117)) ;
    mux21_ni ix1553 (.Y (nx1552), .A0 (Mem_10__3), .A1 (Mem_11__3), .S0 (
             Address[0])) ;
    dff reg_Mem_10__3 (.Q (Mem_10__3), .QB (\$dummy [94]), .D (nx5395), .CLK (
        CLK)) ;
    mux21_ni ix5396 (.Y (nx5395), .A0 (Mem_10__3), .A1 (Din[3]), .S0 (nx9119)) ;
    dff reg_Mem_11__3 (.Q (Mem_11__3), .QB (\$dummy [95]), .D (nx5405), .CLK (
        CLK)) ;
    mux21_ni ix5406 (.Y (nx5405), .A0 (Mem_11__3), .A1 (Din[3]), .S0 (nx9121)) ;
    aoi22 ix7407 (.Y (nx7406), .A0 (nx1502), .A1 (nx340), .B0 (nx1452), .B1 (
          nx266)) ;
    mux21_ni ix1503 (.Y (nx1502), .A0 (nx1474), .A1 (nx1498), .S0 (Address[1])
             ) ;
    mux21_ni ix1475 (.Y (nx1474), .A0 (Mem_12__3), .A1 (Mem_13__3), .S0 (
             Address[0])) ;
    dff reg_Mem_12__3 (.Q (Mem_12__3), .QB (\$dummy [96]), .D (nx5335), .CLK (
        CLK)) ;
    mux21_ni ix5336 (.Y (nx5335), .A0 (Mem_12__3), .A1 (Din[3]), .S0 (nx9109)) ;
    dff reg_Mem_13__3 (.Q (Mem_13__3), .QB (\$dummy [97]), .D (nx5345), .CLK (
        CLK)) ;
    mux21_ni ix5346 (.Y (nx5345), .A0 (Din[3]), .A1 (Mem_13__3), .S0 (nx8997)) ;
    mux21_ni ix1499 (.Y (nx1498), .A0 (Mem_14__3), .A1 (Mem_15__3), .S0 (
             Address[0])) ;
    dff reg_Mem_14__3 (.Q (Mem_14__3), .QB (\$dummy [98]), .D (nx5355), .CLK (
        CLK)) ;
    mux21_ni ix5356 (.Y (nx5355), .A0 (Mem_14__3), .A1 (Din[3]), .S0 (nx9111)) ;
    dff reg_Mem_15__3 (.Q (Mem_15__3), .QB (\$dummy [99]), .D (nx5365), .CLK (
        CLK)) ;
    mux21_ni ix5366 (.Y (nx5365), .A0 (Mem_15__3), .A1 (Din[3]), .S0 (nx9113)) ;
    mux21_ni ix1453 (.Y (nx1452), .A0 (nx1424), .A1 (nx1448), .S0 (Address[1])
             ) ;
    mux21_ni ix1425 (.Y (nx1424), .A0 (Mem_16__3), .A1 (Mem_17__3), .S0 (
             Address[0])) ;
    dff reg_Mem_16__3 (.Q (Mem_16__3), .QB (\$dummy [100]), .D (nx5295), .CLK (
        CLK)) ;
    mux21_ni ix5296 (.Y (nx5295), .A0 (Mem_16__3), .A1 (Din[3]), .S0 (nx9101)) ;
    dff reg_Mem_17__3 (.Q (Mem_17__3), .QB (\$dummy [101]), .D (nx5305), .CLK (
        CLK)) ;
    mux21_ni ix5306 (.Y (nx5305), .A0 (Mem_17__3), .A1 (Din[3]), .S0 (nx9103)) ;
    mux21_ni ix1449 (.Y (nx1448), .A0 (Mem_18__3), .A1 (Mem_19__3), .S0 (
             Address[0])) ;
    dff reg_Mem_18__3 (.Q (Mem_18__3), .QB (\$dummy [102]), .D (nx5315), .CLK (
        CLK)) ;
    mux21_ni ix5316 (.Y (nx5315), .A0 (Mem_18__3), .A1 (Din[3]), .S0 (nx9105)) ;
    dff reg_Mem_19__3 (.Q (Mem_19__3), .QB (\$dummy [103]), .D (nx5325), .CLK (
        CLK)) ;
    mux21_ni ix5326 (.Y (nx5325), .A0 (Mem_19__3), .A1 (Din[3]), .S0 (nx9107)) ;
    aoi22 ix7439 (.Y (nx7438), .A0 (nx1400), .A1 (nx190), .B0 (nx1350), .B1 (
          nx104)) ;
    mux21_ni ix1401 (.Y (nx1400), .A0 (nx1372), .A1 (nx1396), .S0 (Address[1])
             ) ;
    mux21_ni ix1373 (.Y (nx1372), .A0 (Mem_4__3), .A1 (Mem_5__3), .S0 (
             Address[0])) ;
    dff reg_Mem_4__3 (.Q (Mem_4__3), .QB (\$dummy [104]), .D (nx5255), .CLK (CLK
        )) ;
    mux21_ni ix5256 (.Y (nx5255), .A0 (Mem_4__3), .A1 (Din[3]), .S0 (nx9093)) ;
    dff reg_Mem_5__3 (.Q (Mem_5__3), .QB (\$dummy [105]), .D (nx5265), .CLK (CLK
        )) ;
    mux21_ni ix5266 (.Y (nx5265), .A0 (Mem_5__3), .A1 (Din[3]), .S0 (nx9095)) ;
    mux21_ni ix1397 (.Y (nx1396), .A0 (Mem_6__3), .A1 (Mem_7__3), .S0 (
             Address[0])) ;
    dff reg_Mem_6__3 (.Q (Mem_6__3), .QB (\$dummy [106]), .D (nx5275), .CLK (CLK
        )) ;
    mux21_ni ix5276 (.Y (nx5275), .A0 (Mem_6__3), .A1 (Din[3]), .S0 (nx9097)) ;
    dff reg_Mem_7__3 (.Q (Mem_7__3), .QB (\$dummy [107]), .D (nx5285), .CLK (CLK
        )) ;
    mux21_ni ix5286 (.Y (nx5285), .A0 (Mem_7__3), .A1 (Din[3]), .S0 (nx9099)) ;
    mux21_ni ix1351 (.Y (nx1350), .A0 (nx1322), .A1 (nx1346), .S0 (Address[1])
             ) ;
    mux21_ni ix1323 (.Y (nx1322), .A0 (Mem_24__3), .A1 (Mem_25__3), .S0 (
             Address[0])) ;
    dff reg_Mem_24__3 (.Q (Mem_24__3), .QB (\$dummy [108]), .D (nx5215), .CLK (
        CLK)) ;
    mux21_ni ix5216 (.Y (nx5215), .A0 (Mem_24__3), .A1 (Din[3]), .S0 (nx9085)) ;
    dff reg_Mem_25__3 (.Q (Mem_25__3), .QB (\$dummy [109]), .D (nx5225), .CLK (
        CLK)) ;
    mux21_ni ix5226 (.Y (nx5225), .A0 (Mem_25__3), .A1 (Din[3]), .S0 (nx9087)) ;
    mux21_ni ix1347 (.Y (nx1346), .A0 (Mem_26__3), .A1 (Mem_27__3), .S0 (
             Address[0])) ;
    dff reg_Mem_26__3 (.Q (Mem_26__3), .QB (\$dummy [110]), .D (nx5235), .CLK (
        CLK)) ;
    mux21_ni ix5236 (.Y (nx5235), .A0 (Mem_26__3), .A1 (Din[3]), .S0 (nx9089)) ;
    dff reg_Mem_27__3 (.Q (Mem_27__3), .QB (\$dummy [111]), .D (nx5245), .CLK (
        CLK)) ;
    mux21_ni ix5246 (.Y (nx5245), .A0 (Mem_27__3), .A1 (Din[3]), .S0 (nx9091)) ;
    nand03 ix2027 (.Y (Dout[4]), .A0 (nx7471), .A1 (nx7518), .A2 (nx7550)) ;
    aoi222 ix7472 (.Y (nx7471), .A0 (nx2018), .A1 (nx8809), .B0 (nx1968), .B1 (
           nx8805), .C0 (nx1918), .C1 (nx8801)) ;
    mux21_ni ix2019 (.Y (nx2018), .A0 (nx1990), .A1 (nx2014), .S0 (Address[1])
             ) ;
    mux21_ni ix1991 (.Y (nx1990), .A0 (Mem_28__4), .A1 (Mem_29__4), .S0 (
             Address[0])) ;
    dff reg_Mem_28__4 (.Q (Mem_28__4), .QB (\$dummy [112]), .D (nx5735), .CLK (
        CLK)) ;
    mux21_ni ix5736 (.Y (nx5735), .A0 (Din[4]), .A1 (Mem_28__4), .S0 (nx8939)) ;
    dff reg_Mem_29__4 (.Q (Mem_29__4), .QB (\$dummy [113]), .D (nx5745), .CLK (
        CLK)) ;
    mux21_ni ix5746 (.Y (nx5745), .A0 (Din[4]), .A1 (Mem_29__4), .S0 (nx8943)) ;
    mux21_ni ix2015 (.Y (nx2014), .A0 (Mem_30__4), .A1 (Mem_31__4), .S0 (
             Address[0])) ;
    dff reg_Mem_30__4 (.Q (Mem_30__4), .QB (\$dummy [114]), .D (nx5755), .CLK (
        CLK)) ;
    mux21_ni ix5756 (.Y (nx5755), .A0 (Din[4]), .A1 (Mem_30__4), .S0 (nx8947)) ;
    dff reg_Mem_31__4 (.Q (Mem_31__4), .QB (\$dummy [115]), .D (nx5765), .CLK (
        CLK)) ;
    mux21_ni ix5766 (.Y (nx5765), .A0 (Din[4]), .A1 (Mem_31__4), .S0 (nx8955)) ;
    mux21_ni ix1969 (.Y (nx1968), .A0 (nx1940), .A1 (nx1964), .S0 (Address[1])
             ) ;
    mux21_ni ix1941 (.Y (nx1940), .A0 (Mem_20__4), .A1 (Mem_21__4), .S0 (
             Address[0])) ;
    dff reg_Mem_20__4 (.Q (Mem_20__4), .QB (\$dummy [116]), .D (nx5695), .CLK (
        CLK)) ;
    mux21_ni ix5696 (.Y (nx5695), .A0 (Din[4]), .A1 (Mem_20__4), .S0 (nx8967)) ;
    dff reg_Mem_21__4 (.Q (Mem_21__4), .QB (\$dummy [117]), .D (nx5705), .CLK (
        CLK)) ;
    mux21_ni ix5706 (.Y (nx5705), .A0 (Din[4]), .A1 (Mem_21__4), .S0 (nx8977)) ;
    mux21_ni ix1965 (.Y (nx1964), .A0 (Mem_22__4), .A1 (Mem_23__4), .S0 (
             Address[0])) ;
    dff reg_Mem_22__4 (.Q (Mem_22__4), .QB (\$dummy [118]), .D (nx5715), .CLK (
        CLK)) ;
    mux21_ni ix5716 (.Y (nx5715), .A0 (Din[4]), .A1 (Mem_22__4), .S0 (nx8981)) ;
    dff reg_Mem_23__4 (.Q (Mem_23__4), .QB (\$dummy [119]), .D (nx5725), .CLK (
        CLK)) ;
    mux21_ni ix5726 (.Y (nx5725), .A0 (Din[4]), .A1 (Mem_23__4), .S0 (nx8985)) ;
    mux21_ni ix1919 (.Y (nx1918), .A0 (nx1890), .A1 (nx1914), .S0 (Address[1])
             ) ;
    mux21_ni ix1891 (.Y (nx1890), .A0 (Mem_8__4), .A1 (Mem_9__4), .S0 (
             Address[0])) ;
    dff reg_Mem_8__4 (.Q (Mem_8__4), .QB (\$dummy [120]), .D (nx5655), .CLK (CLK
        )) ;
    mux21_ni ix5656 (.Y (nx5655), .A0 (Mem_8__4), .A1 (Din[4]), .S0 (nx9115)) ;
    dff reg_Mem_9__4 (.Q (Mem_9__4), .QB (\$dummy [121]), .D (nx5665), .CLK (CLK
        )) ;
    mux21_ni ix5666 (.Y (nx5665), .A0 (Mem_9__4), .A1 (Din[4]), .S0 (nx9117)) ;
    mux21_ni ix1915 (.Y (nx1914), .A0 (Mem_10__4), .A1 (Mem_11__4), .S0 (
             Address[0])) ;
    dff reg_Mem_10__4 (.Q (Mem_10__4), .QB (\$dummy [122]), .D (nx5675), .CLK (
        CLK)) ;
    mux21_ni ix5676 (.Y (nx5675), .A0 (Mem_10__4), .A1 (Din[4]), .S0 (nx9119)) ;
    dff reg_Mem_11__4 (.Q (Mem_11__4), .QB (\$dummy [123]), .D (nx5685), .CLK (
        CLK)) ;
    mux21_ni ix5686 (.Y (nx5685), .A0 (Mem_11__4), .A1 (Din[4]), .S0 (nx9121)) ;
    aoi22 ix7519 (.Y (nx7518), .A0 (nx1864), .A1 (nx340), .B0 (nx1814), .B1 (
          nx266)) ;
    mux21_ni ix1865 (.Y (nx1864), .A0 (nx1836), .A1 (nx1860), .S0 (Address[1])
             ) ;
    mux21_ni ix1837 (.Y (nx1836), .A0 (Mem_12__4), .A1 (Mem_13__4), .S0 (
             Address[0])) ;
    dff reg_Mem_12__4 (.Q (Mem_12__4), .QB (\$dummy [124]), .D (nx5615), .CLK (
        CLK)) ;
    mux21_ni ix5616 (.Y (nx5615), .A0 (Mem_12__4), .A1 (Din[4]), .S0 (nx9109)) ;
    dff reg_Mem_13__4 (.Q (Mem_13__4), .QB (\$dummy [125]), .D (nx5625), .CLK (
        CLK)) ;
    mux21_ni ix5626 (.Y (nx5625), .A0 (Din[4]), .A1 (Mem_13__4), .S0 (nx8997)) ;
    mux21_ni ix1861 (.Y (nx1860), .A0 (Mem_14__4), .A1 (Mem_15__4), .S0 (
             Address[0])) ;
    dff reg_Mem_14__4 (.Q (Mem_14__4), .QB (\$dummy [126]), .D (nx5635), .CLK (
        CLK)) ;
    mux21_ni ix5636 (.Y (nx5635), .A0 (Mem_14__4), .A1 (Din[4]), .S0 (nx9111)) ;
    dff reg_Mem_15__4 (.Q (Mem_15__4), .QB (\$dummy [127]), .D (nx5645), .CLK (
        CLK)) ;
    mux21_ni ix5646 (.Y (nx5645), .A0 (Mem_15__4), .A1 (Din[4]), .S0 (nx9113)) ;
    mux21_ni ix1815 (.Y (nx1814), .A0 (nx1786), .A1 (nx1810), .S0 (Address[1])
             ) ;
    mux21_ni ix1787 (.Y (nx1786), .A0 (Mem_16__4), .A1 (Mem_17__4), .S0 (
             Address[0])) ;
    dff reg_Mem_16__4 (.Q (Mem_16__4), .QB (\$dummy [128]), .D (nx5575), .CLK (
        CLK)) ;
    mux21_ni ix5576 (.Y (nx5575), .A0 (Mem_16__4), .A1 (Din[4]), .S0 (nx9101)) ;
    dff reg_Mem_17__4 (.Q (Mem_17__4), .QB (\$dummy [129]), .D (nx5585), .CLK (
        CLK)) ;
    mux21_ni ix5586 (.Y (nx5585), .A0 (Mem_17__4), .A1 (Din[4]), .S0 (nx9103)) ;
    mux21_ni ix1811 (.Y (nx1810), .A0 (Mem_18__4), .A1 (Mem_19__4), .S0 (
             Address[0])) ;
    dff reg_Mem_18__4 (.Q (Mem_18__4), .QB (\$dummy [130]), .D (nx5595), .CLK (
        CLK)) ;
    mux21_ni ix5596 (.Y (nx5595), .A0 (Mem_18__4), .A1 (Din[4]), .S0 (nx9105)) ;
    dff reg_Mem_19__4 (.Q (Mem_19__4), .QB (\$dummy [131]), .D (nx5605), .CLK (
        CLK)) ;
    mux21_ni ix5606 (.Y (nx5605), .A0 (Mem_19__4), .A1 (Din[4]), .S0 (nx9107)) ;
    aoi22 ix7551 (.Y (nx7550), .A0 (nx1762), .A1 (nx190), .B0 (nx1712), .B1 (
          nx104)) ;
    mux21_ni ix1763 (.Y (nx1762), .A0 (nx1734), .A1 (nx1758), .S0 (Address[1])
             ) ;
    mux21_ni ix1735 (.Y (nx1734), .A0 (Mem_4__4), .A1 (Mem_5__4), .S0 (
             Address[0])) ;
    dff reg_Mem_4__4 (.Q (Mem_4__4), .QB (\$dummy [132]), .D (nx5535), .CLK (CLK
        )) ;
    mux21_ni ix5536 (.Y (nx5535), .A0 (Mem_4__4), .A1 (Din[4]), .S0 (nx9093)) ;
    dff reg_Mem_5__4 (.Q (Mem_5__4), .QB (\$dummy [133]), .D (nx5545), .CLK (CLK
        )) ;
    mux21_ni ix5546 (.Y (nx5545), .A0 (Mem_5__4), .A1 (Din[4]), .S0 (nx9095)) ;
    mux21_ni ix1759 (.Y (nx1758), .A0 (Mem_6__4), .A1 (Mem_7__4), .S0 (
             Address[0])) ;
    dff reg_Mem_6__4 (.Q (Mem_6__4), .QB (\$dummy [134]), .D (nx5555), .CLK (CLK
        )) ;
    mux21_ni ix5556 (.Y (nx5555), .A0 (Mem_6__4), .A1 (Din[4]), .S0 (nx9097)) ;
    dff reg_Mem_7__4 (.Q (Mem_7__4), .QB (\$dummy [135]), .D (nx5565), .CLK (CLK
        )) ;
    mux21_ni ix5566 (.Y (nx5565), .A0 (Mem_7__4), .A1 (Din[4]), .S0 (nx9099)) ;
    mux21_ni ix1713 (.Y (nx1712), .A0 (nx1684), .A1 (nx1708), .S0 (Address[1])
             ) ;
    mux21_ni ix1685 (.Y (nx1684), .A0 (Mem_24__4), .A1 (Mem_25__4), .S0 (
             Address[0])) ;
    dff reg_Mem_24__4 (.Q (Mem_24__4), .QB (\$dummy [136]), .D (nx5495), .CLK (
        CLK)) ;
    mux21_ni ix5496 (.Y (nx5495), .A0 (Mem_24__4), .A1 (Din[4]), .S0 (nx9085)) ;
    dff reg_Mem_25__4 (.Q (Mem_25__4), .QB (\$dummy [137]), .D (nx5505), .CLK (
        CLK)) ;
    mux21_ni ix5506 (.Y (nx5505), .A0 (Mem_25__4), .A1 (Din[4]), .S0 (nx9087)) ;
    mux21_ni ix1709 (.Y (nx1708), .A0 (Mem_26__4), .A1 (Mem_27__4), .S0 (
             Address[0])) ;
    dff reg_Mem_26__4 (.Q (Mem_26__4), .QB (\$dummy [138]), .D (nx5515), .CLK (
        CLK)) ;
    mux21_ni ix5516 (.Y (nx5515), .A0 (Mem_26__4), .A1 (Din[4]), .S0 (nx9089)) ;
    dff reg_Mem_27__4 (.Q (Mem_27__4), .QB (\$dummy [139]), .D (nx5525), .CLK (
        CLK)) ;
    mux21_ni ix5526 (.Y (nx5525), .A0 (Mem_27__4), .A1 (Din[4]), .S0 (nx9091)) ;
    nand03 ix2389 (.Y (Dout[5]), .A0 (nx7583), .A1 (nx7630), .A2 (nx7662)) ;
    aoi222 ix7584 (.Y (nx7583), .A0 (nx2380), .A1 (nx8809), .B0 (nx2330), .B1 (
           nx8805), .C0 (nx2280), .C1 (nx8801)) ;
    mux21_ni ix2381 (.Y (nx2380), .A0 (nx2352), .A1 (nx2376), .S0 (Address[1])
             ) ;
    mux21_ni ix2353 (.Y (nx2352), .A0 (Mem_28__5), .A1 (Mem_29__5), .S0 (
             Address[0])) ;
    dff reg_Mem_28__5 (.Q (Mem_28__5), .QB (\$dummy [140]), .D (nx6015), .CLK (
        CLK)) ;
    mux21_ni ix6016 (.Y (nx6015), .A0 (Din[5]), .A1 (Mem_28__5), .S0 (nx8939)) ;
    dff reg_Mem_29__5 (.Q (Mem_29__5), .QB (\$dummy [141]), .D (nx6025), .CLK (
        CLK)) ;
    mux21_ni ix6026 (.Y (nx6025), .A0 (Din[5]), .A1 (Mem_29__5), .S0 (nx8943)) ;
    mux21_ni ix2377 (.Y (nx2376), .A0 (Mem_30__5), .A1 (Mem_31__5), .S0 (
             Address[0])) ;
    dff reg_Mem_30__5 (.Q (Mem_30__5), .QB (\$dummy [142]), .D (nx6035), .CLK (
        CLK)) ;
    mux21_ni ix6036 (.Y (nx6035), .A0 (Din[5]), .A1 (Mem_30__5), .S0 (nx8947)) ;
    dff reg_Mem_31__5 (.Q (Mem_31__5), .QB (\$dummy [143]), .D (nx6045), .CLK (
        CLK)) ;
    mux21_ni ix6046 (.Y (nx6045), .A0 (Din[5]), .A1 (Mem_31__5), .S0 (nx8955)) ;
    mux21_ni ix2331 (.Y (nx2330), .A0 (nx2302), .A1 (nx2326), .S0 (Address[1])
             ) ;
    mux21_ni ix2303 (.Y (nx2302), .A0 (Mem_20__5), .A1 (Mem_21__5), .S0 (
             Address[0])) ;
    dff reg_Mem_20__5 (.Q (Mem_20__5), .QB (\$dummy [144]), .D (nx5975), .CLK (
        CLK)) ;
    mux21_ni ix5976 (.Y (nx5975), .A0 (Din[5]), .A1 (Mem_20__5), .S0 (nx8967)) ;
    dff reg_Mem_21__5 (.Q (Mem_21__5), .QB (\$dummy [145]), .D (nx5985), .CLK (
        CLK)) ;
    mux21_ni ix5986 (.Y (nx5985), .A0 (Din[5]), .A1 (Mem_21__5), .S0 (nx8977)) ;
    mux21_ni ix2327 (.Y (nx2326), .A0 (Mem_22__5), .A1 (Mem_23__5), .S0 (
             Address[0])) ;
    dff reg_Mem_22__5 (.Q (Mem_22__5), .QB (\$dummy [146]), .D (nx5995), .CLK (
        CLK)) ;
    mux21_ni ix5996 (.Y (nx5995), .A0 (Din[5]), .A1 (Mem_22__5), .S0 (nx8981)) ;
    dff reg_Mem_23__5 (.Q (Mem_23__5), .QB (\$dummy [147]), .D (nx6005), .CLK (
        CLK)) ;
    mux21_ni ix6006 (.Y (nx6005), .A0 (Din[5]), .A1 (Mem_23__5), .S0 (nx8985)) ;
    mux21_ni ix2281 (.Y (nx2280), .A0 (nx2252), .A1 (nx2276), .S0 (Address[1])
             ) ;
    mux21_ni ix2253 (.Y (nx2252), .A0 (Mem_8__5), .A1 (Mem_9__5), .S0 (
             Address[0])) ;
    dff reg_Mem_8__5 (.Q (Mem_8__5), .QB (\$dummy [148]), .D (nx5935), .CLK (CLK
        )) ;
    mux21_ni ix5936 (.Y (nx5935), .A0 (Mem_8__5), .A1 (Din[5]), .S0 (nx9115)) ;
    dff reg_Mem_9__5 (.Q (Mem_9__5), .QB (\$dummy [149]), .D (nx5945), .CLK (CLK
        )) ;
    mux21_ni ix5946 (.Y (nx5945), .A0 (Mem_9__5), .A1 (Din[5]), .S0 (nx9117)) ;
    mux21_ni ix2277 (.Y (nx2276), .A0 (Mem_10__5), .A1 (Mem_11__5), .S0 (
             Address[0])) ;
    dff reg_Mem_10__5 (.Q (Mem_10__5), .QB (\$dummy [150]), .D (nx5955), .CLK (
        CLK)) ;
    mux21_ni ix5956 (.Y (nx5955), .A0 (Mem_10__5), .A1 (Din[5]), .S0 (nx9119)) ;
    dff reg_Mem_11__5 (.Q (Mem_11__5), .QB (\$dummy [151]), .D (nx5965), .CLK (
        CLK)) ;
    mux21_ni ix5966 (.Y (nx5965), .A0 (Mem_11__5), .A1 (Din[5]), .S0 (nx9121)) ;
    aoi22 ix7631 (.Y (nx7630), .A0 (nx2226), .A1 (nx340), .B0 (nx2176), .B1 (
          nx266)) ;
    mux21_ni ix2227 (.Y (nx2226), .A0 (nx2198), .A1 (nx2222), .S0 (Address[1])
             ) ;
    mux21_ni ix2199 (.Y (nx2198), .A0 (Mem_12__5), .A1 (Mem_13__5), .S0 (
             Address[0])) ;
    dff reg_Mem_12__5 (.Q (Mem_12__5), .QB (\$dummy [152]), .D (nx5895), .CLK (
        CLK)) ;
    mux21_ni ix5896 (.Y (nx5895), .A0 (Mem_12__5), .A1 (Din[5]), .S0 (nx9109)) ;
    dff reg_Mem_13__5 (.Q (Mem_13__5), .QB (\$dummy [153]), .D (nx5905), .CLK (
        CLK)) ;
    mux21_ni ix5906 (.Y (nx5905), .A0 (Din[5]), .A1 (Mem_13__5), .S0 (nx8997)) ;
    mux21_ni ix2223 (.Y (nx2222), .A0 (Mem_14__5), .A1 (Mem_15__5), .S0 (
             Address[0])) ;
    dff reg_Mem_14__5 (.Q (Mem_14__5), .QB (\$dummy [154]), .D (nx5915), .CLK (
        CLK)) ;
    mux21_ni ix5916 (.Y (nx5915), .A0 (Mem_14__5), .A1 (Din[5]), .S0 (nx9111)) ;
    dff reg_Mem_15__5 (.Q (Mem_15__5), .QB (\$dummy [155]), .D (nx5925), .CLK (
        CLK)) ;
    mux21_ni ix5926 (.Y (nx5925), .A0 (Mem_15__5), .A1 (Din[5]), .S0 (nx9113)) ;
    mux21_ni ix2177 (.Y (nx2176), .A0 (nx2148), .A1 (nx2172), .S0 (Address[1])
             ) ;
    mux21_ni ix2149 (.Y (nx2148), .A0 (Mem_16__5), .A1 (Mem_17__5), .S0 (
             Address[0])) ;
    dff reg_Mem_16__5 (.Q (Mem_16__5), .QB (\$dummy [156]), .D (nx5855), .CLK (
        CLK)) ;
    mux21_ni ix5856 (.Y (nx5855), .A0 (Mem_16__5), .A1 (Din[5]), .S0 (nx9101)) ;
    dff reg_Mem_17__5 (.Q (Mem_17__5), .QB (\$dummy [157]), .D (nx5865), .CLK (
        CLK)) ;
    mux21_ni ix5866 (.Y (nx5865), .A0 (Mem_17__5), .A1 (Din[5]), .S0 (nx9103)) ;
    mux21_ni ix2173 (.Y (nx2172), .A0 (Mem_18__5), .A1 (Mem_19__5), .S0 (
             Address[0])) ;
    dff reg_Mem_18__5 (.Q (Mem_18__5), .QB (\$dummy [158]), .D (nx5875), .CLK (
        CLK)) ;
    mux21_ni ix5876 (.Y (nx5875), .A0 (Mem_18__5), .A1 (Din[5]), .S0 (nx9105)) ;
    dff reg_Mem_19__5 (.Q (Mem_19__5), .QB (\$dummy [159]), .D (nx5885), .CLK (
        CLK)) ;
    mux21_ni ix5886 (.Y (nx5885), .A0 (Mem_19__5), .A1 (Din[5]), .S0 (nx9107)) ;
    aoi22 ix7663 (.Y (nx7662), .A0 (nx2124), .A1 (nx190), .B0 (nx2074), .B1 (
          nx104)) ;
    mux21_ni ix2125 (.Y (nx2124), .A0 (nx2096), .A1 (nx2120), .S0 (Address[1])
             ) ;
    mux21_ni ix2097 (.Y (nx2096), .A0 (Mem_4__5), .A1 (Mem_5__5), .S0 (
             Address[0])) ;
    dff reg_Mem_4__5 (.Q (Mem_4__5), .QB (\$dummy [160]), .D (nx5815), .CLK (CLK
        )) ;
    mux21_ni ix5816 (.Y (nx5815), .A0 (Mem_4__5), .A1 (Din[5]), .S0 (nx9093)) ;
    dff reg_Mem_5__5 (.Q (Mem_5__5), .QB (\$dummy [161]), .D (nx5825), .CLK (CLK
        )) ;
    mux21_ni ix5826 (.Y (nx5825), .A0 (Mem_5__5), .A1 (Din[5]), .S0 (nx9095)) ;
    mux21_ni ix2121 (.Y (nx2120), .A0 (Mem_6__5), .A1 (Mem_7__5), .S0 (
             Address[0])) ;
    dff reg_Mem_6__5 (.Q (Mem_6__5), .QB (\$dummy [162]), .D (nx5835), .CLK (CLK
        )) ;
    mux21_ni ix5836 (.Y (nx5835), .A0 (Mem_6__5), .A1 (Din[5]), .S0 (nx9097)) ;
    dff reg_Mem_7__5 (.Q (Mem_7__5), .QB (\$dummy [163]), .D (nx5845), .CLK (CLK
        )) ;
    mux21_ni ix5846 (.Y (nx5845), .A0 (Mem_7__5), .A1 (Din[5]), .S0 (nx9099)) ;
    mux21_ni ix2075 (.Y (nx2074), .A0 (nx2046), .A1 (nx2070), .S0 (Address[1])
             ) ;
    mux21_ni ix2047 (.Y (nx2046), .A0 (Mem_24__5), .A1 (Mem_25__5), .S0 (
             Address[0])) ;
    dff reg_Mem_24__5 (.Q (Mem_24__5), .QB (\$dummy [164]), .D (nx5775), .CLK (
        CLK)) ;
    mux21_ni ix5776 (.Y (nx5775), .A0 (Mem_24__5), .A1 (Din[5]), .S0 (nx9085)) ;
    dff reg_Mem_25__5 (.Q (Mem_25__5), .QB (\$dummy [165]), .D (nx5785), .CLK (
        CLK)) ;
    mux21_ni ix5786 (.Y (nx5785), .A0 (Mem_25__5), .A1 (Din[5]), .S0 (nx9087)) ;
    mux21_ni ix2071 (.Y (nx2070), .A0 (Mem_26__5), .A1 (Mem_27__5), .S0 (
             Address[0])) ;
    dff reg_Mem_26__5 (.Q (Mem_26__5), .QB (\$dummy [166]), .D (nx5795), .CLK (
        CLK)) ;
    mux21_ni ix5796 (.Y (nx5795), .A0 (Mem_26__5), .A1 (Din[5]), .S0 (nx9089)) ;
    dff reg_Mem_27__5 (.Q (Mem_27__5), .QB (\$dummy [167]), .D (nx5805), .CLK (
        CLK)) ;
    mux21_ni ix5806 (.Y (nx5805), .A0 (Mem_27__5), .A1 (Din[5]), .S0 (nx9091)) ;
    nand03 ix2751 (.Y (Dout[6]), .A0 (nx7695), .A1 (nx7742), .A2 (nx7774)) ;
    aoi222 ix7696 (.Y (nx7695), .A0 (nx2742), .A1 (nx8809), .B0 (nx2692), .B1 (
           nx8805), .C0 (nx2642), .C1 (nx8801)) ;
    mux21_ni ix2743 (.Y (nx2742), .A0 (nx2714), .A1 (nx2738), .S0 (Address[1])
             ) ;
    mux21_ni ix2715 (.Y (nx2714), .A0 (Mem_28__6), .A1 (Mem_29__6), .S0 (
             Address[0])) ;
    dff reg_Mem_28__6 (.Q (Mem_28__6), .QB (\$dummy [168]), .D (nx6295), .CLK (
        CLK)) ;
    mux21_ni ix6296 (.Y (nx6295), .A0 (Din[6]), .A1 (Mem_28__6), .S0 (nx8939)) ;
    dff reg_Mem_29__6 (.Q (Mem_29__6), .QB (\$dummy [169]), .D (nx6305), .CLK (
        CLK)) ;
    mux21_ni ix6306 (.Y (nx6305), .A0 (Din[6]), .A1 (Mem_29__6), .S0 (nx8943)) ;
    mux21_ni ix2739 (.Y (nx2738), .A0 (Mem_30__6), .A1 (Mem_31__6), .S0 (
             Address[0])) ;
    dff reg_Mem_30__6 (.Q (Mem_30__6), .QB (\$dummy [170]), .D (nx6315), .CLK (
        CLK)) ;
    mux21_ni ix6316 (.Y (nx6315), .A0 (Din[6]), .A1 (Mem_30__6), .S0 (nx8947)) ;
    dff reg_Mem_31__6 (.Q (Mem_31__6), .QB (\$dummy [171]), .D (nx6325), .CLK (
        CLK)) ;
    mux21_ni ix6326 (.Y (nx6325), .A0 (Din[6]), .A1 (Mem_31__6), .S0 (nx8955)) ;
    mux21_ni ix2693 (.Y (nx2692), .A0 (nx2664), .A1 (nx2688), .S0 (Address[1])
             ) ;
    mux21_ni ix2665 (.Y (nx2664), .A0 (Mem_20__6), .A1 (Mem_21__6), .S0 (
             Address[0])) ;
    dff reg_Mem_20__6 (.Q (Mem_20__6), .QB (\$dummy [172]), .D (nx6255), .CLK (
        CLK)) ;
    mux21_ni ix6256 (.Y (nx6255), .A0 (Din[6]), .A1 (Mem_20__6), .S0 (nx8967)) ;
    dff reg_Mem_21__6 (.Q (Mem_21__6), .QB (\$dummy [173]), .D (nx6265), .CLK (
        CLK)) ;
    mux21_ni ix6266 (.Y (nx6265), .A0 (Din[6]), .A1 (Mem_21__6), .S0 (nx8977)) ;
    mux21_ni ix2689 (.Y (nx2688), .A0 (Mem_22__6), .A1 (Mem_23__6), .S0 (
             Address[0])) ;
    dff reg_Mem_22__6 (.Q (Mem_22__6), .QB (\$dummy [174]), .D (nx6275), .CLK (
        CLK)) ;
    mux21_ni ix6276 (.Y (nx6275), .A0 (Din[6]), .A1 (Mem_22__6), .S0 (nx8981)) ;
    dff reg_Mem_23__6 (.Q (Mem_23__6), .QB (\$dummy [175]), .D (nx6285), .CLK (
        CLK)) ;
    mux21_ni ix6286 (.Y (nx6285), .A0 (Din[6]), .A1 (Mem_23__6), .S0 (nx8985)) ;
    mux21_ni ix2643 (.Y (nx2642), .A0 (nx2614), .A1 (nx2638), .S0 (Address[1])
             ) ;
    mux21_ni ix2615 (.Y (nx2614), .A0 (Mem_8__6), .A1 (Mem_9__6), .S0 (
             Address[0])) ;
    dff reg_Mem_8__6 (.Q (Mem_8__6), .QB (\$dummy [176]), .D (nx6215), .CLK (CLK
        )) ;
    mux21_ni ix6216 (.Y (nx6215), .A0 (Mem_8__6), .A1 (Din[6]), .S0 (nx358)) ;
    dff reg_Mem_9__6 (.Q (Mem_9__6), .QB (\$dummy [177]), .D (nx6225), .CLK (CLK
        )) ;
    mux21_ni ix6226 (.Y (nx6225), .A0 (Mem_9__6), .A1 (Din[6]), .S0 (nx372)) ;
    mux21_ni ix2639 (.Y (nx2638), .A0 (Mem_10__6), .A1 (Mem_11__6), .S0 (
             Address[0])) ;
    dff reg_Mem_10__6 (.Q (Mem_10__6), .QB (\$dummy [178]), .D (nx6235), .CLK (
        CLK)) ;
    mux21_ni ix6236 (.Y (nx6235), .A0 (Mem_10__6), .A1 (Din[6]), .S0 (nx390)) ;
    dff reg_Mem_11__6 (.Q (Mem_11__6), .QB (\$dummy [179]), .D (nx6245), .CLK (
        CLK)) ;
    mux21_ni ix6246 (.Y (nx6245), .A0 (Mem_11__6), .A1 (Din[6]), .S0 (nx402)) ;
    aoi22 ix7743 (.Y (nx7742), .A0 (nx2588), .A1 (nx340), .B0 (nx2538), .B1 (
          nx266)) ;
    mux21_ni ix2589 (.Y (nx2588), .A0 (nx2560), .A1 (nx2584), .S0 (Address[1])
             ) ;
    mux21_ni ix2561 (.Y (nx2560), .A0 (Mem_12__6), .A1 (Mem_13__6), .S0 (
             Address[0])) ;
    dff reg_Mem_12__6 (.Q (Mem_12__6), .QB (\$dummy [180]), .D (nx6175), .CLK (
        CLK)) ;
    mux21_ni ix6176 (.Y (nx6175), .A0 (Mem_12__6), .A1 (Din[6]), .S0 (nx274)) ;
    dff reg_Mem_13__6 (.Q (Mem_13__6), .QB (\$dummy [181]), .D (nx6185), .CLK (
        CLK)) ;
    mux21_ni ix6186 (.Y (nx6185), .A0 (Din[6]), .A1 (Mem_13__6), .S0 (nx8997)) ;
    mux21_ni ix2585 (.Y (nx2584), .A0 (Mem_14__6), .A1 (Mem_15__6), .S0 (
             Address[0])) ;
    dff reg_Mem_14__6 (.Q (Mem_14__6), .QB (\$dummy [182]), .D (nx6195), .CLK (
        CLK)) ;
    mux21_ni ix6196 (.Y (nx6195), .A0 (Mem_14__6), .A1 (Din[6]), .S0 (nx306)) ;
    dff reg_Mem_15__6 (.Q (Mem_15__6), .QB (\$dummy [183]), .D (nx6205), .CLK (
        CLK)) ;
    mux21_ni ix6206 (.Y (nx6205), .A0 (Mem_15__6), .A1 (Din[6]), .S0 (nx318)) ;
    mux21_ni ix2539 (.Y (nx2538), .A0 (nx2510), .A1 (nx2534), .S0 (Address[1])
             ) ;
    mux21_ni ix2511 (.Y (nx2510), .A0 (Mem_16__6), .A1 (Mem_17__6), .S0 (
             Address[0])) ;
    dff reg_Mem_16__6 (.Q (Mem_16__6), .QB (\$dummy [184]), .D (nx6135), .CLK (
        CLK)) ;
    mux21_ni ix6136 (.Y (nx6135), .A0 (Mem_16__6), .A1 (Din[6]), .S0 (nx202)) ;
    dff reg_Mem_17__6 (.Q (Mem_17__6), .QB (\$dummy [185]), .D (nx6145), .CLK (
        CLK)) ;
    mux21_ni ix6146 (.Y (nx6145), .A0 (Mem_17__6), .A1 (Din[6]), .S0 (nx216)) ;
    mux21_ni ix2535 (.Y (nx2534), .A0 (Mem_18__6), .A1 (Mem_19__6), .S0 (
             Address[0])) ;
    dff reg_Mem_18__6 (.Q (Mem_18__6), .QB (\$dummy [186]), .D (nx6155), .CLK (
        CLK)) ;
    mux21_ni ix6156 (.Y (nx6155), .A0 (Mem_18__6), .A1 (Din[6]), .S0 (nx234)) ;
    dff reg_Mem_19__6 (.Q (Mem_19__6), .QB (\$dummy [187]), .D (nx6165), .CLK (
        CLK)) ;
    mux21_ni ix6166 (.Y (nx6165), .A0 (Mem_19__6), .A1 (Din[6]), .S0 (nx246)) ;
    aoi22 ix7775 (.Y (nx7774), .A0 (nx2486), .A1 (nx190), .B0 (nx2436), .B1 (
          nx104)) ;
    mux21_ni ix2487 (.Y (nx2486), .A0 (nx2458), .A1 (nx2482), .S0 (Address[1])
             ) ;
    mux21_ni ix2459 (.Y (nx2458), .A0 (Mem_4__6), .A1 (Mem_5__6), .S0 (
             Address[0])) ;
    dff reg_Mem_4__6 (.Q (Mem_4__6), .QB (\$dummy [188]), .D (nx6095), .CLK (CLK
        )) ;
    mux21_ni ix6096 (.Y (nx6095), .A0 (Mem_4__6), .A1 (Din[6]), .S0 (nx122)) ;
    dff reg_Mem_5__6 (.Q (Mem_5__6), .QB (\$dummy [189]), .D (nx6105), .CLK (CLK
        )) ;
    mux21_ni ix6106 (.Y (nx6105), .A0 (Mem_5__6), .A1 (Din[6]), .S0 (nx136)) ;
    mux21_ni ix2483 (.Y (nx2482), .A0 (Mem_6__6), .A1 (Mem_7__6), .S0 (
             Address[0])) ;
    dff reg_Mem_6__6 (.Q (Mem_6__6), .QB (\$dummy [190]), .D (nx6115), .CLK (CLK
        )) ;
    mux21_ni ix6116 (.Y (nx6115), .A0 (Mem_6__6), .A1 (Din[6]), .S0 (nx154)) ;
    dff reg_Mem_7__6 (.Q (Mem_7__6), .QB (\$dummy [191]), .D (nx6125), .CLK (CLK
        )) ;
    mux21_ni ix6126 (.Y (nx6125), .A0 (Mem_7__6), .A1 (Din[6]), .S0 (nx166)) ;
    mux21_ni ix2437 (.Y (nx2436), .A0 (nx2408), .A1 (nx2432), .S0 (Address[1])
             ) ;
    mux21_ni ix2409 (.Y (nx2408), .A0 (Mem_24__6), .A1 (Mem_25__6), .S0 (
             Address[0])) ;
    dff reg_Mem_24__6 (.Q (Mem_24__6), .QB (\$dummy [192]), .D (nx6055), .CLK (
        CLK)) ;
    mux21_ni ix6056 (.Y (nx6055), .A0 (Mem_24__6), .A1 (Din[6]), .S0 (nx14)) ;
    dff reg_Mem_25__6 (.Q (Mem_25__6), .QB (\$dummy [193]), .D (nx6065), .CLK (
        CLK)) ;
    mux21_ni ix6066 (.Y (nx6065), .A0 (Mem_25__6), .A1 (Din[6]), .S0 (nx32)) ;
    mux21_ni ix2433 (.Y (nx2432), .A0 (Mem_26__6), .A1 (Mem_27__6), .S0 (
             Address[0])) ;
    dff reg_Mem_26__6 (.Q (Mem_26__6), .QB (\$dummy [194]), .D (nx6075), .CLK (
        CLK)) ;
    mux21_ni ix6076 (.Y (nx6075), .A0 (Mem_26__6), .A1 (Din[6]), .S0 (nx54)) ;
    dff reg_Mem_27__6 (.Q (Mem_27__6), .QB (\$dummy [195]), .D (nx6085), .CLK (
        CLK)) ;
    mux21_ni ix6086 (.Y (nx6085), .A0 (Mem_27__6), .A1 (Din[6]), .S0 (nx68)) ;
    nand03 ix3113 (.Y (Dout[7]), .A0 (nx7807), .A1 (nx7854), .A2 (nx7886)) ;
    aoi222 ix7808 (.Y (nx7807), .A0 (nx3104), .A1 (nx8811), .B0 (nx3054), .B1 (
           nx8807), .C0 (nx3004), .C1 (nx8803)) ;
    mux21_ni ix3105 (.Y (nx3104), .A0 (nx3076), .A1 (nx3100), .S0 (Address[1])
             ) ;
    mux21_ni ix3077 (.Y (nx3076), .A0 (Mem_28__7), .A1 (Mem_29__7), .S0 (
             Address[0])) ;
    dff reg_Mem_28__7 (.Q (Mem_28__7), .QB (\$dummy [196]), .D (nx6575), .CLK (
        CLK)) ;
    mux21_ni ix6576 (.Y (nx6575), .A0 (Din[7]), .A1 (Mem_28__7), .S0 (nx8941)) ;
    dff reg_Mem_29__7 (.Q (Mem_29__7), .QB (\$dummy [197]), .D (nx6585), .CLK (
        CLK)) ;
    mux21_ni ix6586 (.Y (nx6585), .A0 (Din[7]), .A1 (Mem_29__7), .S0 (nx8945)) ;
    mux21_ni ix3101 (.Y (nx3100), .A0 (Mem_30__7), .A1 (Mem_31__7), .S0 (
             Address[0])) ;
    dff reg_Mem_30__7 (.Q (Mem_30__7), .QB (\$dummy [198]), .D (nx6595), .CLK (
        CLK)) ;
    mux21_ni ix6596 (.Y (nx6595), .A0 (Din[7]), .A1 (Mem_30__7), .S0 (nx8949)) ;
    dff reg_Mem_31__7 (.Q (Mem_31__7), .QB (\$dummy [199]), .D (nx6605), .CLK (
        CLK)) ;
    mux21_ni ix6606 (.Y (nx6605), .A0 (Din[7]), .A1 (Mem_31__7), .S0 (nx8957)) ;
    mux21_ni ix3055 (.Y (nx3054), .A0 (nx3026), .A1 (nx3050), .S0 (Address[1])
             ) ;
    mux21_ni ix3027 (.Y (nx3026), .A0 (Mem_20__7), .A1 (Mem_21__7), .S0 (
             Address[0])) ;
    dff reg_Mem_20__7 (.Q (Mem_20__7), .QB (\$dummy [200]), .D (nx6535), .CLK (
        CLK)) ;
    mux21_ni ix6536 (.Y (nx6535), .A0 (Din[7]), .A1 (Mem_20__7), .S0 (nx8969)) ;
    dff reg_Mem_21__7 (.Q (Mem_21__7), .QB (\$dummy [201]), .D (nx6545), .CLK (
        CLK)) ;
    mux21_ni ix6546 (.Y (nx6545), .A0 (Din[7]), .A1 (Mem_21__7), .S0 (nx8979)) ;
    mux21_ni ix3051 (.Y (nx3050), .A0 (Mem_22__7), .A1 (Mem_23__7), .S0 (
             Address[0])) ;
    dff reg_Mem_22__7 (.Q (Mem_22__7), .QB (\$dummy [202]), .D (nx6555), .CLK (
        CLK)) ;
    mux21_ni ix6556 (.Y (nx6555), .A0 (Din[7]), .A1 (Mem_22__7), .S0 (nx8983)) ;
    dff reg_Mem_23__7 (.Q (Mem_23__7), .QB (\$dummy [203]), .D (nx6565), .CLK (
        CLK)) ;
    mux21_ni ix6566 (.Y (nx6565), .A0 (Din[7]), .A1 (Mem_23__7), .S0 (nx8987)) ;
    mux21_ni ix3005 (.Y (nx3004), .A0 (nx2976), .A1 (nx3000), .S0 (Address[1])
             ) ;
    mux21_ni ix2977 (.Y (nx2976), .A0 (Mem_8__7), .A1 (Mem_9__7), .S0 (
             Address[0])) ;
    dff reg_Mem_8__7 (.Q (Mem_8__7), .QB (\$dummy [204]), .D (nx6495), .CLK (CLK
        )) ;
    mux21_ni ix6496 (.Y (nx6495), .A0 (Mem_8__7), .A1 (Din[7]), .S0 (nx358)) ;
    dff reg_Mem_9__7 (.Q (Mem_9__7), .QB (\$dummy [205]), .D (nx6505), .CLK (CLK
        )) ;
    mux21_ni ix6506 (.Y (nx6505), .A0 (Mem_9__7), .A1 (Din[7]), .S0 (nx372)) ;
    mux21_ni ix3001 (.Y (nx3000), .A0 (Mem_10__7), .A1 (Mem_11__7), .S0 (
             Address[0])) ;
    dff reg_Mem_10__7 (.Q (Mem_10__7), .QB (\$dummy [206]), .D (nx6515), .CLK (
        CLK)) ;
    mux21_ni ix6516 (.Y (nx6515), .A0 (Mem_10__7), .A1 (Din[7]), .S0 (nx390)) ;
    dff reg_Mem_11__7 (.Q (Mem_11__7), .QB (\$dummy [207]), .D (nx6525), .CLK (
        CLK)) ;
    mux21_ni ix6526 (.Y (nx6525), .A0 (Mem_11__7), .A1 (Din[7]), .S0 (nx402)) ;
    aoi22 ix7855 (.Y (nx7854), .A0 (nx2950), .A1 (nx340), .B0 (nx2900), .B1 (
          nx266)) ;
    mux21_ni ix2951 (.Y (nx2950), .A0 (nx2922), .A1 (nx2946), .S0 (Address[1])
             ) ;
    mux21_ni ix2923 (.Y (nx2922), .A0 (Mem_12__7), .A1 (Mem_13__7), .S0 (
             Address[0])) ;
    dff reg_Mem_12__7 (.Q (Mem_12__7), .QB (\$dummy [208]), .D (nx6455), .CLK (
        CLK)) ;
    mux21_ni ix6456 (.Y (nx6455), .A0 (Mem_12__7), .A1 (Din[7]), .S0 (nx274)) ;
    dff reg_Mem_13__7 (.Q (Mem_13__7), .QB (\$dummy [209]), .D (nx6465), .CLK (
        CLK)) ;
    mux21_ni ix6466 (.Y (nx6465), .A0 (Din[7]), .A1 (Mem_13__7), .S0 (nx8999)) ;
    mux21_ni ix2947 (.Y (nx2946), .A0 (Mem_14__7), .A1 (Mem_15__7), .S0 (
             Address[0])) ;
    dff reg_Mem_14__7 (.Q (Mem_14__7), .QB (\$dummy [210]), .D (nx6475), .CLK (
        CLK)) ;
    mux21_ni ix6476 (.Y (nx6475), .A0 (Mem_14__7), .A1 (Din[7]), .S0 (nx306)) ;
    dff reg_Mem_15__7 (.Q (Mem_15__7), .QB (\$dummy [211]), .D (nx6485), .CLK (
        CLK)) ;
    mux21_ni ix6486 (.Y (nx6485), .A0 (Mem_15__7), .A1 (Din[7]), .S0 (nx318)) ;
    mux21_ni ix2901 (.Y (nx2900), .A0 (nx2872), .A1 (nx2896), .S0 (Address[1])
             ) ;
    mux21_ni ix2873 (.Y (nx2872), .A0 (Mem_16__7), .A1 (Mem_17__7), .S0 (
             Address[0])) ;
    dff reg_Mem_16__7 (.Q (Mem_16__7), .QB (\$dummy [212]), .D (nx6415), .CLK (
        CLK)) ;
    mux21_ni ix6416 (.Y (nx6415), .A0 (Mem_16__7), .A1 (Din[7]), .S0 (nx202)) ;
    dff reg_Mem_17__7 (.Q (Mem_17__7), .QB (\$dummy [213]), .D (nx6425), .CLK (
        CLK)) ;
    mux21_ni ix6426 (.Y (nx6425), .A0 (Mem_17__7), .A1 (Din[7]), .S0 (nx216)) ;
    mux21_ni ix2897 (.Y (nx2896), .A0 (Mem_18__7), .A1 (Mem_19__7), .S0 (
             Address[0])) ;
    dff reg_Mem_18__7 (.Q (Mem_18__7), .QB (\$dummy [214]), .D (nx6435), .CLK (
        CLK)) ;
    mux21_ni ix6436 (.Y (nx6435), .A0 (Mem_18__7), .A1 (Din[7]), .S0 (nx234)) ;
    dff reg_Mem_19__7 (.Q (Mem_19__7), .QB (\$dummy [215]), .D (nx6445), .CLK (
        CLK)) ;
    mux21_ni ix6446 (.Y (nx6445), .A0 (Mem_19__7), .A1 (Din[7]), .S0 (nx246)) ;
    aoi22 ix7887 (.Y (nx7886), .A0 (nx2848), .A1 (nx190), .B0 (nx2798), .B1 (
          nx104)) ;
    mux21_ni ix2849 (.Y (nx2848), .A0 (nx2820), .A1 (nx2844), .S0 (Address[1])
             ) ;
    mux21_ni ix2821 (.Y (nx2820), .A0 (Mem_4__7), .A1 (Mem_5__7), .S0 (
             Address[0])) ;
    dff reg_Mem_4__7 (.Q (Mem_4__7), .QB (\$dummy [216]), .D (nx6375), .CLK (CLK
        )) ;
    mux21_ni ix6376 (.Y (nx6375), .A0 (Mem_4__7), .A1 (Din[7]), .S0 (nx122)) ;
    dff reg_Mem_5__7 (.Q (Mem_5__7), .QB (\$dummy [217]), .D (nx6385), .CLK (CLK
        )) ;
    mux21_ni ix6386 (.Y (nx6385), .A0 (Mem_5__7), .A1 (Din[7]), .S0 (nx136)) ;
    mux21_ni ix2845 (.Y (nx2844), .A0 (Mem_6__7), .A1 (Mem_7__7), .S0 (
             Address[0])) ;
    dff reg_Mem_6__7 (.Q (Mem_6__7), .QB (\$dummy [218]), .D (nx6395), .CLK (CLK
        )) ;
    mux21_ni ix6396 (.Y (nx6395), .A0 (Mem_6__7), .A1 (Din[7]), .S0 (nx154)) ;
    dff reg_Mem_7__7 (.Q (Mem_7__7), .QB (\$dummy [219]), .D (nx6405), .CLK (CLK
        )) ;
    mux21_ni ix6406 (.Y (nx6405), .A0 (Mem_7__7), .A1 (Din[7]), .S0 (nx166)) ;
    mux21_ni ix2799 (.Y (nx2798), .A0 (nx2770), .A1 (nx2794), .S0 (Address[1])
             ) ;
    mux21_ni ix2771 (.Y (nx2770), .A0 (Mem_24__7), .A1 (Mem_25__7), .S0 (
             Address[0])) ;
    dff reg_Mem_24__7 (.Q (Mem_24__7), .QB (\$dummy [220]), .D (nx6335), .CLK (
        CLK)) ;
    mux21_ni ix6336 (.Y (nx6335), .A0 (Mem_24__7), .A1 (Din[7]), .S0 (nx14)) ;
    dff reg_Mem_25__7 (.Q (Mem_25__7), .QB (\$dummy [221]), .D (nx6345), .CLK (
        CLK)) ;
    mux21_ni ix6346 (.Y (nx6345), .A0 (Mem_25__7), .A1 (Din[7]), .S0 (nx32)) ;
    mux21_ni ix2795 (.Y (nx2794), .A0 (Mem_26__7), .A1 (Mem_27__7), .S0 (
             Address[0])) ;
    dff reg_Mem_26__7 (.Q (Mem_26__7), .QB (\$dummy [222]), .D (nx6355), .CLK (
        CLK)) ;
    mux21_ni ix6356 (.Y (nx6355), .A0 (Mem_26__7), .A1 (Din[7]), .S0 (nx54)) ;
    dff reg_Mem_27__7 (.Q (Mem_27__7), .QB (\$dummy [223]), .D (nx6365), .CLK (
        CLK)) ;
    mux21_ni ix6366 (.Y (nx6365), .A0 (Mem_27__7), .A1 (Din[7]), .S0 (nx68)) ;
    nand04 ix3425 (.Y (Dout[8]), .A0 (nx7919), .A1 (nx7947), .A2 (nx7957), .A3 (
           nx7970)) ;
    aoi222 ix7920 (.Y (nx7919), .A0 (nx3392), .A1 (nx8831), .B0 (nx3406), .B1 (
           nx8835), .C0 (nx3376), .C1 (nx8827)) ;
    mux21_ni ix3393 (.Y (nx3392), .A0 (Mem_25__0), .A1 (Mem_24__0), .S0 (
             Address[0])) ;
    and03 ix3397 (.Y (nx3396), .A0 (nx3188), .A1 (nx9053), .A2 (nx8813)) ;
    xnor2 ix7927 (.Y (nx7926), .A0 (Address[3]), .A1 (nx3122)) ;
    xnor2_2x ix3127 (.Y (nx3126), .A0 (nx7929), .A1 (Address[4])) ;
    nand02 ix7930 (.Y (nx7929), .A0 (Address[3]), .A1 (nx3122)) ;
    mux21_ni ix3407 (.Y (nx3406), .A0 (Mem_5__0), .A1 (Mem_4__0), .S0 (
             Address[0])) ;
    nor03_2x ix3415 (.Y (nx3414), .A0 (nx7934), .A1 (nx3148), .A2 (nx9053)) ;
    mux21_ni ix3377 (.Y (nx3376), .A0 (Mem_9__0), .A1 (Mem_8__0), .S0 (
             Address[0])) ;
    nor03_2x ix3383 (.Y (nx3382), .A0 (nx7939), .A1 (nx9053), .A2 (nx9081)) ;
    aoi22 ix7948 (.Y (nx7947), .A0 (nx3342), .A1 (nx3344), .B0 (nx3354), .B1 (
          nx8823)) ;
    mux21_ni ix3343 (.Y (nx3342), .A0 (Mem_21__0), .A1 (Mem_20__0), .S0 (
             Address[0])) ;
    nor02_2x ix3345 (.Y (nx3344), .A0 (nx7951), .A1 (nx7934)) ;
    nand02 ix7952 (.Y (nx7951), .A0 (nx9013), .A1 (nx9053)) ;
    mux21_ni ix3355 (.Y (nx3354), .A0 (Mem_31__0), .A1 (Mem_30__0), .S0 (
             Address[0])) ;
    aoi22 ix7958 (.Y (nx7957), .A0 (nx3294), .A1 (nx3300), .B0 (Mem_3__0), .B1 (
          nx8819)) ;
    mux21_ni ix3295 (.Y (nx3294), .A0 (Mem_13__0), .A1 (Mem_12__0), .S0 (
             Address[0])) ;
    nor03_2x ix3301 (.Y (nx3300), .A0 (nx7934), .A1 (nx9013), .A2 (nx9053)) ;
    dff reg_Mem_3__0 (.Q (Mem_3__0), .QB (\$dummy [224]), .D (nx6615), .CLK (CLK
        )) ;
    mux21_ni ix6616 (.Y (nx6615), .A0 (Din[0]), .A1 (Mem_3__0), .S0 (nx9015)) ;
    nand03 ix7964 (.Y (nx7963), .A0 (nx3308), .A1 (WR), .A2 (nx9049)) ;
    nor03_2x ix3309 (.Y (nx3308), .A0 (Address[4]), .A1 (Address[2]), .A2 (
             Address[3])) ;
    and04 ix7971 (.Y (nx7970), .A0 (nx7972), .A1 (nx7979), .A2 (nx7985), .A3 (
          nx7991)) ;
    aoi22 ix7973 (.Y (nx7972), .A0 (nx3272), .A1 (nx3278), .B0 (nx3260), .B1 (
          nx3262)) ;
    mux21_ni ix3273 (.Y (nx3272), .A0 (Mem_29__0), .A1 (Mem_28__0), .S0 (
             Address[0])) ;
    nor03_2x ix3279 (.Y (nx3278), .A0 (nx7934), .A1 (nx9013), .A2 (nx7955)) ;
    mux21_ni ix3261 (.Y (nx3260), .A0 (Mem_11__0), .A1 (Mem_10__0), .S0 (
             Address[0])) ;
    and02 ix3263 (.Y (nx3262), .A0 (nx3136), .A1 (nx3188)) ;
    aoi22 ix7980 (.Y (nx7979), .A0 (nx3224), .A1 (nx3232), .B0 (nx3242), .B1 (
          nx3248)) ;
    mux21_ni ix3225 (.Y (nx3224), .A0 (Mem_19__0), .A1 (Mem_18__0), .S0 (
             Address[0])) ;
    nor03_2x ix3233 (.Y (nx3232), .A0 (nx7951), .A1 (nx8817), .A2 (nx8813)) ;
    mux21_ni ix3243 (.Y (nx3242), .A0 (Mem_7__0), .A1 (Mem_6__0), .S0 (
             Address[0])) ;
    aoi22 ix7986 (.Y (nx7985), .A0 (nx3204), .A1 (nx3210), .B0 (nx3184), .B1 (
          nx3194)) ;
    mux21_ni ix3205 (.Y (nx3204), .A0 (Mem_17__0), .A1 (Mem_16__0), .S0 (
             Address[0])) ;
    nor03_2x ix3211 (.Y (nx3210), .A0 (nx7951), .A1 (nx8817), .A2 (nx9081)) ;
    mux21_ni ix3185 (.Y (nx3184), .A0 (Mem_27__0), .A1 (Mem_26__0), .S0 (
             Address[0])) ;
    aoi22 ix7992 (.Y (nx7991), .A0 (nx3120), .A1 (nx3152), .B0 (nx3162), .B1 (
          nx3172)) ;
    mux21_ni ix3121 (.Y (nx3120), .A0 (Mem_15__0), .A1 (Mem_14__0), .S0 (
             Address[0])) ;
    nor03_2x ix3153 (.Y (nx3152), .A0 (nx7968), .A1 (nx9079), .A2 (nx9013)) ;
    mux21_ni ix3163 (.Y (nx3162), .A0 (Mem_23__0), .A1 (Mem_22__0), .S0 (
             Address[0])) ;
    nor03_2x ix3173 (.Y (nx3172), .A0 (nx7951), .A1 (nx9079), .A2 (nx8813)) ;
    nand04 ix3601 (.Y (Dout[9]), .A0 (nx7998), .A1 (nx8003), .A2 (nx8007), .A3 (
           nx8013)) ;
    aoi222 ix7999 (.Y (nx7998), .A0 (nx3580), .A1 (nx8831), .B0 (nx3590), .B1 (
           nx8835), .C0 (nx3570), .C1 (nx8827)) ;
    mux21_ni ix3581 (.Y (nx3580), .A0 (Mem_25__1), .A1 (Mem_24__1), .S0 (
             Address[0])) ;
    mux21_ni ix3591 (.Y (nx3590), .A0 (Mem_5__1), .A1 (Mem_4__1), .S0 (
             Address[0])) ;
    mux21_ni ix3571 (.Y (nx3570), .A0 (Mem_9__1), .A1 (Mem_8__1), .S0 (
             Address[0])) ;
    aoi22 ix8004 (.Y (nx8003), .A0 (nx3546), .A1 (nx3344), .B0 (nx3556), .B1 (
          nx8823)) ;
    mux21_ni ix3547 (.Y (nx3546), .A0 (Mem_21__1), .A1 (Mem_20__1), .S0 (
             Address[0])) ;
    mux21_ni ix3557 (.Y (nx3556), .A0 (Mem_31__1), .A1 (Mem_30__1), .S0 (
             Address[0])) ;
    aoi22 ix8008 (.Y (nx8007), .A0 (nx3526), .A1 (nx3300), .B0 (Mem_3__1), .B1 (
          nx8819)) ;
    mux21_ni ix3527 (.Y (nx3526), .A0 (Mem_13__1), .A1 (Mem_12__1), .S0 (
             Address[0])) ;
    dff reg_Mem_3__1 (.Q (Mem_3__1), .QB (\$dummy [225]), .D (nx6625), .CLK (CLK
        )) ;
    mux21_ni ix6626 (.Y (nx6625), .A0 (Din[1]), .A1 (Mem_3__1), .S0 (nx9015)) ;
    and04 ix8014 (.Y (nx8013), .A0 (nx8015), .A1 (nx8019), .A2 (nx8023), .A3 (
          nx8027)) ;
    aoi22 ix8016 (.Y (nx8015), .A0 (nx3510), .A1 (nx3278), .B0 (nx3500), .B1 (
          nx3262)) ;
    mux21_ni ix3511 (.Y (nx3510), .A0 (Mem_29__1), .A1 (Mem_28__1), .S0 (
             Address[0])) ;
    mux21_ni ix3501 (.Y (nx3500), .A0 (Mem_11__1), .A1 (Mem_10__1), .S0 (
             Address[0])) ;
    aoi22 ix8020 (.Y (nx8019), .A0 (nx3478), .A1 (nx3232), .B0 (nx3488), .B1 (
          nx3248)) ;
    mux21_ni ix3479 (.Y (nx3478), .A0 (Mem_19__1), .A1 (Mem_18__1), .S0 (
             Address[0])) ;
    mux21_ni ix3489 (.Y (nx3488), .A0 (Mem_7__1), .A1 (Mem_6__1), .S0 (
             Address[0])) ;
    aoi22 ix8024 (.Y (nx8023), .A0 (nx3464), .A1 (nx3210), .B0 (nx3454), .B1 (
          nx3194)) ;
    mux21_ni ix3465 (.Y (nx3464), .A0 (Mem_17__1), .A1 (Mem_16__1), .S0 (
             Address[0])) ;
    mux21_ni ix3455 (.Y (nx3454), .A0 (Mem_27__1), .A1 (Mem_26__1), .S0 (
             Address[0])) ;
    aoi22 ix8028 (.Y (nx8027), .A0 (nx3432), .A1 (nx3152), .B0 (nx3442), .B1 (
          nx3172)) ;
    mux21_ni ix3433 (.Y (nx3432), .A0 (Mem_15__1), .A1 (Mem_14__1), .S0 (
             Address[0])) ;
    mux21_ni ix3443 (.Y (nx3442), .A0 (Mem_23__1), .A1 (Mem_22__1), .S0 (
             Address[0])) ;
    nand04 ix3777 (.Y (Dout[10]), .A0 (nx8032), .A1 (nx8037), .A2 (nx8041), .A3 (
           nx8047)) ;
    aoi222 ix8033 (.Y (nx8032), .A0 (nx3756), .A1 (nx8831), .B0 (nx3766), .B1 (
           nx8835), .C0 (nx3746), .C1 (nx8827)) ;
    mux21_ni ix3757 (.Y (nx3756), .A0 (Mem_25__2), .A1 (Mem_24__2), .S0 (
             Address[0])) ;
    mux21_ni ix3767 (.Y (nx3766), .A0 (Mem_5__2), .A1 (Mem_4__2), .S0 (
             Address[0])) ;
    mux21_ni ix3747 (.Y (nx3746), .A0 (Mem_9__2), .A1 (Mem_8__2), .S0 (
             Address[0])) ;
    aoi22 ix8038 (.Y (nx8037), .A0 (nx3722), .A1 (nx3344), .B0 (nx3732), .B1 (
          nx8823)) ;
    mux21_ni ix3723 (.Y (nx3722), .A0 (Mem_21__2), .A1 (Mem_20__2), .S0 (
             Address[0])) ;
    mux21_ni ix3733 (.Y (nx3732), .A0 (Mem_31__2), .A1 (Mem_30__2), .S0 (
             Address[0])) ;
    aoi22 ix8042 (.Y (nx8041), .A0 (nx3702), .A1 (nx3300), .B0 (Mem_3__2), .B1 (
          nx8819)) ;
    mux21_ni ix3703 (.Y (nx3702), .A0 (Mem_13__2), .A1 (Mem_12__2), .S0 (
             Address[0])) ;
    dff reg_Mem_3__2 (.Q (Mem_3__2), .QB (\$dummy [226]), .D (nx6635), .CLK (CLK
        )) ;
    mux21_ni ix6636 (.Y (nx6635), .A0 (Din[2]), .A1 (Mem_3__2), .S0 (nx9015)) ;
    and04 ix8048 (.Y (nx8047), .A0 (nx8049), .A1 (nx8053), .A2 (nx8057), .A3 (
          nx8061)) ;
    aoi22 ix8050 (.Y (nx8049), .A0 (nx3686), .A1 (nx3278), .B0 (nx3676), .B1 (
          nx3262)) ;
    mux21_ni ix3687 (.Y (nx3686), .A0 (Mem_29__2), .A1 (Mem_28__2), .S0 (
             Address[0])) ;
    mux21_ni ix3677 (.Y (nx3676), .A0 (Mem_11__2), .A1 (Mem_10__2), .S0 (
             Address[0])) ;
    aoi22 ix8054 (.Y (nx8053), .A0 (nx3654), .A1 (nx3232), .B0 (nx3664), .B1 (
          nx3248)) ;
    mux21_ni ix3655 (.Y (nx3654), .A0 (Mem_19__2), .A1 (Mem_18__2), .S0 (
             Address[0])) ;
    mux21_ni ix3665 (.Y (nx3664), .A0 (Mem_7__2), .A1 (Mem_6__2), .S0 (
             Address[0])) ;
    aoi22 ix8058 (.Y (nx8057), .A0 (nx3640), .A1 (nx3210), .B0 (nx3630), .B1 (
          nx3194)) ;
    mux21_ni ix3641 (.Y (nx3640), .A0 (Mem_17__2), .A1 (Mem_16__2), .S0 (
             Address[0])) ;
    mux21_ni ix3631 (.Y (nx3630), .A0 (Mem_27__2), .A1 (Mem_26__2), .S0 (
             Address[0])) ;
    aoi22 ix8062 (.Y (nx8061), .A0 (nx3608), .A1 (nx3152), .B0 (nx3618), .B1 (
          nx3172)) ;
    mux21_ni ix3609 (.Y (nx3608), .A0 (Mem_15__2), .A1 (Mem_14__2), .S0 (
             Address[0])) ;
    mux21_ni ix3619 (.Y (nx3618), .A0 (Mem_23__2), .A1 (Mem_22__2), .S0 (
             Address[0])) ;
    nand04 ix3953 (.Y (Dout[11]), .A0 (nx8066), .A1 (nx8071), .A2 (nx8075), .A3 (
           nx8081)) ;
    aoi222 ix8067 (.Y (nx8066), .A0 (nx3932), .A1 (nx8831), .B0 (nx3942), .B1 (
           nx8835), .C0 (nx3922), .C1 (nx8827)) ;
    mux21_ni ix3933 (.Y (nx3932), .A0 (Mem_25__3), .A1 (Mem_24__3), .S0 (
             Address[0])) ;
    mux21_ni ix3943 (.Y (nx3942), .A0 (Mem_5__3), .A1 (Mem_4__3), .S0 (
             Address[0])) ;
    mux21_ni ix3923 (.Y (nx3922), .A0 (Mem_9__3), .A1 (Mem_8__3), .S0 (
             Address[0])) ;
    aoi22 ix8072 (.Y (nx8071), .A0 (nx3898), .A1 (nx3344), .B0 (nx3908), .B1 (
          nx8823)) ;
    mux21_ni ix3899 (.Y (nx3898), .A0 (Mem_21__3), .A1 (Mem_20__3), .S0 (
             Address[0])) ;
    mux21_ni ix3909 (.Y (nx3908), .A0 (Mem_31__3), .A1 (Mem_30__3), .S0 (
             Address[0])) ;
    aoi22 ix8076 (.Y (nx8075), .A0 (nx3878), .A1 (nx3300), .B0 (Mem_3__3), .B1 (
          nx8819)) ;
    mux21_ni ix3879 (.Y (nx3878), .A0 (Mem_13__3), .A1 (Mem_12__3), .S0 (
             Address[0])) ;
    dff reg_Mem_3__3 (.Q (Mem_3__3), .QB (\$dummy [227]), .D (nx6645), .CLK (CLK
        )) ;
    mux21_ni ix6646 (.Y (nx6645), .A0 (Din[3]), .A1 (Mem_3__3), .S0 (nx9015)) ;
    and04 ix8082 (.Y (nx8081), .A0 (nx8083), .A1 (nx8087), .A2 (nx8091), .A3 (
          nx8095)) ;
    aoi22 ix8084 (.Y (nx8083), .A0 (nx3862), .A1 (nx3278), .B0 (nx3852), .B1 (
          nx3262)) ;
    mux21_ni ix3863 (.Y (nx3862), .A0 (Mem_29__3), .A1 (Mem_28__3), .S0 (
             Address[0])) ;
    mux21_ni ix3853 (.Y (nx3852), .A0 (Mem_11__3), .A1 (Mem_10__3), .S0 (
             Address[0])) ;
    aoi22 ix8088 (.Y (nx8087), .A0 (nx3830), .A1 (nx3232), .B0 (nx3840), .B1 (
          nx3248)) ;
    mux21_ni ix3831 (.Y (nx3830), .A0 (Mem_19__3), .A1 (Mem_18__3), .S0 (
             Address[0])) ;
    mux21_ni ix3841 (.Y (nx3840), .A0 (Mem_7__3), .A1 (Mem_6__3), .S0 (
             Address[0])) ;
    aoi22 ix8092 (.Y (nx8091), .A0 (nx3816), .A1 (nx3210), .B0 (nx3806), .B1 (
          nx3194)) ;
    mux21_ni ix3817 (.Y (nx3816), .A0 (Mem_17__3), .A1 (Mem_16__3), .S0 (
             Address[0])) ;
    mux21_ni ix3807 (.Y (nx3806), .A0 (Mem_27__3), .A1 (Mem_26__3), .S0 (
             Address[0])) ;
    aoi22 ix8096 (.Y (nx8095), .A0 (nx3784), .A1 (nx3152), .B0 (nx3794), .B1 (
          nx3172)) ;
    mux21_ni ix3785 (.Y (nx3784), .A0 (Mem_15__3), .A1 (Mem_14__3), .S0 (
             Address[0])) ;
    mux21_ni ix3795 (.Y (nx3794), .A0 (Mem_23__3), .A1 (Mem_22__3), .S0 (
             Address[0])) ;
    nand04 ix4129 (.Y (Dout[12]), .A0 (nx8100), .A1 (nx8105), .A2 (nx8109), .A3 (
           nx8115)) ;
    aoi222 ix8101 (.Y (nx8100), .A0 (nx4108), .A1 (nx8831), .B0 (nx4118), .B1 (
           nx8835), .C0 (nx4098), .C1 (nx8827)) ;
    mux21_ni ix4109 (.Y (nx4108), .A0 (Mem_25__4), .A1 (Mem_24__4), .S0 (
             Address[0])) ;
    mux21_ni ix4119 (.Y (nx4118), .A0 (Mem_5__4), .A1 (Mem_4__4), .S0 (
             Address[0])) ;
    mux21_ni ix4099 (.Y (nx4098), .A0 (Mem_9__4), .A1 (Mem_8__4), .S0 (
             Address[0])) ;
    aoi22 ix8106 (.Y (nx8105), .A0 (nx4074), .A1 (nx3344), .B0 (nx4084), .B1 (
          nx8823)) ;
    mux21_ni ix4075 (.Y (nx4074), .A0 (Mem_21__4), .A1 (Mem_20__4), .S0 (
             Address[0])) ;
    mux21_ni ix4085 (.Y (nx4084), .A0 (Mem_31__4), .A1 (Mem_30__4), .S0 (
             Address[0])) ;
    aoi22 ix8110 (.Y (nx8109), .A0 (nx4054), .A1 (nx3300), .B0 (Mem_3__4), .B1 (
          nx8819)) ;
    mux21_ni ix4055 (.Y (nx4054), .A0 (Mem_13__4), .A1 (Mem_12__4), .S0 (
             Address[0])) ;
    dff reg_Mem_3__4 (.Q (Mem_3__4), .QB (\$dummy [228]), .D (nx6655), .CLK (CLK
        )) ;
    mux21_ni ix6656 (.Y (nx6655), .A0 (Din[4]), .A1 (Mem_3__4), .S0 (nx9015)) ;
    and04 ix8116 (.Y (nx8115), .A0 (nx8117), .A1 (nx8121), .A2 (nx8125), .A3 (
          nx8129)) ;
    aoi22 ix8118 (.Y (nx8117), .A0 (nx4038), .A1 (nx3278), .B0 (nx4028), .B1 (
          nx3262)) ;
    mux21_ni ix4039 (.Y (nx4038), .A0 (Mem_29__4), .A1 (Mem_28__4), .S0 (
             Address[0])) ;
    mux21_ni ix4029 (.Y (nx4028), .A0 (Mem_11__4), .A1 (Mem_10__4), .S0 (
             Address[0])) ;
    aoi22 ix8122 (.Y (nx8121), .A0 (nx4006), .A1 (nx3232), .B0 (nx4016), .B1 (
          nx3248)) ;
    mux21_ni ix4007 (.Y (nx4006), .A0 (Mem_19__4), .A1 (Mem_18__4), .S0 (
             Address[0])) ;
    mux21_ni ix4017 (.Y (nx4016), .A0 (Mem_7__4), .A1 (Mem_6__4), .S0 (
             Address[0])) ;
    aoi22 ix8126 (.Y (nx8125), .A0 (nx3992), .A1 (nx3210), .B0 (nx3982), .B1 (
          nx3194)) ;
    mux21_ni ix3993 (.Y (nx3992), .A0 (Mem_17__4), .A1 (Mem_16__4), .S0 (
             Address[0])) ;
    mux21_ni ix3983 (.Y (nx3982), .A0 (Mem_27__4), .A1 (Mem_26__4), .S0 (
             Address[0])) ;
    aoi22 ix8130 (.Y (nx8129), .A0 (nx3960), .A1 (nx3152), .B0 (nx3970), .B1 (
          nx3172)) ;
    mux21_ni ix3961 (.Y (nx3960), .A0 (Mem_15__4), .A1 (Mem_14__4), .S0 (
             Address[0])) ;
    mux21_ni ix3971 (.Y (nx3970), .A0 (Mem_23__4), .A1 (Mem_22__4), .S0 (
             Address[0])) ;
    nand04 ix4305 (.Y (Dout[13]), .A0 (nx8134), .A1 (nx8139), .A2 (nx8143), .A3 (
           nx8149)) ;
    aoi222 ix8135 (.Y (nx8134), .A0 (nx4284), .A1 (nx8831), .B0 (nx4294), .B1 (
           nx8835), .C0 (nx4274), .C1 (nx8827)) ;
    mux21_ni ix4285 (.Y (nx4284), .A0 (Mem_25__5), .A1 (Mem_24__5), .S0 (
             Address[0])) ;
    mux21_ni ix4295 (.Y (nx4294), .A0 (Mem_5__5), .A1 (Mem_4__5), .S0 (
             Address[0])) ;
    mux21_ni ix4275 (.Y (nx4274), .A0 (Mem_9__5), .A1 (Mem_8__5), .S0 (
             Address[0])) ;
    aoi22 ix8140 (.Y (nx8139), .A0 (nx4250), .A1 (nx3344), .B0 (nx4260), .B1 (
          nx8823)) ;
    mux21_ni ix4251 (.Y (nx4250), .A0 (Mem_21__5), .A1 (Mem_20__5), .S0 (
             Address[0])) ;
    mux21_ni ix4261 (.Y (nx4260), .A0 (Mem_31__5), .A1 (Mem_30__5), .S0 (
             Address[0])) ;
    aoi22 ix8144 (.Y (nx8143), .A0 (nx4230), .A1 (nx3300), .B0 (Mem_3__5), .B1 (
          nx8819)) ;
    mux21_ni ix4231 (.Y (nx4230), .A0 (Mem_13__5), .A1 (Mem_12__5), .S0 (
             Address[0])) ;
    dff reg_Mem_3__5 (.Q (Mem_3__5), .QB (\$dummy [229]), .D (nx6665), .CLK (CLK
        )) ;
    mux21_ni ix6666 (.Y (nx6665), .A0 (Din[5]), .A1 (Mem_3__5), .S0 (nx9015)) ;
    and04 ix8150 (.Y (nx8149), .A0 (nx8151), .A1 (nx8155), .A2 (nx8159), .A3 (
          nx8163)) ;
    aoi22 ix8152 (.Y (nx8151), .A0 (nx4214), .A1 (nx3278), .B0 (nx4204), .B1 (
          nx3262)) ;
    mux21_ni ix4215 (.Y (nx4214), .A0 (Mem_29__5), .A1 (Mem_28__5), .S0 (
             Address[0])) ;
    mux21_ni ix4205 (.Y (nx4204), .A0 (Mem_11__5), .A1 (Mem_10__5), .S0 (
             Address[0])) ;
    aoi22 ix8156 (.Y (nx8155), .A0 (nx4182), .A1 (nx3232), .B0 (nx4192), .B1 (
          nx3248)) ;
    mux21_ni ix4183 (.Y (nx4182), .A0 (Mem_19__5), .A1 (Mem_18__5), .S0 (
             Address[0])) ;
    mux21_ni ix4193 (.Y (nx4192), .A0 (Mem_7__5), .A1 (Mem_6__5), .S0 (
             Address[0])) ;
    aoi22 ix8160 (.Y (nx8159), .A0 (nx4168), .A1 (nx3210), .B0 (nx4158), .B1 (
          nx3194)) ;
    mux21_ni ix4169 (.Y (nx4168), .A0 (Mem_17__5), .A1 (Mem_16__5), .S0 (
             Address[0])) ;
    mux21_ni ix4159 (.Y (nx4158), .A0 (Mem_27__5), .A1 (Mem_26__5), .S0 (
             Address[0])) ;
    aoi22 ix8164 (.Y (nx8163), .A0 (nx4136), .A1 (nx3152), .B0 (nx4146), .B1 (
          nx3172)) ;
    mux21_ni ix4137 (.Y (nx4136), .A0 (Mem_15__5), .A1 (Mem_14__5), .S0 (
             Address[0])) ;
    mux21_ni ix4147 (.Y (nx4146), .A0 (Mem_23__5), .A1 (Mem_22__5), .S0 (
             Address[0])) ;
    nand04 ix4481 (.Y (Dout[14]), .A0 (nx8168), .A1 (nx8173), .A2 (nx8177), .A3 (
           nx8183)) ;
    aoi222 ix8169 (.Y (nx8168), .A0 (nx4460), .A1 (nx8831), .B0 (nx4470), .B1 (
           nx8835), .C0 (nx4450), .C1 (nx8827)) ;
    mux21_ni ix4461 (.Y (nx4460), .A0 (Mem_25__6), .A1 (Mem_24__6), .S0 (
             Address[0])) ;
    mux21_ni ix4471 (.Y (nx4470), .A0 (Mem_5__6), .A1 (Mem_4__6), .S0 (
             Address[0])) ;
    mux21_ni ix4451 (.Y (nx4450), .A0 (Mem_9__6), .A1 (Mem_8__6), .S0 (
             Address[0])) ;
    aoi22 ix8174 (.Y (nx8173), .A0 (nx4426), .A1 (nx3344), .B0 (nx4436), .B1 (
          nx8823)) ;
    mux21_ni ix4427 (.Y (nx4426), .A0 (Mem_21__6), .A1 (Mem_20__6), .S0 (
             Address[0])) ;
    mux21_ni ix4437 (.Y (nx4436), .A0 (Mem_31__6), .A1 (Mem_30__6), .S0 (
             Address[0])) ;
    aoi22 ix8178 (.Y (nx8177), .A0 (nx4406), .A1 (nx3300), .B0 (Mem_3__6), .B1 (
          nx8819)) ;
    mux21_ni ix4407 (.Y (nx4406), .A0 (Mem_13__6), .A1 (Mem_12__6), .S0 (
             Address[0])) ;
    dff reg_Mem_3__6 (.Q (Mem_3__6), .QB (\$dummy [230]), .D (nx6675), .CLK (CLK
        )) ;
    mux21_ni ix6676 (.Y (nx6675), .A0 (Din[6]), .A1 (Mem_3__6), .S0 (nx9015)) ;
    and04 ix8184 (.Y (nx8183), .A0 (nx8185), .A1 (nx8189), .A2 (nx8193), .A3 (
          nx8197)) ;
    aoi22 ix8186 (.Y (nx8185), .A0 (nx4390), .A1 (nx3278), .B0 (nx4380), .B1 (
          nx3262)) ;
    mux21_ni ix4391 (.Y (nx4390), .A0 (Mem_29__6), .A1 (Mem_28__6), .S0 (
             Address[0])) ;
    mux21_ni ix4381 (.Y (nx4380), .A0 (Mem_11__6), .A1 (Mem_10__6), .S0 (
             Address[0])) ;
    aoi22 ix8190 (.Y (nx8189), .A0 (nx4358), .A1 (nx3232), .B0 (nx4368), .B1 (
          nx3248)) ;
    mux21_ni ix4359 (.Y (nx4358), .A0 (Mem_19__6), .A1 (Mem_18__6), .S0 (
             Address[0])) ;
    mux21_ni ix4369 (.Y (nx4368), .A0 (Mem_7__6), .A1 (Mem_6__6), .S0 (
             Address[0])) ;
    aoi22 ix8194 (.Y (nx8193), .A0 (nx4344), .A1 (nx3210), .B0 (nx4334), .B1 (
          nx3194)) ;
    mux21_ni ix4348 (.Y (nx4344), .A0 (Mem_17__6), .A1 (Mem_16__6), .S0 (
             Address[0])) ;
    mux21_ni ix4335 (.Y (nx4334), .A0 (Mem_27__6), .A1 (Mem_26__6), .S0 (
             Address[0])) ;
    aoi22 ix8198 (.Y (nx8197), .A0 (nx4312), .A1 (nx3152), .B0 (nx4322), .B1 (
          nx3172)) ;
    mux21_ni ix4313 (.Y (nx4312), .A0 (Mem_15__6), .A1 (Mem_14__6), .S0 (
             Address[0])) ;
    mux21_ni ix4323 (.Y (nx4322), .A0 (Mem_23__6), .A1 (Mem_22__6), .S0 (
             Address[0])) ;
    nand04 ix4657 (.Y (Dout[15]), .A0 (nx8202), .A1 (nx8207), .A2 (nx8211), .A3 (
           nx8217)) ;
    aoi222 ix8203 (.Y (nx8202), .A0 (nx4636), .A1 (nx8833), .B0 (nx4646), .B1 (
           nx8837), .C0 (nx4626), .C1 (nx8829)) ;
    mux21_ni ix4637 (.Y (nx4636), .A0 (Mem_25__7), .A1 (Mem_24__7), .S0 (
             Address[0])) ;
    mux21_ni ix4647 (.Y (nx4646), .A0 (Mem_5__7), .A1 (Mem_4__7), .S0 (
             Address[0])) ;
    mux21_ni ix4627 (.Y (nx4626), .A0 (Mem_9__7), .A1 (Mem_8__7), .S0 (
             Address[0])) ;
    aoi22 ix8208 (.Y (nx8207), .A0 (nx4602), .A1 (nx3344), .B0 (nx4612), .B1 (
          nx8825)) ;
    mux21_ni ix4603 (.Y (nx4602), .A0 (Mem_21__7), .A1 (Mem_20__7), .S0 (
             Address[0])) ;
    mux21_ni ix4613 (.Y (nx4612), .A0 (Mem_31__7), .A1 (Mem_30__7), .S0 (
             Address[0])) ;
    aoi22 ix8212 (.Y (nx8211), .A0 (nx4582), .A1 (nx3300), .B0 (Mem_3__7), .B1 (
          nx8821)) ;
    mux21_ni ix4583 (.Y (nx4582), .A0 (Mem_13__7), .A1 (Mem_12__7), .S0 (
             Address[0])) ;
    dff reg_Mem_3__7 (.Q (Mem_3__7), .QB (\$dummy [231]), .D (nx6685), .CLK (CLK
        )) ;
    mux21_ni ix6686 (.Y (nx6685), .A0 (Din[7]), .A1 (Mem_3__7), .S0 (nx9017)) ;
    and04 ix8218 (.Y (nx8217), .A0 (nx8219), .A1 (nx8223), .A2 (nx8227), .A3 (
          nx8231)) ;
    aoi22 ix8220 (.Y (nx8219), .A0 (nx4566), .A1 (nx3278), .B0 (nx4556), .B1 (
          nx3262)) ;
    mux21_ni ix4567 (.Y (nx4566), .A0 (Mem_29__7), .A1 (Mem_28__7), .S0 (
             Address[0])) ;
    mux21_ni ix4557 (.Y (nx4556), .A0 (Mem_11__7), .A1 (Mem_10__7), .S0 (
             Address[0])) ;
    aoi22 ix8224 (.Y (nx8223), .A0 (nx4534), .A1 (nx3232), .B0 (nx4544), .B1 (
          nx3248)) ;
    mux21_ni ix4535 (.Y (nx4534), .A0 (Mem_19__7), .A1 (Mem_18__7), .S0 (
             Address[0])) ;
    mux21_ni ix4545 (.Y (nx4544), .A0 (Mem_7__7), .A1 (Mem_6__7), .S0 (
             Address[0])) ;
    aoi22 ix8228 (.Y (nx8227), .A0 (nx4520), .A1 (nx3210), .B0 (nx4510), .B1 (
          nx3194)) ;
    mux21_ni ix4521 (.Y (nx4520), .A0 (Mem_17__7), .A1 (Mem_16__7), .S0 (
             Address[0])) ;
    mux21_ni ix4511 (.Y (nx4510), .A0 (Mem_27__7), .A1 (Mem_26__7), .S0 (
             Address[0])) ;
    aoi22 ix8232 (.Y (nx8231), .A0 (nx4488), .A1 (nx3152), .B0 (nx4498), .B1 (
          nx3172)) ;
    mux21_ni ix4489 (.Y (nx4488), .A0 (Mem_15__7), .A1 (Mem_14__7), .S0 (
             Address[0])) ;
    mux21_ni ix4499 (.Y (nx4498), .A0 (Mem_23__7), .A1 (Mem_22__7), .S0 (
             Address[0])) ;
    nand04 ix4841 (.Y (Dout[16]), .A0 (nx8236), .A1 (nx8241), .A2 (nx8245), .A3 (
           nx8249)) ;
    aoi222 ix8237 (.Y (nx8236), .A0 (nx256), .A1 (nx8887), .B0 (nx226), .B1 (
           nx8895), .C0 (nx298), .C1 (nx8891)) ;
    nor04 ix4815 (.Y (nx4814), .A0 (Address[3]), .A1 (Address[2]), .A2 (
          Address[1]), .A3 (nx8959)) ;
    nor04 ix4823 (.Y (nx4822), .A0 (nx8951), .A1 (nx8963), .A2 (Address[2]), .A3 (
          Address[4])) ;
    aoi22 ix8242 (.Y (nx8241), .A0 (nx176), .A1 (nx8879), .B0 (nx42), .B1 (
          nx8883)) ;
    nor04 ix4799 (.Y (nx4798), .A0 (Address[1]), .A1 (nx8973), .A2 (Address[3])
          , .A3 (Address[4])) ;
    aoi22 ix8246 (.Y (nx8245), .A0 (nx328), .A1 (nx8871), .B0 (nx382), .B1 (
          nx8875)) ;
    nor04 ix4783 (.Y (nx4782), .A0 (Address[1]), .A1 (nx8973), .A2 (nx8963), .A3 (
          Address[4])) ;
    nor04 ix4793 (.Y (nx4792), .A0 (nx8951), .A1 (Address[3]), .A2 (nx8973), .A3 (
          Address[4])) ;
    and04 ix8250 (.Y (nx8249), .A0 (nx8251), .A1 (nx8255), .A2 (nx8259), .A3 (
          nx8263)) ;
    aoi22 ix8252 (.Y (nx8251), .A0 (nx486), .A1 (nx8867), .B0 (nx560), .B1 (
          nx8863)) ;
    nor04 ix4769 (.Y (nx4768), .A0 (Address[3]), .A1 (nx8973), .A2 (Address[1])
          , .A3 (nx8959)) ;
    aoi22 ix8256 (.Y (nx8255), .A0 (nx456), .A1 (nx8859), .B0 (nx530), .B1 (
          nx8855)) ;
    nor04 ix4753 (.Y (nx4752), .A0 (Address[3]), .A1 (Address[2]), .A2 (nx8951)
          , .A3 (nx8961)) ;
    aoi22 ix8260 (.Y (nx8259), .A0 (nx78), .A1 (nx8851), .B0 (nx146), .B1 (
          nx8847)) ;
    nor04 ix4731 (.Y (nx4730), .A0 (Address[1]), .A1 (Address[2]), .A2 (nx8965)
          , .A3 (nx8961)) ;
    nor04 ix4725 (.Y (nx4724), .A0 (Address[3]), .A1 (Address[2]), .A2 (nx8951)
          , .A3 (Address[4])) ;
    aoi22 ix8264 (.Y (nx8263), .A0 (nx412), .A1 (nx8843), .B0 (nx4676), .B1 (
          nx8839)) ;
    nor04 ix4717 (.Y (nx4716), .A0 (Address[1]), .A1 (Address[2]), .A2 (nx8965)
          , .A3 (Address[4])) ;
    mux21_ni ix4677 (.Y (nx4676), .A0 (Mem_2__0), .A1 (Mem_3__0), .S0 (
             Address[0])) ;
    dff reg_Mem_2__0 (.Q (Mem_2__0), .QB (\$dummy [232]), .D (nx6695), .CLK (CLK
        )) ;
    mux21_ni ix6696 (.Y (nx6695), .A0 (Din[0]), .A1 (Mem_2__0), .S0 (nx9019)) ;
    nand03 ix8270 (.Y (nx8269), .A0 (nx3308), .A1 (WR), .A2 (nx9075)) ;
    nor04 ix4709 (.Y (nx4708), .A0 (Address[1]), .A1 (Address[2]), .A2 (
          Address[3]), .A3 (Address[4])) ;
    nand04 ix4913 (.Y (Dout[17]), .A0 (nx8274), .A1 (nx8276), .A2 (nx8278), .A3 (
           nx8280)) ;
    aoi222 ix8275 (.Y (nx8274), .A0 (nx724), .A1 (nx8887), .B0 (nx700), .B1 (
           nx8895), .C0 (nx750), .C1 (nx8891)) ;
    aoi22 ix8277 (.Y (nx8276), .A0 (nx672), .A1 (nx8879), .B0 (nx598), .B1 (
          nx8883)) ;
    aoi22 ix8279 (.Y (nx8278), .A0 (nx774), .A1 (nx8871), .B0 (nx804), .B1 (
          nx8875)) ;
    and04 ix8281 (.Y (nx8280), .A0 (nx8282), .A1 (nx8284), .A2 (nx8286), .A3 (
          nx8288)) ;
    aoi22 ix8283 (.Y (nx8282), .A0 (nx878), .A1 (nx8867), .B0 (nx928), .B1 (
          nx8863)) ;
    aoi22 ix8285 (.Y (nx8284), .A0 (nx854), .A1 (nx8859), .B0 (nx904), .B1 (
          nx8855)) ;
    aoi22 ix8287 (.Y (nx8286), .A0 (nx622), .A1 (nx8851), .B0 (nx648), .B1 (
          nx8847)) ;
    aoi22 ix8289 (.Y (nx8288), .A0 (nx828), .A1 (nx8843), .B0 (nx4854), .B1 (
          nx8839)) ;
    mux21_ni ix4855 (.Y (nx4854), .A0 (Mem_2__1), .A1 (Mem_3__1), .S0 (
             Address[0])) ;
    dff reg_Mem_2__1 (.Q (Mem_2__1), .QB (\$dummy [233]), .D (nx6705), .CLK (CLK
        )) ;
    mux21_ni ix6706 (.Y (nx6705), .A0 (Din[1]), .A1 (Mem_2__1), .S0 (nx9019)) ;
    nand04 ix4985 (.Y (Dout[18]), .A0 (nx8295), .A1 (nx8297), .A2 (nx8299), .A3 (
           nx8301)) ;
    aoi222 ix8296 (.Y (nx8295), .A0 (nx1086), .A1 (nx8887), .B0 (nx1062), .B1 (
           nx8895), .C0 (nx1112), .C1 (nx8891)) ;
    aoi22 ix8298 (.Y (nx8297), .A0 (nx1034), .A1 (nx8879), .B0 (nx960), .B1 (
          nx8883)) ;
    aoi22 ix8300 (.Y (nx8299), .A0 (nx1136), .A1 (nx8871), .B0 (nx1166), .B1 (
          nx8875)) ;
    and04 ix8302 (.Y (nx8301), .A0 (nx8303), .A1 (nx8305), .A2 (nx8307), .A3 (
          nx8309)) ;
    aoi22 ix8304 (.Y (nx8303), .A0 (nx1240), .A1 (nx8867), .B0 (nx1290), .B1 (
          nx8863)) ;
    aoi22 ix8306 (.Y (nx8305), .A0 (nx1216), .A1 (nx8859), .B0 (nx1266), .B1 (
          nx8855)) ;
    aoi22 ix8308 (.Y (nx8307), .A0 (nx984), .A1 (nx8851), .B0 (nx1010), .B1 (
          nx8847)) ;
    aoi22 ix8310 (.Y (nx8309), .A0 (nx1190), .A1 (nx8843), .B0 (nx4926), .B1 (
          nx8839)) ;
    mux21_ni ix4927 (.Y (nx4926), .A0 (Mem_2__2), .A1 (Mem_3__2), .S0 (
             Address[0])) ;
    dff reg_Mem_2__2 (.Q (Mem_2__2), .QB (\$dummy [234]), .D (nx6715), .CLK (CLK
        )) ;
    mux21_ni ix6716 (.Y (nx6715), .A0 (Din[2]), .A1 (Mem_2__2), .S0 (nx9019)) ;
    nand04 ix5057 (.Y (Dout[19]), .A0 (nx8316), .A1 (nx8318), .A2 (nx8320), .A3 (
           nx8322)) ;
    aoi222 ix8317 (.Y (nx8316), .A0 (nx1448), .A1 (nx8887), .B0 (nx1424), .B1 (
           nx8895), .C0 (nx1474), .C1 (nx8891)) ;
    aoi22 ix8319 (.Y (nx8318), .A0 (nx1396), .A1 (nx8879), .B0 (nx1322), .B1 (
          nx8883)) ;
    aoi22 ix8321 (.Y (nx8320), .A0 (nx1498), .A1 (nx8871), .B0 (nx1528), .B1 (
          nx8875)) ;
    and04 ix8323 (.Y (nx8322), .A0 (nx8324), .A1 (nx8326), .A2 (nx8328), .A3 (
          nx8330)) ;
    aoi22 ix8325 (.Y (nx8324), .A0 (nx1602), .A1 (nx8867), .B0 (nx1652), .B1 (
          nx8863)) ;
    aoi22 ix8327 (.Y (nx8326), .A0 (nx1578), .A1 (nx8859), .B0 (nx1628), .B1 (
          nx8855)) ;
    aoi22 ix8329 (.Y (nx8328), .A0 (nx1346), .A1 (nx8851), .B0 (nx1372), .B1 (
          nx8847)) ;
    aoi22 ix8331 (.Y (nx8330), .A0 (nx1552), .A1 (nx8843), .B0 (nx4998), .B1 (
          nx8839)) ;
    mux21_ni ix4999 (.Y (nx4998), .A0 (Mem_2__3), .A1 (Mem_3__3), .S0 (
             Address[0])) ;
    dff reg_Mem_2__3 (.Q (Mem_2__3), .QB (\$dummy [235]), .D (nx6725), .CLK (CLK
        )) ;
    mux21_ni ix6726 (.Y (nx6725), .A0 (Din[3]), .A1 (Mem_2__3), .S0 (nx9019)) ;
    nand04 ix5129 (.Y (Dout[20]), .A0 (nx8337), .A1 (nx8339), .A2 (nx8341), .A3 (
           nx8343)) ;
    aoi222 ix8338 (.Y (nx8337), .A0 (nx1810), .A1 (nx8887), .B0 (nx1786), .B1 (
           nx8895), .C0 (nx1836), .C1 (nx8891)) ;
    aoi22 ix8340 (.Y (nx8339), .A0 (nx1758), .A1 (nx8879), .B0 (nx1684), .B1 (
          nx8883)) ;
    aoi22 ix8342 (.Y (nx8341), .A0 (nx1860), .A1 (nx8871), .B0 (nx1890), .B1 (
          nx8875)) ;
    and04 ix8344 (.Y (nx8343), .A0 (nx8345), .A1 (nx8347), .A2 (nx8349), .A3 (
          nx8351)) ;
    aoi22 ix8346 (.Y (nx8345), .A0 (nx1964), .A1 (nx8867), .B0 (nx2014), .B1 (
          nx8863)) ;
    aoi22 ix8348 (.Y (nx8347), .A0 (nx1940), .A1 (nx8859), .B0 (nx1990), .B1 (
          nx8855)) ;
    aoi22 ix8350 (.Y (nx8349), .A0 (nx1708), .A1 (nx8851), .B0 (nx1734), .B1 (
          nx8847)) ;
    aoi22 ix8352 (.Y (nx8351), .A0 (nx1914), .A1 (nx8843), .B0 (nx5070), .B1 (
          nx8839)) ;
    mux21_ni ix5071 (.Y (nx5070), .A0 (Mem_2__4), .A1 (Mem_3__4), .S0 (
             Address[0])) ;
    dff reg_Mem_2__4 (.Q (Mem_2__4), .QB (\$dummy [236]), .D (nx6735), .CLK (CLK
        )) ;
    mux21_ni ix6736 (.Y (nx6735), .A0 (Din[4]), .A1 (Mem_2__4), .S0 (nx9019)) ;
    nand04 ix5201 (.Y (Dout[21]), .A0 (nx8358), .A1 (nx8360), .A2 (nx8362), .A3 (
           nx8364)) ;
    aoi222 ix8359 (.Y (nx8358), .A0 (nx2172), .A1 (nx8887), .B0 (nx2148), .B1 (
           nx8895), .C0 (nx2198), .C1 (nx8891)) ;
    aoi22 ix8361 (.Y (nx8360), .A0 (nx2120), .A1 (nx8879), .B0 (nx2046), .B1 (
          nx8883)) ;
    aoi22 ix8363 (.Y (nx8362), .A0 (nx2222), .A1 (nx8871), .B0 (nx2252), .B1 (
          nx8875)) ;
    and04 ix8365 (.Y (nx8364), .A0 (nx8366), .A1 (nx8368), .A2 (nx8370), .A3 (
          nx8372)) ;
    aoi22 ix8367 (.Y (nx8366), .A0 (nx2326), .A1 (nx8867), .B0 (nx2376), .B1 (
          nx8863)) ;
    aoi22 ix8369 (.Y (nx8368), .A0 (nx2302), .A1 (nx8859), .B0 (nx2352), .B1 (
          nx8855)) ;
    aoi22 ix8371 (.Y (nx8370), .A0 (nx2070), .A1 (nx8851), .B0 (nx2096), .B1 (
          nx8847)) ;
    aoi22 ix8373 (.Y (nx8372), .A0 (nx2276), .A1 (nx8843), .B0 (nx5142), .B1 (
          nx8839)) ;
    mux21_ni ix5143 (.Y (nx5142), .A0 (Mem_2__5), .A1 (Mem_3__5), .S0 (
             Address[0])) ;
    dff reg_Mem_2__5 (.Q (Mem_2__5), .QB (\$dummy [237]), .D (nx6745), .CLK (CLK
        )) ;
    mux21_ni ix6746 (.Y (nx6745), .A0 (Din[5]), .A1 (Mem_2__5), .S0 (nx9019)) ;
    nand04 ix5273 (.Y (Dout[22]), .A0 (nx8379), .A1 (nx8381), .A2 (nx8383), .A3 (
           nx8385)) ;
    aoi222 ix8380 (.Y (nx8379), .A0 (nx2534), .A1 (nx8887), .B0 (nx2510), .B1 (
           nx8895), .C0 (nx2560), .C1 (nx8891)) ;
    aoi22 ix8382 (.Y (nx8381), .A0 (nx2482), .A1 (nx8879), .B0 (nx2408), .B1 (
          nx8883)) ;
    aoi22 ix8384 (.Y (nx8383), .A0 (nx2584), .A1 (nx8871), .B0 (nx2614), .B1 (
          nx8875)) ;
    and04 ix8386 (.Y (nx8385), .A0 (nx8387), .A1 (nx8389), .A2 (nx8391), .A3 (
          nx8393)) ;
    aoi22 ix8388 (.Y (nx8387), .A0 (nx2688), .A1 (nx8867), .B0 (nx2738), .B1 (
          nx8863)) ;
    aoi22 ix8390 (.Y (nx8389), .A0 (nx2664), .A1 (nx8859), .B0 (nx2714), .B1 (
          nx8855)) ;
    aoi22 ix8392 (.Y (nx8391), .A0 (nx2432), .A1 (nx8851), .B0 (nx2458), .B1 (
          nx8847)) ;
    aoi22 ix8394 (.Y (nx8393), .A0 (nx2638), .A1 (nx8843), .B0 (nx5214), .B1 (
          nx8839)) ;
    mux21_ni ix5215 (.Y (nx5214), .A0 (Mem_2__6), .A1 (Mem_3__6), .S0 (
             Address[0])) ;
    dff reg_Mem_2__6 (.Q (Mem_2__6), .QB (\$dummy [238]), .D (nx6755), .CLK (CLK
        )) ;
    mux21_ni ix6756 (.Y (nx6755), .A0 (Din[6]), .A1 (Mem_2__6), .S0 (nx9019)) ;
    nand04 ix5345 (.Y (Dout[23]), .A0 (nx8400), .A1 (nx8402), .A2 (nx8404), .A3 (
           nx8406)) ;
    aoi222 ix8401 (.Y (nx8400), .A0 (nx2896), .A1 (nx8889), .B0 (nx2872), .B1 (
           nx8897), .C0 (nx2922), .C1 (nx8893)) ;
    aoi22 ix8403 (.Y (nx8402), .A0 (nx2844), .A1 (nx8881), .B0 (nx2770), .B1 (
          nx8885)) ;
    aoi22 ix8405 (.Y (nx8404), .A0 (nx2946), .A1 (nx8873), .B0 (nx2976), .B1 (
          nx8877)) ;
    and04 ix8407 (.Y (nx8406), .A0 (nx8408), .A1 (nx8410), .A2 (nx8412), .A3 (
          nx8414)) ;
    aoi22 ix8409 (.Y (nx8408), .A0 (nx3050), .A1 (nx8869), .B0 (nx3100), .B1 (
          nx8865)) ;
    aoi22 ix8411 (.Y (nx8410), .A0 (nx3026), .A1 (nx8861), .B0 (nx3076), .B1 (
          nx8857)) ;
    aoi22 ix8413 (.Y (nx8412), .A0 (nx2794), .A1 (nx8853), .B0 (nx2820), .B1 (
          nx8849)) ;
    aoi22 ix8415 (.Y (nx8414), .A0 (nx3000), .A1 (nx8845), .B0 (nx5286), .B1 (
          nx8841)) ;
    mux21_ni ix5287 (.Y (nx5286), .A0 (Mem_2__7), .A1 (Mem_3__7), .S0 (
             Address[0])) ;
    dff reg_Mem_2__7 (.Q (Mem_2__7), .QB (\$dummy [239]), .D (nx6765), .CLK (CLK
        )) ;
    mux21_ni ix6766 (.Y (nx6765), .A0 (Din[7]), .A1 (Mem_2__7), .S0 (nx9021)) ;
    or02 ix5553 (.Y (Dout[24]), .A0 (nx5550), .A1 (nx5466)) ;
    nand04 ix5551 (.Y (nx5550), .A0 (nx8422), .A1 (nx8442), .A2 (nx8452), .A3 (
           nx8466)) ;
    aoi22 ix8423 (.Y (nx8422), .A0 (nx3260), .A1 (nx5542), .B0 (nx3376), .B1 (
          nx5538)) ;
    and02 ix5543 (.Y (nx5542), .A0 (nx5406), .A1 (nx5434)) ;
    nor02_2x ix5407 (.Y (nx5406), .A0 (nx9081), .A1 (nx5366)) ;
    xnor2_2x ix5367 (.Y (nx5366), .A0 (Address[4]), .A1 (nx8427)) ;
    nand02 ix8428 (.Y (nx8427), .A0 (Address[3]), .A1 (nx5346)) ;
    aoi21 ix5353 (.Y (nx5352), .A0 (nx8993), .A1 (nx8975), .B0 (nx5346)) ;
    xnor2 ix8433 (.Y (nx8432), .A0 (Address[3]), .A1 (nx5346)) ;
    nor03_2x ix5539 (.Y (nx5538), .A0 (nx8435), .A1 (nx8815), .A2 (nx5366)) ;
    aoi22 ix8443 (.Y (nx8442), .A0 (nx3184), .A1 (nx9059), .B0 (nx3120), .B1 (
          nx5526)) ;
    nand02 ix8446 (.Y (nx8445), .A0 (nx8815), .A1 (nx5366)) ;
    aoi22 ix8453 (.Y (nx8452), .A0 (Mem_1__0), .A1 (nx8921), .B0 (nx3354), .B1 (
          nx5512)) ;
    dff reg_Mem_1__0 (.Q (Mem_1__0), .QB (\$dummy [240]), .D (nx6775), .CLK (CLK
        )) ;
    mux21_ni ix6776 (.Y (nx6775), .A0 (Din[0]), .A1 (Mem_1__0), .S0 (nx9025)) ;
    nand02 ix8457 (.Y (nx8456), .A0 (WR), .A1 (nx9123)) ;
    nor04 ix5507 (.Y (nx5506), .A0 (Address[0]), .A1 (Address[1]), .A2 (nx5366)
          , .A3 (nx8463)) ;
    nor03_2x ix5513 (.Y (nx5512), .A0 (nx8445), .A1 (nx8437), .A2 (nx9023)) ;
    aoi22 ix8467 (.Y (nx8466), .A0 (nx3162), .A1 (nx5472), .B0 (Mem_2__0), .B1 (
          nx8915)) ;
    nor03_2x ix5473 (.Y (nx5472), .A0 (nx8445), .A1 (nx8437), .A2 (nx5364)) ;
    nor04 ix5479 (.Y (nx5478), .A0 (nx8463), .A1 (nx6958), .A2 (Address[1]), .A3 (
          Address[4])) ;
    nand04 ix5467 (.Y (nx5466), .A0 (nx8471), .A1 (nx8475), .A2 (nx8481), .A3 (
           nx8485)) ;
    aoi22 ix8472 (.Y (nx8471), .A0 (nx3242), .A1 (nx5458), .B0 (nx3204), .B1 (
          nx5450)) ;
    and03 ix5459 (.Y (nx5458), .A0 (nx5406), .A1 (nx9057), .A2 (nx9023)) ;
    nor03_2x ix5451 (.Y (nx5450), .A0 (nx8463), .A1 (nx8815), .A2 (nx8450)) ;
    aoi22 ix8476 (.Y (nx8475), .A0 (nx3272), .A1 (nx5428), .B0 (nx3392), .B1 (
          nx5440)) ;
    nor03_2x ix5429 (.Y (nx5428), .A0 (nx8478), .A1 (nx9023), .A2 (nx8450)) ;
    nand02 ix8479 (.Y (nx8478), .A0 (nx9081), .A1 (nx9057)) ;
    aoi22 ix8482 (.Y (nx8481), .A0 (nx3224), .A1 (nx5418), .B0 (Mem_3__0), .B1 (
          nx8911)) ;
    nor02_2x ix5419 (.Y (nx5418), .A0 (nx8463), .A1 (nx8445)) ;
    nor04 ix5413 (.Y (nx5412), .A0 (Address[2]), .A1 (Address[0]), .A2 (
          Address[3]), .A3 (nx8448)) ;
    aoi222 ix8486 (.Y (nx8485), .A0 (nx3294), .A1 (nx8899), .B0 (nx3406), .B1 (
           nx8903), .C0 (nx3342), .C1 (nx8907)) ;
    nor03_2x ix5373 (.Y (nx5372), .A0 (nx8478), .A1 (nx9023), .A2 (nx5366)) ;
    nor03_2x ix5383 (.Y (nx5382), .A0 (nx8478), .A1 (nx5364), .A2 (nx5366)) ;
    nor03_2x ix5391 (.Y (nx5390), .A0 (nx8478), .A1 (nx5364), .A2 (nx8450)) ;
    or02 ix5625 (.Y (Dout[25]), .A0 (nx5622), .A1 (nx5586)) ;
    nand04 ix5623 (.Y (nx5622), .A0 (nx8492), .A1 (nx8494), .A2 (nx8496), .A3 (
           nx8501)) ;
    aoi22 ix8493 (.Y (nx8492), .A0 (nx3500), .A1 (nx5542), .B0 (nx3570), .B1 (
          nx5538)) ;
    aoi22 ix8495 (.Y (nx8494), .A0 (nx3454), .A1 (nx9059), .B0 (nx3432), .B1 (
          nx5526)) ;
    aoi22 ix8497 (.Y (nx8496), .A0 (Mem_1__1), .A1 (nx8921), .B0 (nx3556), .B1 (
          nx5512)) ;
    dff reg_Mem_1__1 (.Q (Mem_1__1), .QB (\$dummy [241]), .D (nx6785), .CLK (CLK
        )) ;
    mux21_ni ix6786 (.Y (nx6785), .A0 (Din[1]), .A1 (Mem_1__1), .S0 (nx9025)) ;
    aoi22 ix8502 (.Y (nx8501), .A0 (nx3442), .A1 (nx5472), .B0 (Mem_2__1), .B1 (
          nx8915)) ;
    nand04 ix5587 (.Y (nx5586), .A0 (nx8504), .A1 (nx8506), .A2 (nx8508), .A3 (
           nx8510)) ;
    aoi22 ix8505 (.Y (nx8504), .A0 (nx3488), .A1 (nx5458), .B0 (nx3464), .B1 (
          nx5450)) ;
    aoi22 ix8507 (.Y (nx8506), .A0 (nx3510), .A1 (nx5428), .B0 (nx3580), .B1 (
          nx5440)) ;
    aoi22 ix8509 (.Y (nx8508), .A0 (nx3478), .A1 (nx5418), .B0 (Mem_3__1), .B1 (
          nx8911)) ;
    aoi222 ix8511 (.Y (nx8510), .A0 (nx3526), .A1 (nx8899), .B0 (nx3590), .B1 (
           nx8903), .C0 (nx3546), .C1 (nx8907)) ;
    or02 ix5697 (.Y (Dout[26]), .A0 (nx5694), .A1 (nx5658)) ;
    nand04 ix5695 (.Y (nx5694), .A0 (nx8514), .A1 (nx8516), .A2 (nx8518), .A3 (
           nx8523)) ;
    aoi22 ix8515 (.Y (nx8514), .A0 (nx3676), .A1 (nx5542), .B0 (nx3746), .B1 (
          nx5538)) ;
    aoi22 ix8517 (.Y (nx8516), .A0 (nx3630), .A1 (nx9059), .B0 (nx3608), .B1 (
          nx5526)) ;
    aoi22 ix8519 (.Y (nx8518), .A0 (Mem_1__2), .A1 (nx8921), .B0 (nx3732), .B1 (
          nx5512)) ;
    dff reg_Mem_1__2 (.Q (Mem_1__2), .QB (\$dummy [242]), .D (nx6795), .CLK (CLK
        )) ;
    mux21_ni ix6796 (.Y (nx6795), .A0 (Din[2]), .A1 (Mem_1__2), .S0 (nx9025)) ;
    aoi22 ix8524 (.Y (nx8523), .A0 (nx3618), .A1 (nx5472), .B0 (Mem_2__2), .B1 (
          nx8915)) ;
    nand04 ix5659 (.Y (nx5658), .A0 (nx8526), .A1 (nx8528), .A2 (nx8530), .A3 (
           nx8532)) ;
    aoi22 ix8527 (.Y (nx8526), .A0 (nx3664), .A1 (nx5458), .B0 (nx3640), .B1 (
          nx5450)) ;
    aoi22 ix8529 (.Y (nx8528), .A0 (nx3686), .A1 (nx5428), .B0 (nx3756), .B1 (
          nx5440)) ;
    aoi22 ix8531 (.Y (nx8530), .A0 (nx3654), .A1 (nx5418), .B0 (Mem_3__2), .B1 (
          nx8911)) ;
    aoi222 ix8533 (.Y (nx8532), .A0 (nx3702), .A1 (nx8899), .B0 (nx3766), .B1 (
           nx8903), .C0 (nx3722), .C1 (nx8907)) ;
    or02 ix5769 (.Y (Dout[27]), .A0 (nx5766), .A1 (nx5730)) ;
    nand04 ix5767 (.Y (nx5766), .A0 (nx8536), .A1 (nx8538), .A2 (nx8540), .A3 (
           nx8545)) ;
    aoi22 ix8537 (.Y (nx8536), .A0 (nx3852), .A1 (nx5542), .B0 (nx3922), .B1 (
          nx5538)) ;
    aoi22 ix8539 (.Y (nx8538), .A0 (nx3806), .A1 (nx9059), .B0 (nx3784), .B1 (
          nx5526)) ;
    aoi22 ix8541 (.Y (nx8540), .A0 (Mem_1__3), .A1 (nx8921), .B0 (nx3908), .B1 (
          nx5512)) ;
    dff reg_Mem_1__3 (.Q (Mem_1__3), .QB (\$dummy [243]), .D (nx6805), .CLK (CLK
        )) ;
    mux21_ni ix6806 (.Y (nx6805), .A0 (Din[3]), .A1 (Mem_1__3), .S0 (nx9025)) ;
    aoi22 ix8546 (.Y (nx8545), .A0 (nx3794), .A1 (nx5472), .B0 (Mem_2__3), .B1 (
          nx8915)) ;
    nand04 ix5731 (.Y (nx5730), .A0 (nx8548), .A1 (nx8550), .A2 (nx8552), .A3 (
           nx8554)) ;
    aoi22 ix8549 (.Y (nx8548), .A0 (nx3840), .A1 (nx5458), .B0 (nx3816), .B1 (
          nx5450)) ;
    aoi22 ix8551 (.Y (nx8550), .A0 (nx3862), .A1 (nx5428), .B0 (nx3932), .B1 (
          nx5440)) ;
    aoi22 ix8553 (.Y (nx8552), .A0 (nx3830), .A1 (nx5418), .B0 (Mem_3__3), .B1 (
          nx8911)) ;
    aoi222 ix8555 (.Y (nx8554), .A0 (nx3878), .A1 (nx8899), .B0 (nx3942), .B1 (
           nx8903), .C0 (nx3898), .C1 (nx8907)) ;
    or02 ix5841 (.Y (Dout[28]), .A0 (nx5838), .A1 (nx5802)) ;
    nand04 ix5839 (.Y (nx5838), .A0 (nx8558), .A1 (nx8560), .A2 (nx8562), .A3 (
           nx8567)) ;
    aoi22 ix8559 (.Y (nx8558), .A0 (nx4028), .A1 (nx5542), .B0 (nx4098), .B1 (
          nx5538)) ;
    aoi22 ix8561 (.Y (nx8560), .A0 (nx3982), .A1 (nx9059), .B0 (nx3960), .B1 (
          nx5526)) ;
    aoi22 ix8563 (.Y (nx8562), .A0 (Mem_1__4), .A1 (nx8921), .B0 (nx4084), .B1 (
          nx5512)) ;
    dff reg_Mem_1__4 (.Q (Mem_1__4), .QB (\$dummy [244]), .D (nx6815), .CLK (CLK
        )) ;
    mux21_ni ix6816 (.Y (nx6815), .A0 (Din[4]), .A1 (Mem_1__4), .S0 (nx9025)) ;
    aoi22 ix8568 (.Y (nx8567), .A0 (nx3970), .A1 (nx5472), .B0 (Mem_2__4), .B1 (
          nx8915)) ;
    nand04 ix5803 (.Y (nx5802), .A0 (nx8570), .A1 (nx8572), .A2 (nx8574), .A3 (
           nx8576)) ;
    aoi22 ix8571 (.Y (nx8570), .A0 (nx4016), .A1 (nx5458), .B0 (nx3992), .B1 (
          nx5450)) ;
    aoi22 ix8573 (.Y (nx8572), .A0 (nx4038), .A1 (nx5428), .B0 (nx4108), .B1 (
          nx5440)) ;
    aoi22 ix8575 (.Y (nx8574), .A0 (nx4006), .A1 (nx5418), .B0 (Mem_3__4), .B1 (
          nx8911)) ;
    aoi222 ix8577 (.Y (nx8576), .A0 (nx4054), .A1 (nx8899), .B0 (nx4118), .B1 (
           nx8903), .C0 (nx4074), .C1 (nx8907)) ;
    or02 ix5913 (.Y (Dout[29]), .A0 (nx5910), .A1 (nx5874)) ;
    nand04 ix5911 (.Y (nx5910), .A0 (nx8580), .A1 (nx8582), .A2 (nx8584), .A3 (
           nx8589)) ;
    aoi22 ix8581 (.Y (nx8580), .A0 (nx4204), .A1 (nx5542), .B0 (nx4274), .B1 (
          nx5538)) ;
    aoi22 ix8583 (.Y (nx8582), .A0 (nx4158), .A1 (nx9059), .B0 (nx4136), .B1 (
          nx5526)) ;
    aoi22 ix8585 (.Y (nx8584), .A0 (Mem_1__5), .A1 (nx8921), .B0 (nx4260), .B1 (
          nx5512)) ;
    dff reg_Mem_1__5 (.Q (Mem_1__5), .QB (\$dummy [245]), .D (nx6825), .CLK (CLK
        )) ;
    mux21_ni ix6826 (.Y (nx6825), .A0 (Din[5]), .A1 (Mem_1__5), .S0 (nx9025)) ;
    aoi22 ix8590 (.Y (nx8589), .A0 (nx4146), .A1 (nx5472), .B0 (Mem_2__5), .B1 (
          nx8915)) ;
    nand04 ix5875 (.Y (nx5874), .A0 (nx8592), .A1 (nx8594), .A2 (nx8596), .A3 (
           nx8598)) ;
    aoi22 ix8593 (.Y (nx8592), .A0 (nx4192), .A1 (nx5458), .B0 (nx4168), .B1 (
          nx5450)) ;
    aoi22 ix8595 (.Y (nx8594), .A0 (nx4214), .A1 (nx5428), .B0 (nx4284), .B1 (
          nx5440)) ;
    aoi22 ix8597 (.Y (nx8596), .A0 (nx4182), .A1 (nx5418), .B0 (Mem_3__5), .B1 (
          nx8911)) ;
    aoi222 ix8599 (.Y (nx8598), .A0 (nx4230), .A1 (nx8899), .B0 (nx4294), .B1 (
           nx8903), .C0 (nx4250), .C1 (nx8907)) ;
    or02 ix5985 (.Y (Dout[30]), .A0 (nx5982), .A1 (nx5946)) ;
    nand04 ix5983 (.Y (nx5982), .A0 (nx8602), .A1 (nx8604), .A2 (nx8606), .A3 (
           nx8611)) ;
    aoi22 ix8603 (.Y (nx8602), .A0 (nx4380), .A1 (nx5542), .B0 (nx4450), .B1 (
          nx5538)) ;
    aoi22 ix8605 (.Y (nx8604), .A0 (nx4334), .A1 (nx9059), .B0 (nx4312), .B1 (
          nx5526)) ;
    aoi22 ix8607 (.Y (nx8606), .A0 (Mem_1__6), .A1 (nx8921), .B0 (nx4436), .B1 (
          nx5512)) ;
    dff reg_Mem_1__6 (.Q (Mem_1__6), .QB (\$dummy [246]), .D (nx6835), .CLK (CLK
        )) ;
    mux21_ni ix6836 (.Y (nx6835), .A0 (Din[6]), .A1 (Mem_1__6), .S0 (nx9025)) ;
    aoi22 ix8612 (.Y (nx8611), .A0 (nx4322), .A1 (nx5472), .B0 (Mem_2__6), .B1 (
          nx8915)) ;
    nand04 ix5947 (.Y (nx5946), .A0 (nx8614), .A1 (nx8616), .A2 (nx8618), .A3 (
           nx8620)) ;
    aoi22 ix8615 (.Y (nx8614), .A0 (nx4368), .A1 (nx5458), .B0 (nx4344), .B1 (
          nx5450)) ;
    aoi22 ix8617 (.Y (nx8616), .A0 (nx4390), .A1 (nx5428), .B0 (nx4460), .B1 (
          nx5440)) ;
    aoi22 ix8619 (.Y (nx8618), .A0 (nx4358), .A1 (nx5418), .B0 (Mem_3__6), .B1 (
          nx8911)) ;
    aoi222 ix8621 (.Y (nx8620), .A0 (nx4406), .A1 (nx8899), .B0 (nx4470), .B1 (
           nx8903), .C0 (nx4426), .C1 (nx8907)) ;
    or02 ix6057 (.Y (Dout[31]), .A0 (nx6054), .A1 (nx6018)) ;
    nand04 ix6055 (.Y (nx6054), .A0 (nx8624), .A1 (nx8626), .A2 (nx8628), .A3 (
           nx8633)) ;
    aoi22 ix8625 (.Y (nx8624), .A0 (nx4556), .A1 (nx5542), .B0 (nx4626), .B1 (
          nx5538)) ;
    aoi22 ix8627 (.Y (nx8626), .A0 (nx4510), .A1 (nx9061), .B0 (nx4488), .B1 (
          nx5526)) ;
    aoi22 ix8629 (.Y (nx8628), .A0 (Mem_1__7), .A1 (nx8923), .B0 (nx4612), .B1 (
          nx5512)) ;
    dff reg_Mem_1__7 (.Q (Mem_1__7), .QB (\$dummy [247]), .D (nx6845), .CLK (CLK
        )) ;
    mux21_ni ix6846 (.Y (nx6845), .A0 (Din[7]), .A1 (Mem_1__7), .S0 (nx9027)) ;
    aoi22 ix8634 (.Y (nx8633), .A0 (nx4498), .A1 (nx5472), .B0 (Mem_2__7), .B1 (
          nx8917)) ;
    nand04 ix6019 (.Y (nx6018), .A0 (nx8636), .A1 (nx8638), .A2 (nx8640), .A3 (
           nx8642)) ;
    aoi22 ix8637 (.Y (nx8636), .A0 (nx4544), .A1 (nx5458), .B0 (nx4520), .B1 (
          nx5450)) ;
    aoi22 ix8639 (.Y (nx8638), .A0 (nx4566), .A1 (nx5428), .B0 (nx4636), .B1 (
          nx5440)) ;
    aoi22 ix8641 (.Y (nx8640), .A0 (nx4534), .A1 (nx5418), .B0 (Mem_3__7), .B1 (
          nx8913)) ;
    aoi222 ix8643 (.Y (nx8642), .A0 (nx4582), .A1 (nx8901), .B0 (nx4646), .B1 (
           nx8905), .C0 (nx4602), .C1 (nx8909)) ;
    nand04 ix6123 (.Y (Dout[32]), .A0 (nx8645), .A1 (nx8647), .A2 (nx8655), .A3 (
           nx8659)) ;
    aoi22 ix8646 (.Y (nx8645), .A0 (nx332), .A1 (nx8761), .B0 (nx180), .B1 (
          nx8763)) ;
    aoi222 ix8648 (.Y (nx8647), .A0 (Mem_0__0), .A1 (nx9125), .B0 (Mem_1__0), .B1 (
           nx9123), .C0 (nx416), .C1 (nx8789)) ;
    dff reg_Mem_0__0 (.Q (Mem_0__0), .QB (\$dummy [248]), .D (nx6855), .CLK (CLK
        )) ;
    mux21_ni ix6856 (.Y (nx6855), .A0 (Din[0]), .A1 (Mem_0__0), .S0 (nx9029)) ;
    nand02 ix8652 (.Y (nx8651), .A0 (WR), .A1 (nx9125)) ;
    aoi22 ix8656 (.Y (nx8655), .A0 (nx564), .A1 (nx9063), .B0 (nx260), .B1 (
          nx6080)) ;
    nor03_2x ix6081 (.Y (nx6080), .A0 (nx8961), .A1 (Address[2]), .A2 (
             Address[3])) ;
    aoi222 ix8660 (.Y (nx8659), .A0 (nx4676), .A1 (nx8925), .B0 (nx82), .B1 (
           nx8933), .C0 (nx490), .C1 (nx8929)) ;
    nor03_2x ix6071 (.Y (nx6070), .A0 (nx8961), .A1 (Address[2]), .A2 (nx8965)
             ) ;
    nor03_2x ix6065 (.Y (nx6064), .A0 (nx8961), .A1 (nx8975), .A2 (Address[3])
             ) ;
    nand04 ix6167 (.Y (Dout[33]), .A0 (nx8665), .A1 (nx8667), .A2 (nx8672), .A3 (
           nx8674)) ;
    aoi22 ix8666 (.Y (nx8665), .A0 (nx778), .A1 (nx8761), .B0 (nx676), .B1 (
          nx8763)) ;
    aoi222 ix8668 (.Y (nx8667), .A0 (Mem_0__1), .A1 (nx9125), .B0 (Mem_1__1), .B1 (
           nx9123), .C0 (nx832), .C1 (nx8789)) ;
    dff reg_Mem_0__1 (.Q (Mem_0__1), .QB (\$dummy [249]), .D (nx6865), .CLK (CLK
        )) ;
    mux21_ni ix6866 (.Y (nx6865), .A0 (Din[1]), .A1 (Mem_0__1), .S0 (nx9029)) ;
    aoi22 ix8673 (.Y (nx8672), .A0 (nx932), .A1 (nx9063), .B0 (nx728), .B1 (
          nx6080)) ;
    aoi222 ix8675 (.Y (nx8674), .A0 (nx4854), .A1 (nx8925), .B0 (nx626), .B1 (
           nx8933), .C0 (nx882), .C1 (nx8929)) ;
    nand04 ix6211 (.Y (Dout[34]), .A0 (nx8677), .A1 (nx8679), .A2 (nx8684), .A3 (
           nx8686)) ;
    aoi22 ix8678 (.Y (nx8677), .A0 (nx1140), .A1 (nx8761), .B0 (nx1038), .B1 (
          nx8763)) ;
    aoi222 ix8680 (.Y (nx8679), .A0 (Mem_0__2), .A1 (nx9125), .B0 (Mem_1__2), .B1 (
           nx9123), .C0 (nx1194), .C1 (nx8789)) ;
    dff reg_Mem_0__2 (.Q (Mem_0__2), .QB (\$dummy [250]), .D (nx6875), .CLK (CLK
        )) ;
    mux21_ni ix6876 (.Y (nx6875), .A0 (Din[2]), .A1 (Mem_0__2), .S0 (nx9029)) ;
    aoi22 ix8685 (.Y (nx8684), .A0 (nx1294), .A1 (nx9063), .B0 (nx1090), .B1 (
          nx6080)) ;
    aoi222 ix8687 (.Y (nx8686), .A0 (nx4926), .A1 (nx8925), .B0 (nx988), .B1 (
           nx8933), .C0 (nx1244), .C1 (nx8929)) ;
    nand04 ix6255 (.Y (Dout[35]), .A0 (nx8689), .A1 (nx8691), .A2 (nx8696), .A3 (
           nx8698)) ;
    aoi22 ix8690 (.Y (nx8689), .A0 (nx1502), .A1 (nx8761), .B0 (nx1400), .B1 (
          nx8763)) ;
    aoi222 ix8692 (.Y (nx8691), .A0 (Mem_0__3), .A1 (nx9125), .B0 (Mem_1__3), .B1 (
           nx9123), .C0 (nx1556), .C1 (nx8789)) ;
    dff reg_Mem_0__3 (.Q (Mem_0__3), .QB (\$dummy [251]), .D (nx6885), .CLK (CLK
        )) ;
    mux21_ni ix6886 (.Y (nx6885), .A0 (Din[3]), .A1 (Mem_0__3), .S0 (nx9029)) ;
    aoi22 ix8697 (.Y (nx8696), .A0 (nx1656), .A1 (nx9063), .B0 (nx1452), .B1 (
          nx6080)) ;
    aoi222 ix8699 (.Y (nx8698), .A0 (nx4998), .A1 (nx8925), .B0 (nx1350), .B1 (
           nx8933), .C0 (nx1606), .C1 (nx8929)) ;
    nand04 ix6299 (.Y (Dout[36]), .A0 (nx8701), .A1 (nx8703), .A2 (nx8708), .A3 (
           nx8710)) ;
    aoi22 ix8702 (.Y (nx8701), .A0 (nx1864), .A1 (nx8761), .B0 (nx1762), .B1 (
          nx8763)) ;
    aoi222 ix8704 (.Y (nx8703), .A0 (Mem_0__4), .A1 (nx9125), .B0 (Mem_1__4), .B1 (
           nx9123), .C0 (nx1918), .C1 (nx8789)) ;
    dff reg_Mem_0__4 (.Q (Mem_0__4), .QB (\$dummy [252]), .D (nx6895), .CLK (CLK
        )) ;
    mux21_ni ix6896 (.Y (nx6895), .A0 (Din[4]), .A1 (Mem_0__4), .S0 (nx9029)) ;
    aoi22 ix8709 (.Y (nx8708), .A0 (nx2018), .A1 (nx9063), .B0 (nx1814), .B1 (
          nx6080)) ;
    aoi222 ix8711 (.Y (nx8710), .A0 (nx5070), .A1 (nx8925), .B0 (nx1712), .B1 (
           nx8933), .C0 (nx1968), .C1 (nx8929)) ;
    nand04 ix6343 (.Y (Dout[37]), .A0 (nx8713), .A1 (nx8715), .A2 (nx8720), .A3 (
           nx8722)) ;
    aoi22 ix8714 (.Y (nx8713), .A0 (nx2226), .A1 (nx88), .B0 (nx2124), .B1 (
          nx8763)) ;
    aoi222 ix8716 (.Y (nx8715), .A0 (Mem_0__5), .A1 (nx6098), .B0 (Mem_1__5), .B1 (
           nx9123), .C0 (nx2280), .C1 (nx8789)) ;
    dff reg_Mem_0__5 (.Q (Mem_0__5), .QB (\$dummy [253]), .D (nx6905), .CLK (CLK
        )) ;
    mux21_ni ix6906 (.Y (nx6905), .A0 (Din[5]), .A1 (Mem_0__5), .S0 (nx9029)) ;
    aoi22 ix8721 (.Y (nx8720), .A0 (nx2380), .A1 (nx9063), .B0 (nx2176), .B1 (
          nx6080)) ;
    aoi222 ix8723 (.Y (nx8722), .A0 (nx5142), .A1 (nx8925), .B0 (nx2074), .B1 (
           nx8933), .C0 (nx2330), .C1 (nx8929)) ;
    nand04 ix6387 (.Y (Dout[38]), .A0 (nx8725), .A1 (nx8727), .A2 (nx8732), .A3 (
           nx8734)) ;
    aoi22 ix8726 (.Y (nx8725), .A0 (nx2588), .A1 (nx88), .B0 (nx2486), .B1 (
          nx8765)) ;
    aoi222 ix8728 (.Y (nx8727), .A0 (Mem_0__6), .A1 (nx6098), .B0 (Mem_1__6), .B1 (
           nx5486), .C0 (nx2642), .C1 (nx8791)) ;
    dff reg_Mem_0__6 (.Q (Mem_0__6), .QB (\$dummy [254]), .D (nx6915), .CLK (CLK
        )) ;
    mux21_ni ix6916 (.Y (nx6915), .A0 (Din[6]), .A1 (Mem_0__6), .S0 (nx9029)) ;
    aoi22 ix8733 (.Y (nx8732), .A0 (nx2742), .A1 (nx9063), .B0 (nx2538), .B1 (
          nx6080)) ;
    aoi222 ix8735 (.Y (nx8734), .A0 (nx5214), .A1 (nx8925), .B0 (nx2436), .B1 (
           nx8933), .C0 (nx2692), .C1 (nx8929)) ;
    nand04 ix6431 (.Y (Dout[39]), .A0 (nx8737), .A1 (nx8739), .A2 (nx8744), .A3 (
           nx8746)) ;
    aoi22 ix8738 (.Y (nx8737), .A0 (nx2950), .A1 (nx88), .B0 (nx2848), .B1 (
          nx8765)) ;
    aoi222 ix8740 (.Y (nx8739), .A0 (Mem_0__7), .A1 (nx6098), .B0 (Mem_1__7), .B1 (
           nx5486), .C0 (nx3004), .C1 (nx8791)) ;
    dff reg_Mem_0__7 (.Q (Mem_0__7), .QB (\$dummy [255]), .D (nx6925), .CLK (CLK
        )) ;
    mux21_ni ix6926 (.Y (nx6925), .A0 (Din[7]), .A1 (Mem_0__7), .S0 (nx9031)) ;
    aoi22 ix8745 (.Y (nx8744), .A0 (nx3104), .A1 (nx9065), .B0 (nx2900), .B1 (
          nx6080)) ;
    aoi222 ix8747 (.Y (nx8746), .A0 (nx5286), .A1 (nx8927), .B0 (nx2798), .B1 (
           nx8935), .C0 (nx3054), .C1 (nx8931)) ;
    inv01 ix8436 (.Y (nx8435), .A (nx5434)) ;
    inv01 ix8449 (.Y (nx8448), .A (nx5406)) ;
    inv02 ix8451 (.Y (nx8450), .A (nx5366)) ;
    inv02 ix5365 (.Y (nx5364), .A (nx8432)) ;
    inv01 ix8438 (.Y (nx8437), .A (nx5352)) ;
    inv01 ix7940 (.Y (nx7939), .A (nx3188)) ;
    inv02 ix3149 (.Y (nx3148), .A (nx7926)) ;
    inv01 ix7969 (.Y (nx7968), .A (nx3136)) ;
    inv01 ix7956 (.Y (nx7955), .A (nx3126)) ;
    inv01 ix67 (.Y (nx66), .A (nx7033)) ;
    nor02_2x ix8760 (.Y (nx8761), .A0 (Address[4]), .A1 (nx6947)) ;
    buf02 ix8762 (.Y (nx8763), .A (nx116)) ;
    buf02 ix8764 (.Y (nx8765), .A (nx116)) ;
    buf02 ix8788 (.Y (nx8789), .A (nx352)) ;
    buf02 ix8790 (.Y (nx8791), .A (nx352)) ;
    buf02 ix8800 (.Y (nx8801), .A (nx422)) ;
    buf02 ix8802 (.Y (nx8803), .A (nx422)) ;
    buf02 ix8804 (.Y (nx8805), .A (nx498)) ;
    buf02 ix8806 (.Y (nx8807), .A (nx498)) ;
    buf02 ix8808 (.Y (nx8809), .A (nx570)) ;
    buf02 ix8810 (.Y (nx8811), .A (nx570)) ;
    inv02 ix8812 (.Y (nx8813), .A (nx7945)) ;
    inv02 ix8814 (.Y (nx8815), .A (nx9081)) ;
    inv02 ix8816 (.Y (nx8817), .A (nx7941)) ;
    buf02 ix8818 (.Y (nx8819), .A (nx3330)) ;
    buf02 ix8820 (.Y (nx8821), .A (nx3330)) ;
    buf02 ix8822 (.Y (nx8823), .A (nx3362)) ;
    buf02 ix8824 (.Y (nx8825), .A (nx3362)) ;
    buf02 ix8826 (.Y (nx8827), .A (nx3382)) ;
    buf02 ix8828 (.Y (nx8829), .A (nx3382)) ;
    buf02 ix8830 (.Y (nx8831), .A (nx3396)) ;
    buf02 ix8832 (.Y (nx8833), .A (nx3396)) ;
    buf02 ix8834 (.Y (nx8835), .A (nx3414)) ;
    buf02 ix8836 (.Y (nx8837), .A (nx3414)) ;
    buf02 ix8838 (.Y (nx8839), .A (nx4708)) ;
    buf02 ix8840 (.Y (nx8841), .A (nx4708)) ;
    buf02 ix8842 (.Y (nx8843), .A (nx4716)) ;
    buf02 ix8844 (.Y (nx8845), .A (nx4716)) ;
    buf02 ix8846 (.Y (nx8847), .A (nx4724)) ;
    buf02 ix8848 (.Y (nx8849), .A (nx4724)) ;
    buf02 ix8850 (.Y (nx8851), .A (nx4730)) ;
    buf02 ix8852 (.Y (nx8853), .A (nx4730)) ;
    buf02 ix8854 (.Y (nx8855), .A (nx4742)) ;
    buf02 ix8856 (.Y (nx8857), .A (nx4742)) ;
    buf02 ix8858 (.Y (nx8859), .A (nx4752)) ;
    buf02 ix8860 (.Y (nx8861), .A (nx4752)) ;
    buf02 ix8862 (.Y (nx8863), .A (nx4764)) ;
    buf02 ix8864 (.Y (nx8865), .A (nx4764)) ;
    buf02 ix8866 (.Y (nx8867), .A (nx4768)) ;
    buf02 ix8868 (.Y (nx8869), .A (nx4768)) ;
    buf02 ix8870 (.Y (nx8871), .A (nx4782)) ;
    buf02 ix8872 (.Y (nx8873), .A (nx4782)) ;
    buf02 ix8874 (.Y (nx8875), .A (nx4792)) ;
    buf02 ix8876 (.Y (nx8877), .A (nx4792)) ;
    buf02 ix8878 (.Y (nx8879), .A (nx4798)) ;
    buf02 ix8880 (.Y (nx8881), .A (nx4798)) ;
    buf02 ix8882 (.Y (nx8883), .A (nx4806)) ;
    buf02 ix8884 (.Y (nx8885), .A (nx4806)) ;
    buf02 ix8886 (.Y (nx8887), .A (nx4814)) ;
    buf02 ix8888 (.Y (nx8889), .A (nx4814)) ;
    buf02 ix8890 (.Y (nx8891), .A (nx4822)) ;
    buf02 ix8892 (.Y (nx8893), .A (nx4822)) ;
    buf02 ix8894 (.Y (nx8895), .A (nx4830)) ;
    buf02 ix8896 (.Y (nx8897), .A (nx4830)) ;
    buf02 ix8898 (.Y (nx8899), .A (nx5372)) ;
    buf02 ix8900 (.Y (nx8901), .A (nx5372)) ;
    buf02 ix8902 (.Y (nx8903), .A (nx5382)) ;
    buf02 ix8904 (.Y (nx8905), .A (nx5382)) ;
    buf02 ix8906 (.Y (nx8907), .A (nx5390)) ;
    buf02 ix8908 (.Y (nx8909), .A (nx5390)) ;
    buf02 ix8910 (.Y (nx8911), .A (nx5412)) ;
    buf02 ix8912 (.Y (nx8913), .A (nx5412)) ;
    buf02 ix8914 (.Y (nx8915), .A (nx5478)) ;
    buf02 ix8916 (.Y (nx8917), .A (nx5478)) ;
    buf02 ix8920 (.Y (nx8921), .A (nx5506)) ;
    buf02 ix8922 (.Y (nx8923), .A (nx5506)) ;
    buf02 ix8924 (.Y (nx8925), .A (nx6058)) ;
    buf02 ix8926 (.Y (nx8927), .A (nx6058)) ;
    buf02 ix8928 (.Y (nx8929), .A (nx6064)) ;
    buf02 ix8930 (.Y (nx8931), .A (nx6064)) ;
    buf02 ix8932 (.Y (nx8933), .A (nx6070)) ;
    buf02 ix8934 (.Y (nx8935), .A (nx6070)) ;
    buf02 ix8938 (.Y (nx8939), .A (nx6942)) ;
    buf02 ix8940 (.Y (nx8941), .A (nx6942)) ;
    buf02 ix8942 (.Y (nx8943), .A (nx6954)) ;
    buf02 ix8944 (.Y (nx8945), .A (nx6954)) ;
    buf02 ix8946 (.Y (nx8947), .A (nx6964)) ;
    buf02 ix8948 (.Y (nx8949), .A (nx6964)) ;
    inv02 ix8950 (.Y (nx8951), .A (Address[1])) ;
    buf02 ix8954 (.Y (nx8955), .A (nx6973)) ;
    buf02 ix8956 (.Y (nx8957), .A (nx6973)) ;
    inv04 ix8958 (.Y (nx8959), .A (Address[4])) ;
    inv04 ix8960 (.Y (nx8961), .A (Address[4])) ;
    inv04 ix8962 (.Y (nx8963), .A (Address[3])) ;
    inv04 ix8964 (.Y (nx8965), .A (Address[3])) ;
    buf02 ix8966 (.Y (nx8967), .A (nx6986)) ;
    buf02 ix8968 (.Y (nx8969), .A (nx6986)) ;
    inv02 ix8970 (.Y (nx8971), .A (Address[2])) ;
    inv02 ix8972 (.Y (nx8973), .A (Address[2])) ;
    inv02 ix8974 (.Y (nx8975), .A (Address[2])) ;
    buf02 ix8976 (.Y (nx8977), .A (nx6994)) ;
    buf02 ix8978 (.Y (nx8979), .A (nx6994)) ;
    buf02 ix8980 (.Y (nx8981), .A (nx7000)) ;
    buf02 ix8982 (.Y (nx8983), .A (nx7000)) ;
    buf02 ix8984 (.Y (nx8985), .A (nx7005)) ;
    buf02 ix8986 (.Y (nx8987), .A (nx7005)) ;
    buf02 ix8988 (.Y (nx8989), .A (nx7015)) ;
    buf02 ix8990 (.Y (nx8991), .A (nx7015)) ;
    inv02 ix8992 (.Y (nx8993), .A (nx9049)) ;
    buf02 ix8996 (.Y (nx8997), .A (nx7050)) ;
    buf02 ix8998 (.Y (nx8999), .A (nx7050)) ;
    buf02 ix9000 (.Y (nx9001), .A (nx7068)) ;
    buf02 ix9002 (.Y (nx9003), .A (nx7068)) ;
    buf02 ix9004 (.Y (nx9005), .A (nx7094)) ;
    buf02 ix9006 (.Y (nx9007), .A (nx7094)) ;
    buf02 ix9008 (.Y (nx9009), .A (nx7117)) ;
    buf02 ix9010 (.Y (nx9011), .A (nx7117)) ;
    inv02 ix9012 (.Y (nx9013), .A (nx3148)) ;
    buf02 ix9014 (.Y (nx9015), .A (nx7963)) ;
    buf02 ix9016 (.Y (nx9017), .A (nx7963)) ;
    buf02 ix9018 (.Y (nx9019), .A (nx8269)) ;
    buf02 ix9020 (.Y (nx9021), .A (nx8269)) ;
    inv02 ix9022 (.Y (nx9023), .A (nx5364)) ;
    buf02 ix9024 (.Y (nx9025), .A (nx8456)) ;
    buf02 ix9026 (.Y (nx9027), .A (nx8456)) ;
    buf02 ix9028 (.Y (nx9029), .A (nx8651)) ;
    buf02 ix9030 (.Y (nx9031), .A (nx8651)) ;
    nor02ii ix6957 (.Y (nx6956), .A0 (Address[1]), .A1 (Address[0])) ;
    nor02ii ix359 (.Y (nx358), .A0 (nx8989), .A1 (nx9067)) ;
    nor02ii ix373 (.Y (nx372), .A0 (nx8989), .A1 (nx9071)) ;
    nor02ii ix391 (.Y (nx390), .A0 (nx8989), .A1 (nx9075)) ;
    nor02ii ix51 (.Y (nx6966), .A0 (Address[0]), .A1 (Address[1])) ;
    nor02ii ix403 (.Y (nx402), .A0 (nx8989), .A1 (nx9049)) ;
    nor02ii ix275 (.Y (nx274), .A0 (nx7044), .A1 (nx9067)) ;
    nor02ii ix307 (.Y (nx306), .A0 (nx7044), .A1 (nx9075)) ;
    nor02ii ix319 (.Y (nx318), .A0 (nx7044), .A1 (nx9049)) ;
    nor02ii ix203 (.Y (nx202), .A0 (nx9001), .A1 (nx9067)) ;
    nor02ii ix217 (.Y (nx216), .A0 (nx9001), .A1 (nx9071)) ;
    nor02ii ix235 (.Y (nx234), .A0 (nx9001), .A1 (nx9075)) ;
    nor02ii ix247 (.Y (nx246), .A0 (nx9001), .A1 (nx9049)) ;
    nor02ii ix123 (.Y (nx122), .A0 (nx9005), .A1 (nx9067)) ;
    nor02ii ix137 (.Y (nx136), .A0 (nx9005), .A1 (nx9071)) ;
    nor02ii ix155 (.Y (nx154), .A0 (nx9005), .A1 (nx9075)) ;
    nor02ii ix167 (.Y (nx166), .A0 (nx9005), .A1 (nx9051)) ;
    nor02ii ix15 (.Y (nx14), .A0 (nx9009), .A1 (nx9067)) ;
    nor02ii ix33 (.Y (nx32), .A0 (nx9009), .A1 (nx9071)) ;
    nor02ii ix55 (.Y (nx54), .A0 (nx9009), .A1 (nx9077)) ;
    nor02ii ix69 (.Y (nx68), .A0 (nx9009), .A1 (nx9051)) ;
    and02 ix3189 (.Y (nx3188), .A0 (nx9079), .A1 (nx3148)) ;
    ao21 ix3143 (.Y (nx7941), .A0 (nx9069), .A1 (nx8971), .B0 (nx3122)) ;
    nor02ii ix3123 (.Y (nx3122), .A0 (nx9069), .A1 (Address[2])) ;
    or02 ix3131 (.Y (nx7945), .A0 (nx9069), .A1 (nx9051)) ;
    or02 ix7935 (.Y (nx7934), .A0 (nx9079), .A1 (nx9081)) ;
    and04 ix3363 (.Y (nx3362), .A0 (nx8817), .A1 (nx3148), .A2 (nx9053), .A3 (
          nx9081)) ;
    and04 ix3331 (.Y (nx3330), .A0 (nx6958), .A1 (nx9079), .A2 (nx7926), .A3 (
          nx3136)) ;
    nor02ii ix3137 (.Y (nx3136), .A0 (nx9053), .A1 (nx9083)) ;
    nor03_2x ix3249 (.Y (nx3248), .A0 (nx7968), .A1 (nx9079), .A2 (nx3148)) ;
    and03 ix3195 (.Y (nx3194), .A0 (nx3188), .A1 (nx9055), .A2 (nx9083)) ;
    and04 ix4831 (.Y (nx4830), .A0 (Address[3]), .A1 (Address[2]), .A2 (
          Address[1]), .A3 (nx8959)) ;
    and04 ix4807 (.Y (nx4806), .A0 (Address[1]), .A1 (nx8963), .A2 (Address[2])
          , .A3 (Address[4])) ;
    and04 ix4765 (.Y (nx4764), .A0 (nx8951), .A1 (Address[2]), .A2 (Address[3])
          , .A3 (Address[4])) ;
    and04 ix4743 (.Y (nx4742), .A0 (Address[1]), .A1 (Address[3]), .A2 (nx8971)
          , .A3 (Address[4])) ;
    and02 ix5347 (.Y (nx5346), .A0 (Address[2]), .A1 (nx9051)) ;
    nor02ii ix5435 (.Y (nx5434), .A0 (nx9057), .A1 (nx5364)) ;
    nor02ii ix5521 (.Y (nx5520), .A0 (nx8445), .A1 (nx5434)) ;
    and03 ix5527 (.Y (nx5526), .A0 (nx5406), .A1 (nx9057), .A2 (nx5364)) ;
    and02 ix5487 (.Y (nx5486), .A0 (nx9073), .A1 (nx3308)) ;
    or02 ix8464 (.Y (nx8463), .A0 (nx9057), .A1 (nx5364)) ;
    and03 ix5441 (.Y (nx5440), .A0 (nx5434), .A1 (nx9083), .A2 (nx5366)) ;
    and02 ix6099 (.Y (nx6098), .A0 (nx9069), .A1 (nx3308)) ;
    nor02ii ix6085 (.Y (nx6084), .A0 (nx6947), .A1 (Address[4])) ;
    and02 ix6059 (.Y (nx6058), .A0 (Address[1]), .A1 (nx3308)) ;
    nor02ii ix8752 (.Y (nx8753), .A0 (nx9009), .A1 (nx9069)) ;
    nor02ii ix8754 (.Y (nx8755), .A0 (nx9009), .A1 (nx9073)) ;
    nor02ii ix8756 (.Y (nx8757), .A0 (nx9009), .A1 (nx9077)) ;
    nor02ii ix8758 (.Y (nx8759), .A0 (nx9011), .A1 (nx9051)) ;
    nor02ii ix8766 (.Y (nx8767), .A0 (nx9005), .A1 (nx9069)) ;
    nor02ii ix8768 (.Y (nx8769), .A0 (nx9005), .A1 (nx9073)) ;
    nor02ii ix8770 (.Y (nx8771), .A0 (nx9005), .A1 (nx9077)) ;
    nor02ii ix8772 (.Y (nx8773), .A0 (nx9007), .A1 (nx9051)) ;
    nor02ii ix8774 (.Y (nx8775), .A0 (nx9001), .A1 (nx9069)) ;
    nor02ii ix8776 (.Y (nx8777), .A0 (nx9001), .A1 (nx9073)) ;
    nor02ii ix8778 (.Y (nx8779), .A0 (nx9001), .A1 (nx9077)) ;
    nor02ii ix8780 (.Y (nx8781), .A0 (nx9003), .A1 (nx9051)) ;
    nor02ii ix8782 (.Y (nx8783), .A0 (nx7044), .A1 (nx6944)) ;
    nor02ii ix8784 (.Y (nx8785), .A0 (nx7044), .A1 (nx9077)) ;
    nor02ii ix8786 (.Y (nx8787), .A0 (nx7044), .A1 (nx66)) ;
    nor02ii ix8792 (.Y (nx8793), .A0 (nx8989), .A1 (nx6944)) ;
    nor02ii ix8794 (.Y (nx8795), .A0 (nx8989), .A1 (nx9073)) ;
    nor02ii ix8796 (.Y (nx8797), .A0 (nx8989), .A1 (nx9077)) ;
    nor02ii ix8798 (.Y (nx8799), .A0 (nx8991), .A1 (nx66)) ;
    and02 ix8918 (.Y (nx8919), .A0 (nx9073), .A1 (nx3308)) ;
    and02 ix8936 (.Y (nx8937), .A0 (nx6944), .A1 (nx3308)) ;
    inv01 ix9048 (.Y (nx9049), .A (nx7033)) ;
    inv01 ix9050 (.Y (nx9051), .A (nx7033)) ;
    inv02 ix9052 (.Y (nx9053), .A (nx7955)) ;
    inv02 ix9054 (.Y (nx9055), .A (nx7955)) ;
    inv01 ix9056 (.Y (nx9057), .A (nx8437)) ;
    buf02 ix9058 (.Y (nx9059), .A (nx5520)) ;
    buf02 ix9060 (.Y (nx9061), .A (nx5520)) ;
    buf02 ix9062 (.Y (nx9063), .A (nx6084)) ;
    buf02 ix9064 (.Y (nx9065), .A (nx6084)) ;
    nor02_2x ix9066 (.Y (nx9067), .A0 (Address[1]), .A1 (Address[0])) ;
    nor02_2x ix9068 (.Y (nx9069), .A0 (Address[1]), .A1 (Address[0])) ;
    buf02 ix9070 (.Y (nx9071), .A (nx6956)) ;
    buf02 ix9072 (.Y (nx9073), .A (nx6956)) ;
    buf02 ix9074 (.Y (nx9075), .A (nx6966)) ;
    buf02 ix9076 (.Y (nx9077), .A (nx6966)) ;
    inv02 ix9078 (.Y (nx9079), .A (nx8817)) ;
    inv02 ix9080 (.Y (nx9081), .A (nx8813)) ;
    inv02 ix9082 (.Y (nx9083), .A (nx8813)) ;
    buf02 ix9084 (.Y (nx9085), .A (nx8753)) ;
    buf02 ix9086 (.Y (nx9087), .A (nx8755)) ;
    buf02 ix9088 (.Y (nx9089), .A (nx8757)) ;
    buf02 ix9090 (.Y (nx9091), .A (nx8759)) ;
    buf02 ix9092 (.Y (nx9093), .A (nx8767)) ;
    buf02 ix9094 (.Y (nx9095), .A (nx8769)) ;
    buf02 ix9096 (.Y (nx9097), .A (nx8771)) ;
    buf02 ix9098 (.Y (nx9099), .A (nx8773)) ;
    buf02 ix9100 (.Y (nx9101), .A (nx8775)) ;
    buf02 ix9102 (.Y (nx9103), .A (nx8777)) ;
    buf02 ix9104 (.Y (nx9105), .A (nx8779)) ;
    buf02 ix9106 (.Y (nx9107), .A (nx8781)) ;
    buf02 ix9108 (.Y (nx9109), .A (nx8783)) ;
    buf02 ix9110 (.Y (nx9111), .A (nx8785)) ;
    buf02 ix9112 (.Y (nx9113), .A (nx8787)) ;
    buf02 ix9114 (.Y (nx9115), .A (nx8793)) ;
    buf02 ix9116 (.Y (nx9117), .A (nx8795)) ;
    buf02 ix9118 (.Y (nx9119), .A (nx8797)) ;
    buf02 ix9120 (.Y (nx9121), .A (nx8799)) ;
    buf02 ix9122 (.Y (nx9123), .A (nx8919)) ;
    buf02 ix9124 (.Y (nx9125), .A (nx8937)) ;
endmodule

