//
// Verilog description for cell accelerator, 
// Wed May  9 07:36:06 2018
//
// LeonardoSpectrum Level 3, 2017a.2 
//


module accelerator ( CLK, RST, Start, FilterSize, Instr, FilterDin_0__0__7, 
                     FilterDin_0__0__6, FilterDin_0__0__5, FilterDin_0__0__4, 
                     FilterDin_0__0__3, FilterDin_0__0__2, FilterDin_0__0__1, 
                     FilterDin_0__0__0, FilterDin_0__1__7, FilterDin_0__1__6, 
                     FilterDin_0__1__5, FilterDin_0__1__4, FilterDin_0__1__3, 
                     FilterDin_0__1__2, FilterDin_0__1__1, FilterDin_0__1__0, 
                     FilterDin_0__2__7, FilterDin_0__2__6, FilterDin_0__2__5, 
                     FilterDin_0__2__4, FilterDin_0__2__3, FilterDin_0__2__2, 
                     FilterDin_0__2__1, FilterDin_0__2__0, FilterDin_0__3__7, 
                     FilterDin_0__3__6, FilterDin_0__3__5, FilterDin_0__3__4, 
                     FilterDin_0__3__3, FilterDin_0__3__2, FilterDin_0__3__1, 
                     FilterDin_0__3__0, FilterDin_0__4__7, FilterDin_0__4__6, 
                     FilterDin_0__4__5, FilterDin_0__4__4, FilterDin_0__4__3, 
                     FilterDin_0__4__2, FilterDin_0__4__1, FilterDin_0__4__0, 
                     FilterDin_1__0__7, FilterDin_1__0__6, FilterDin_1__0__5, 
                     FilterDin_1__0__4, FilterDin_1__0__3, FilterDin_1__0__2, 
                     FilterDin_1__0__1, FilterDin_1__0__0, FilterDin_1__1__7, 
                     FilterDin_1__1__6, FilterDin_1__1__5, FilterDin_1__1__4, 
                     FilterDin_1__1__3, FilterDin_1__1__2, FilterDin_1__1__1, 
                     FilterDin_1__1__0, FilterDin_1__2__7, FilterDin_1__2__6, 
                     FilterDin_1__2__5, FilterDin_1__2__4, FilterDin_1__2__3, 
                     FilterDin_1__2__2, FilterDin_1__2__1, FilterDin_1__2__0, 
                     FilterDin_1__3__7, FilterDin_1__3__6, FilterDin_1__3__5, 
                     FilterDin_1__3__4, FilterDin_1__3__3, FilterDin_1__3__2, 
                     FilterDin_1__3__1, FilterDin_1__3__0, FilterDin_1__4__7, 
                     FilterDin_1__4__6, FilterDin_1__4__5, FilterDin_1__4__4, 
                     FilterDin_1__4__3, FilterDin_1__4__2, FilterDin_1__4__1, 
                     FilterDin_1__4__0, FilterDin_2__0__7, FilterDin_2__0__6, 
                     FilterDin_2__0__5, FilterDin_2__0__4, FilterDin_2__0__3, 
                     FilterDin_2__0__2, FilterDin_2__0__1, FilterDin_2__0__0, 
                     FilterDin_2__1__7, FilterDin_2__1__6, FilterDin_2__1__5, 
                     FilterDin_2__1__4, FilterDin_2__1__3, FilterDin_2__1__2, 
                     FilterDin_2__1__1, FilterDin_2__1__0, FilterDin_2__2__7, 
                     FilterDin_2__2__6, FilterDin_2__2__5, FilterDin_2__2__4, 
                     FilterDin_2__2__3, FilterDin_2__2__2, FilterDin_2__2__1, 
                     FilterDin_2__2__0, FilterDin_2__3__7, FilterDin_2__3__6, 
                     FilterDin_2__3__5, FilterDin_2__3__4, FilterDin_2__3__3, 
                     FilterDin_2__3__2, FilterDin_2__3__1, FilterDin_2__3__0, 
                     FilterDin_2__4__7, FilterDin_2__4__6, FilterDin_2__4__5, 
                     FilterDin_2__4__4, FilterDin_2__4__3, FilterDin_2__4__2, 
                     FilterDin_2__4__1, FilterDin_2__4__0, FilterDin_3__0__7, 
                     FilterDin_3__0__6, FilterDin_3__0__5, FilterDin_3__0__4, 
                     FilterDin_3__0__3, FilterDin_3__0__2, FilterDin_3__0__1, 
                     FilterDin_3__0__0, FilterDin_3__1__7, FilterDin_3__1__6, 
                     FilterDin_3__1__5, FilterDin_3__1__4, FilterDin_3__1__3, 
                     FilterDin_3__1__2, FilterDin_3__1__1, FilterDin_3__1__0, 
                     FilterDin_3__2__7, FilterDin_3__2__6, FilterDin_3__2__5, 
                     FilterDin_3__2__4, FilterDin_3__2__3, FilterDin_3__2__2, 
                     FilterDin_3__2__1, FilterDin_3__2__0, FilterDin_3__3__7, 
                     FilterDin_3__3__6, FilterDin_3__3__5, FilterDin_3__3__4, 
                     FilterDin_3__3__3, FilterDin_3__3__2, FilterDin_3__3__1, 
                     FilterDin_3__3__0, FilterDin_3__4__7, FilterDin_3__4__6, 
                     FilterDin_3__4__5, FilterDin_3__4__4, FilterDin_3__4__3, 
                     FilterDin_3__4__2, FilterDin_3__4__1, FilterDin_3__4__0, 
                     FilterDin_4__0__7, FilterDin_4__0__6, FilterDin_4__0__5, 
                     FilterDin_4__0__4, FilterDin_4__0__3, FilterDin_4__0__2, 
                     FilterDin_4__0__1, FilterDin_4__0__0, FilterDin_4__1__7, 
                     FilterDin_4__1__6, FilterDin_4__1__5, FilterDin_4__1__4, 
                     FilterDin_4__1__3, FilterDin_4__1__2, FilterDin_4__1__1, 
                     FilterDin_4__1__0, FilterDin_4__2__7, FilterDin_4__2__6, 
                     FilterDin_4__2__5, FilterDin_4__2__4, FilterDin_4__2__3, 
                     FilterDin_4__2__2, FilterDin_4__2__1, FilterDin_4__2__0, 
                     FilterDin_4__3__7, FilterDin_4__3__6, FilterDin_4__3__5, 
                     FilterDin_4__3__4, FilterDin_4__3__3, FilterDin_4__3__2, 
                     FilterDin_4__3__1, FilterDin_4__3__0, FilterDin_4__4__7, 
                     FilterDin_4__4__6, FilterDin_4__4__5, FilterDin_4__4__4, 
                     FilterDin_4__4__3, FilterDin_4__4__2, FilterDin_4__4__1, 
                     FilterDin_4__4__0, WindowDin_0__0__7, WindowDin_0__0__6, 
                     WindowDin_0__0__5, WindowDin_0__0__4, WindowDin_0__0__3, 
                     WindowDin_0__0__2, WindowDin_0__0__1, WindowDin_0__0__0, 
                     WindowDin_0__1__7, WindowDin_0__1__6, WindowDin_0__1__5, 
                     WindowDin_0__1__4, WindowDin_0__1__3, WindowDin_0__1__2, 
                     WindowDin_0__1__1, WindowDin_0__1__0, WindowDin_0__2__7, 
                     WindowDin_0__2__6, WindowDin_0__2__5, WindowDin_0__2__4, 
                     WindowDin_0__2__3, WindowDin_0__2__2, WindowDin_0__2__1, 
                     WindowDin_0__2__0, WindowDin_0__3__7, WindowDin_0__3__6, 
                     WindowDin_0__3__5, WindowDin_0__3__4, WindowDin_0__3__3, 
                     WindowDin_0__3__2, WindowDin_0__3__1, WindowDin_0__3__0, 
                     WindowDin_0__4__7, WindowDin_0__4__6, WindowDin_0__4__5, 
                     WindowDin_0__4__4, WindowDin_0__4__3, WindowDin_0__4__2, 
                     WindowDin_0__4__1, WindowDin_0__4__0, WindowDin_1__0__7, 
                     WindowDin_1__0__6, WindowDin_1__0__5, WindowDin_1__0__4, 
                     WindowDin_1__0__3, WindowDin_1__0__2, WindowDin_1__0__1, 
                     WindowDin_1__0__0, WindowDin_1__1__7, WindowDin_1__1__6, 
                     WindowDin_1__1__5, WindowDin_1__1__4, WindowDin_1__1__3, 
                     WindowDin_1__1__2, WindowDin_1__1__1, WindowDin_1__1__0, 
                     WindowDin_1__2__7, WindowDin_1__2__6, WindowDin_1__2__5, 
                     WindowDin_1__2__4, WindowDin_1__2__3, WindowDin_1__2__2, 
                     WindowDin_1__2__1, WindowDin_1__2__0, WindowDin_1__3__7, 
                     WindowDin_1__3__6, WindowDin_1__3__5, WindowDin_1__3__4, 
                     WindowDin_1__3__3, WindowDin_1__3__2, WindowDin_1__3__1, 
                     WindowDin_1__3__0, WindowDin_1__4__7, WindowDin_1__4__6, 
                     WindowDin_1__4__5, WindowDin_1__4__4, WindowDin_1__4__3, 
                     WindowDin_1__4__2, WindowDin_1__4__1, WindowDin_1__4__0, 
                     WindowDin_2__0__7, WindowDin_2__0__6, WindowDin_2__0__5, 
                     WindowDin_2__0__4, WindowDin_2__0__3, WindowDin_2__0__2, 
                     WindowDin_2__0__1, WindowDin_2__0__0, WindowDin_2__1__7, 
                     WindowDin_2__1__6, WindowDin_2__1__5, WindowDin_2__1__4, 
                     WindowDin_2__1__3, WindowDin_2__1__2, WindowDin_2__1__1, 
                     WindowDin_2__1__0, WindowDin_2__2__7, WindowDin_2__2__6, 
                     WindowDin_2__2__5, WindowDin_2__2__4, WindowDin_2__2__3, 
                     WindowDin_2__2__2, WindowDin_2__2__1, WindowDin_2__2__0, 
                     WindowDin_2__3__7, WindowDin_2__3__6, WindowDin_2__3__5, 
                     WindowDin_2__3__4, WindowDin_2__3__3, WindowDin_2__3__2, 
                     WindowDin_2__3__1, WindowDin_2__3__0, WindowDin_2__4__7, 
                     WindowDin_2__4__6, WindowDin_2__4__5, WindowDin_2__4__4, 
                     WindowDin_2__4__3, WindowDin_2__4__2, WindowDin_2__4__1, 
                     WindowDin_2__4__0, WindowDin_3__0__7, WindowDin_3__0__6, 
                     WindowDin_3__0__5, WindowDin_3__0__4, WindowDin_3__0__3, 
                     WindowDin_3__0__2, WindowDin_3__0__1, WindowDin_3__0__0, 
                     WindowDin_3__1__7, WindowDin_3__1__6, WindowDin_3__1__5, 
                     WindowDin_3__1__4, WindowDin_3__1__3, WindowDin_3__1__2, 
                     WindowDin_3__1__1, WindowDin_3__1__0, WindowDin_3__2__7, 
                     WindowDin_3__2__6, WindowDin_3__2__5, WindowDin_3__2__4, 
                     WindowDin_3__2__3, WindowDin_3__2__2, WindowDin_3__2__1, 
                     WindowDin_3__2__0, WindowDin_3__3__7, WindowDin_3__3__6, 
                     WindowDin_3__3__5, WindowDin_3__3__4, WindowDin_3__3__3, 
                     WindowDin_3__3__2, WindowDin_3__3__1, WindowDin_3__3__0, 
                     WindowDin_3__4__7, WindowDin_3__4__6, WindowDin_3__4__5, 
                     WindowDin_3__4__4, WindowDin_3__4__3, WindowDin_3__4__2, 
                     WindowDin_3__4__1, WindowDin_3__4__0, WindowDin_4__0__7, 
                     WindowDin_4__0__6, WindowDin_4__0__5, WindowDin_4__0__4, 
                     WindowDin_4__0__3, WindowDin_4__0__2, WindowDin_4__0__1, 
                     WindowDin_4__0__0, WindowDin_4__1__7, WindowDin_4__1__6, 
                     WindowDin_4__1__5, WindowDin_4__1__4, WindowDin_4__1__3, 
                     WindowDin_4__1__2, WindowDin_4__1__1, WindowDin_4__1__0, 
                     WindowDin_4__2__7, WindowDin_4__2__6, WindowDin_4__2__5, 
                     WindowDin_4__2__4, WindowDin_4__2__3, WindowDin_4__2__2, 
                     WindowDin_4__2__1, WindowDin_4__2__0, WindowDin_4__3__7, 
                     WindowDin_4__3__6, WindowDin_4__3__5, WindowDin_4__3__4, 
                     WindowDin_4__3__3, WindowDin_4__3__2, WindowDin_4__3__1, 
                     WindowDin_4__3__0, WindowDin_4__4__7, WindowDin_4__4__6, 
                     WindowDin_4__4__5, WindowDin_4__4__4, WindowDin_4__4__3, 
                     WindowDin_4__4__2, WindowDin_4__4__1, WindowDin_4__4__0, 
                     Done, Result ) ;

    input CLK ;
    input RST ;
    input Start ;
    input FilterSize ;
    input Instr ;
    input FilterDin_0__0__7 ;
    input FilterDin_0__0__6 ;
    input FilterDin_0__0__5 ;
    input FilterDin_0__0__4 ;
    input FilterDin_0__0__3 ;
    input FilterDin_0__0__2 ;
    input FilterDin_0__0__1 ;
    input FilterDin_0__0__0 ;
    input FilterDin_0__1__7 ;
    input FilterDin_0__1__6 ;
    input FilterDin_0__1__5 ;
    input FilterDin_0__1__4 ;
    input FilterDin_0__1__3 ;
    input FilterDin_0__1__2 ;
    input FilterDin_0__1__1 ;
    input FilterDin_0__1__0 ;
    input FilterDin_0__2__7 ;
    input FilterDin_0__2__6 ;
    input FilterDin_0__2__5 ;
    input FilterDin_0__2__4 ;
    input FilterDin_0__2__3 ;
    input FilterDin_0__2__2 ;
    input FilterDin_0__2__1 ;
    input FilterDin_0__2__0 ;
    input FilterDin_0__3__7 ;
    input FilterDin_0__3__6 ;
    input FilterDin_0__3__5 ;
    input FilterDin_0__3__4 ;
    input FilterDin_0__3__3 ;
    input FilterDin_0__3__2 ;
    input FilterDin_0__3__1 ;
    input FilterDin_0__3__0 ;
    input FilterDin_0__4__7 ;
    input FilterDin_0__4__6 ;
    input FilterDin_0__4__5 ;
    input FilterDin_0__4__4 ;
    input FilterDin_0__4__3 ;
    input FilterDin_0__4__2 ;
    input FilterDin_0__4__1 ;
    input FilterDin_0__4__0 ;
    input FilterDin_1__0__7 ;
    input FilterDin_1__0__6 ;
    input FilterDin_1__0__5 ;
    input FilterDin_1__0__4 ;
    input FilterDin_1__0__3 ;
    input FilterDin_1__0__2 ;
    input FilterDin_1__0__1 ;
    input FilterDin_1__0__0 ;
    input FilterDin_1__1__7 ;
    input FilterDin_1__1__6 ;
    input FilterDin_1__1__5 ;
    input FilterDin_1__1__4 ;
    input FilterDin_1__1__3 ;
    input FilterDin_1__1__2 ;
    input FilterDin_1__1__1 ;
    input FilterDin_1__1__0 ;
    input FilterDin_1__2__7 ;
    input FilterDin_1__2__6 ;
    input FilterDin_1__2__5 ;
    input FilterDin_1__2__4 ;
    input FilterDin_1__2__3 ;
    input FilterDin_1__2__2 ;
    input FilterDin_1__2__1 ;
    input FilterDin_1__2__0 ;
    input FilterDin_1__3__7 ;
    input FilterDin_1__3__6 ;
    input FilterDin_1__3__5 ;
    input FilterDin_1__3__4 ;
    input FilterDin_1__3__3 ;
    input FilterDin_1__3__2 ;
    input FilterDin_1__3__1 ;
    input FilterDin_1__3__0 ;
    input FilterDin_1__4__7 ;
    input FilterDin_1__4__6 ;
    input FilterDin_1__4__5 ;
    input FilterDin_1__4__4 ;
    input FilterDin_1__4__3 ;
    input FilterDin_1__4__2 ;
    input FilterDin_1__4__1 ;
    input FilterDin_1__4__0 ;
    input FilterDin_2__0__7 ;
    input FilterDin_2__0__6 ;
    input FilterDin_2__0__5 ;
    input FilterDin_2__0__4 ;
    input FilterDin_2__0__3 ;
    input FilterDin_2__0__2 ;
    input FilterDin_2__0__1 ;
    input FilterDin_2__0__0 ;
    input FilterDin_2__1__7 ;
    input FilterDin_2__1__6 ;
    input FilterDin_2__1__5 ;
    input FilterDin_2__1__4 ;
    input FilterDin_2__1__3 ;
    input FilterDin_2__1__2 ;
    input FilterDin_2__1__1 ;
    input FilterDin_2__1__0 ;
    input FilterDin_2__2__7 ;
    input FilterDin_2__2__6 ;
    input FilterDin_2__2__5 ;
    input FilterDin_2__2__4 ;
    input FilterDin_2__2__3 ;
    input FilterDin_2__2__2 ;
    input FilterDin_2__2__1 ;
    input FilterDin_2__2__0 ;
    input FilterDin_2__3__7 ;
    input FilterDin_2__3__6 ;
    input FilterDin_2__3__5 ;
    input FilterDin_2__3__4 ;
    input FilterDin_2__3__3 ;
    input FilterDin_2__3__2 ;
    input FilterDin_2__3__1 ;
    input FilterDin_2__3__0 ;
    input FilterDin_2__4__7 ;
    input FilterDin_2__4__6 ;
    input FilterDin_2__4__5 ;
    input FilterDin_2__4__4 ;
    input FilterDin_2__4__3 ;
    input FilterDin_2__4__2 ;
    input FilterDin_2__4__1 ;
    input FilterDin_2__4__0 ;
    input FilterDin_3__0__7 ;
    input FilterDin_3__0__6 ;
    input FilterDin_3__0__5 ;
    input FilterDin_3__0__4 ;
    input FilterDin_3__0__3 ;
    input FilterDin_3__0__2 ;
    input FilterDin_3__0__1 ;
    input FilterDin_3__0__0 ;
    input FilterDin_3__1__7 ;
    input FilterDin_3__1__6 ;
    input FilterDin_3__1__5 ;
    input FilterDin_3__1__4 ;
    input FilterDin_3__1__3 ;
    input FilterDin_3__1__2 ;
    input FilterDin_3__1__1 ;
    input FilterDin_3__1__0 ;
    input FilterDin_3__2__7 ;
    input FilterDin_3__2__6 ;
    input FilterDin_3__2__5 ;
    input FilterDin_3__2__4 ;
    input FilterDin_3__2__3 ;
    input FilterDin_3__2__2 ;
    input FilterDin_3__2__1 ;
    input FilterDin_3__2__0 ;
    input FilterDin_3__3__7 ;
    input FilterDin_3__3__6 ;
    input FilterDin_3__3__5 ;
    input FilterDin_3__3__4 ;
    input FilterDin_3__3__3 ;
    input FilterDin_3__3__2 ;
    input FilterDin_3__3__1 ;
    input FilterDin_3__3__0 ;
    input FilterDin_3__4__7 ;
    input FilterDin_3__4__6 ;
    input FilterDin_3__4__5 ;
    input FilterDin_3__4__4 ;
    input FilterDin_3__4__3 ;
    input FilterDin_3__4__2 ;
    input FilterDin_3__4__1 ;
    input FilterDin_3__4__0 ;
    input FilterDin_4__0__7 ;
    input FilterDin_4__0__6 ;
    input FilterDin_4__0__5 ;
    input FilterDin_4__0__4 ;
    input FilterDin_4__0__3 ;
    input FilterDin_4__0__2 ;
    input FilterDin_4__0__1 ;
    input FilterDin_4__0__0 ;
    input FilterDin_4__1__7 ;
    input FilterDin_4__1__6 ;
    input FilterDin_4__1__5 ;
    input FilterDin_4__1__4 ;
    input FilterDin_4__1__3 ;
    input FilterDin_4__1__2 ;
    input FilterDin_4__1__1 ;
    input FilterDin_4__1__0 ;
    input FilterDin_4__2__7 ;
    input FilterDin_4__2__6 ;
    input FilterDin_4__2__5 ;
    input FilterDin_4__2__4 ;
    input FilterDin_4__2__3 ;
    input FilterDin_4__2__2 ;
    input FilterDin_4__2__1 ;
    input FilterDin_4__2__0 ;
    input FilterDin_4__3__7 ;
    input FilterDin_4__3__6 ;
    input FilterDin_4__3__5 ;
    input FilterDin_4__3__4 ;
    input FilterDin_4__3__3 ;
    input FilterDin_4__3__2 ;
    input FilterDin_4__3__1 ;
    input FilterDin_4__3__0 ;
    input FilterDin_4__4__7 ;
    input FilterDin_4__4__6 ;
    input FilterDin_4__4__5 ;
    input FilterDin_4__4__4 ;
    input FilterDin_4__4__3 ;
    input FilterDin_4__4__2 ;
    input FilterDin_4__4__1 ;
    input FilterDin_4__4__0 ;
    input WindowDin_0__0__7 ;
    input WindowDin_0__0__6 ;
    input WindowDin_0__0__5 ;
    input WindowDin_0__0__4 ;
    input WindowDin_0__0__3 ;
    input WindowDin_0__0__2 ;
    input WindowDin_0__0__1 ;
    input WindowDin_0__0__0 ;
    input WindowDin_0__1__7 ;
    input WindowDin_0__1__6 ;
    input WindowDin_0__1__5 ;
    input WindowDin_0__1__4 ;
    input WindowDin_0__1__3 ;
    input WindowDin_0__1__2 ;
    input WindowDin_0__1__1 ;
    input WindowDin_0__1__0 ;
    input WindowDin_0__2__7 ;
    input WindowDin_0__2__6 ;
    input WindowDin_0__2__5 ;
    input WindowDin_0__2__4 ;
    input WindowDin_0__2__3 ;
    input WindowDin_0__2__2 ;
    input WindowDin_0__2__1 ;
    input WindowDin_0__2__0 ;
    input WindowDin_0__3__7 ;
    input WindowDin_0__3__6 ;
    input WindowDin_0__3__5 ;
    input WindowDin_0__3__4 ;
    input WindowDin_0__3__3 ;
    input WindowDin_0__3__2 ;
    input WindowDin_0__3__1 ;
    input WindowDin_0__3__0 ;
    input WindowDin_0__4__7 ;
    input WindowDin_0__4__6 ;
    input WindowDin_0__4__5 ;
    input WindowDin_0__4__4 ;
    input WindowDin_0__4__3 ;
    input WindowDin_0__4__2 ;
    input WindowDin_0__4__1 ;
    input WindowDin_0__4__0 ;
    input WindowDin_1__0__7 ;
    input WindowDin_1__0__6 ;
    input WindowDin_1__0__5 ;
    input WindowDin_1__0__4 ;
    input WindowDin_1__0__3 ;
    input WindowDin_1__0__2 ;
    input WindowDin_1__0__1 ;
    input WindowDin_1__0__0 ;
    input WindowDin_1__1__7 ;
    input WindowDin_1__1__6 ;
    input WindowDin_1__1__5 ;
    input WindowDin_1__1__4 ;
    input WindowDin_1__1__3 ;
    input WindowDin_1__1__2 ;
    input WindowDin_1__1__1 ;
    input WindowDin_1__1__0 ;
    input WindowDin_1__2__7 ;
    input WindowDin_1__2__6 ;
    input WindowDin_1__2__5 ;
    input WindowDin_1__2__4 ;
    input WindowDin_1__2__3 ;
    input WindowDin_1__2__2 ;
    input WindowDin_1__2__1 ;
    input WindowDin_1__2__0 ;
    input WindowDin_1__3__7 ;
    input WindowDin_1__3__6 ;
    input WindowDin_1__3__5 ;
    input WindowDin_1__3__4 ;
    input WindowDin_1__3__3 ;
    input WindowDin_1__3__2 ;
    input WindowDin_1__3__1 ;
    input WindowDin_1__3__0 ;
    input WindowDin_1__4__7 ;
    input WindowDin_1__4__6 ;
    input WindowDin_1__4__5 ;
    input WindowDin_1__4__4 ;
    input WindowDin_1__4__3 ;
    input WindowDin_1__4__2 ;
    input WindowDin_1__4__1 ;
    input WindowDin_1__4__0 ;
    input WindowDin_2__0__7 ;
    input WindowDin_2__0__6 ;
    input WindowDin_2__0__5 ;
    input WindowDin_2__0__4 ;
    input WindowDin_2__0__3 ;
    input WindowDin_2__0__2 ;
    input WindowDin_2__0__1 ;
    input WindowDin_2__0__0 ;
    input WindowDin_2__1__7 ;
    input WindowDin_2__1__6 ;
    input WindowDin_2__1__5 ;
    input WindowDin_2__1__4 ;
    input WindowDin_2__1__3 ;
    input WindowDin_2__1__2 ;
    input WindowDin_2__1__1 ;
    input WindowDin_2__1__0 ;
    input WindowDin_2__2__7 ;
    input WindowDin_2__2__6 ;
    input WindowDin_2__2__5 ;
    input WindowDin_2__2__4 ;
    input WindowDin_2__2__3 ;
    input WindowDin_2__2__2 ;
    input WindowDin_2__2__1 ;
    input WindowDin_2__2__0 ;
    input WindowDin_2__3__7 ;
    input WindowDin_2__3__6 ;
    input WindowDin_2__3__5 ;
    input WindowDin_2__3__4 ;
    input WindowDin_2__3__3 ;
    input WindowDin_2__3__2 ;
    input WindowDin_2__3__1 ;
    input WindowDin_2__3__0 ;
    input WindowDin_2__4__7 ;
    input WindowDin_2__4__6 ;
    input WindowDin_2__4__5 ;
    input WindowDin_2__4__4 ;
    input WindowDin_2__4__3 ;
    input WindowDin_2__4__2 ;
    input WindowDin_2__4__1 ;
    input WindowDin_2__4__0 ;
    input WindowDin_3__0__7 ;
    input WindowDin_3__0__6 ;
    input WindowDin_3__0__5 ;
    input WindowDin_3__0__4 ;
    input WindowDin_3__0__3 ;
    input WindowDin_3__0__2 ;
    input WindowDin_3__0__1 ;
    input WindowDin_3__0__0 ;
    input WindowDin_3__1__7 ;
    input WindowDin_3__1__6 ;
    input WindowDin_3__1__5 ;
    input WindowDin_3__1__4 ;
    input WindowDin_3__1__3 ;
    input WindowDin_3__1__2 ;
    input WindowDin_3__1__1 ;
    input WindowDin_3__1__0 ;
    input WindowDin_3__2__7 ;
    input WindowDin_3__2__6 ;
    input WindowDin_3__2__5 ;
    input WindowDin_3__2__4 ;
    input WindowDin_3__2__3 ;
    input WindowDin_3__2__2 ;
    input WindowDin_3__2__1 ;
    input WindowDin_3__2__0 ;
    input WindowDin_3__3__7 ;
    input WindowDin_3__3__6 ;
    input WindowDin_3__3__5 ;
    input WindowDin_3__3__4 ;
    input WindowDin_3__3__3 ;
    input WindowDin_3__3__2 ;
    input WindowDin_3__3__1 ;
    input WindowDin_3__3__0 ;
    input WindowDin_3__4__7 ;
    input WindowDin_3__4__6 ;
    input WindowDin_3__4__5 ;
    input WindowDin_3__4__4 ;
    input WindowDin_3__4__3 ;
    input WindowDin_3__4__2 ;
    input WindowDin_3__4__1 ;
    input WindowDin_3__4__0 ;
    input WindowDin_4__0__7 ;
    input WindowDin_4__0__6 ;
    input WindowDin_4__0__5 ;
    input WindowDin_4__0__4 ;
    input WindowDin_4__0__3 ;
    input WindowDin_4__0__2 ;
    input WindowDin_4__0__1 ;
    input WindowDin_4__0__0 ;
    input WindowDin_4__1__7 ;
    input WindowDin_4__1__6 ;
    input WindowDin_4__1__5 ;
    input WindowDin_4__1__4 ;
    input WindowDin_4__1__3 ;
    input WindowDin_4__1__2 ;
    input WindowDin_4__1__1 ;
    input WindowDin_4__1__0 ;
    input WindowDin_4__2__7 ;
    input WindowDin_4__2__6 ;
    input WindowDin_4__2__5 ;
    input WindowDin_4__2__4 ;
    input WindowDin_4__2__3 ;
    input WindowDin_4__2__2 ;
    input WindowDin_4__2__1 ;
    input WindowDin_4__2__0 ;
    input WindowDin_4__3__7 ;
    input WindowDin_4__3__6 ;
    input WindowDin_4__3__5 ;
    input WindowDin_4__3__4 ;
    input WindowDin_4__3__3 ;
    input WindowDin_4__3__2 ;
    input WindowDin_4__3__1 ;
    input WindowDin_4__3__0 ;
    input WindowDin_4__4__7 ;
    input WindowDin_4__4__6 ;
    input WindowDin_4__4__5 ;
    input WindowDin_4__4__4 ;
    input WindowDin_4__4__3 ;
    input WindowDin_4__4__2 ;
    input WindowDin_4__4__1 ;
    input WindowDin_4__4__0 ;
    output Done ;
    output [7:0]Result ;

    wire LoopingAndResultNotReady, L1FirstOperands_0__15, L1FirstOperands_0__14, 
         L1FirstOperands_0__13, L1FirstOperands_0__12, L1FirstOperands_0__11, 
         L1FirstOperands_0__10, L1FirstOperands_0__9, L1FirstOperands_0__8, 
         L1FirstOperands_0__7, L1FirstOperands_0__6, L1FirstOperands_0__5, 
         L1FirstOperands_0__4, L1FirstOperands_0__3, L1FirstOperands_0__2, 
         L1FirstOperands_0__1, L1FirstOperands_0__0, L1FirstOperands_2__15, 
         L1FirstOperands_2__14, L1FirstOperands_2__13, L1FirstOperands_2__12, 
         L1FirstOperands_2__11, L1FirstOperands_2__10, L1FirstOperands_2__9, 
         L1FirstOperands_2__8, L1FirstOperands_2__7, L1FirstOperands_2__6, 
         L1FirstOperands_2__5, L1FirstOperands_2__4, L1FirstOperands_2__3, 
         L1FirstOperands_2__2, L1FirstOperands_2__1, L1FirstOperands_2__0, 
         L1FirstOperands_3__15, L1FirstOperands_3__14, L1FirstOperands_3__13, 
         L1FirstOperands_3__12, L1FirstOperands_3__11, L1FirstOperands_3__10, 
         L1FirstOperands_3__9, L1FirstOperands_3__8, L1FirstOperands_3__7, 
         L1FirstOperands_3__6, L1FirstOperands_3__5, L1FirstOperands_3__4, 
         L1FirstOperands_3__3, L1FirstOperands_3__2, L1FirstOperands_3__1, 
         L1FirstOperands_3__0, L1FirstOperands_4__15, L1FirstOperands_4__14, 
         L1FirstOperands_4__13, L1FirstOperands_4__12, L1FirstOperands_4__11, 
         L1FirstOperands_4__10, L1FirstOperands_4__9, L1FirstOperands_4__8, 
         L1FirstOperands_4__7, L1FirstOperands_4__6, L1FirstOperands_4__5, 
         L1FirstOperands_4__4, L1FirstOperands_4__3, L1FirstOperands_4__2, 
         L1FirstOperands_4__1, L1FirstOperands_4__0, L1FirstOperands_6__15, 
         L1FirstOperands_6__14, L1FirstOperands_6__13, L1FirstOperands_6__12, 
         L1FirstOperands_6__11, L1FirstOperands_6__10, L1FirstOperands_6__9, 
         L1FirstOperands_6__8, L1FirstOperands_6__7, L1FirstOperands_6__6, 
         L1FirstOperands_6__5, L1FirstOperands_6__4, L1FirstOperands_6__3, 
         L1FirstOperands_6__2, L1FirstOperands_6__1, L1FirstOperands_6__0, 
         L1FirstOperands_7__15, L1FirstOperands_7__14, L1FirstOperands_7__13, 
         L1FirstOperands_7__12, L1FirstOperands_7__11, L1FirstOperands_7__10, 
         L1FirstOperands_7__9, L1FirstOperands_7__8, L1FirstOperands_7__7, 
         L1FirstOperands_7__6, L1FirstOperands_7__5, L1FirstOperands_7__4, 
         L1FirstOperands_7__3, L1FirstOperands_7__2, L1FirstOperands_7__1, 
         L1FirstOperands_7__0, L1FirstOperands_8__15, L1FirstOperands_8__14, 
         L1FirstOperands_8__13, L1FirstOperands_8__12, L1FirstOperands_8__11, 
         L1FirstOperands_8__10, L1FirstOperands_8__9, L1FirstOperands_8__8, 
         L1FirstOperands_8__7, L1FirstOperands_8__6, L1FirstOperands_8__5, 
         L1FirstOperands_8__4, L1FirstOperands_8__3, L1FirstOperands_8__2, 
         L1FirstOperands_8__1, L1FirstOperands_8__0, L1FirstOperands_10__15, 
         L1FirstOperands_10__14, L1FirstOperands_10__13, L1FirstOperands_10__12, 
         L1FirstOperands_10__11, L1FirstOperands_10__10, L1FirstOperands_10__9, 
         L1FirstOperands_10__8, L1FirstOperands_10__7, L1FirstOperands_10__6, 
         L1FirstOperands_10__5, L1FirstOperands_10__4, L1FirstOperands_10__3, 
         L1FirstOperands_10__2, L1FirstOperands_10__1, L1FirstOperands_10__0, 
         L1FirstOperands_11__15, L1FirstOperands_11__14, L1FirstOperands_11__13, 
         L1FirstOperands_11__12, L1FirstOperands_11__11, L1FirstOperands_11__10, 
         L1FirstOperands_11__9, L1FirstOperands_11__8, L1FirstOperands_11__7, 
         L1FirstOperands_11__6, L1FirstOperands_11__5, L1FirstOperands_11__4, 
         L1FirstOperands_11__3, L1FirstOperands_11__2, L1FirstOperands_11__1, 
         L1FirstOperands_11__0, L1ResultsLarge_0__16, L1ResultsLarge_0__15, 
         L1ResultsLarge_0__14, L1ResultsLarge_0__13, L1ResultsLarge_0__12, 
         L1ResultsLarge_0__11, L1ResultsLarge_0__10, L1ResultsLarge_0__9, 
         L1ResultsLarge_0__8, L1ResultsLarge_0__7, L1ResultsLarge_0__6, 
         L1ResultsLarge_0__5, L1ResultsLarge_0__4, L1ResultsLarge_0__3, 
         L1ResultsLarge_0__2, L1ResultsLarge_0__1, L1ResultsLarge_0__0, 
         L1ResultsLarge_1__16, L1ResultsLarge_1__15, L1ResultsLarge_1__14, 
         L1ResultsLarge_1__13, L1ResultsLarge_1__12, L1ResultsLarge_1__11, 
         L1ResultsLarge_1__10, L1ResultsLarge_1__9, L1ResultsLarge_1__8, 
         L1ResultsLarge_1__7, L1ResultsLarge_1__6, L1ResultsLarge_1__5, 
         L1ResultsLarge_1__4, L1ResultsLarge_1__3, L1ResultsLarge_1__2, 
         L1ResultsLarge_1__1, L1ResultsLarge_1__0, L1ResultsLarge_2__16, 
         L1ResultsLarge_2__15, L1ResultsLarge_2__14, L1ResultsLarge_2__13, 
         L1ResultsLarge_2__12, L1ResultsLarge_2__11, L1ResultsLarge_2__10, 
         L1ResultsLarge_2__9, L1ResultsLarge_2__8, L1ResultsLarge_2__7, 
         L1ResultsLarge_2__6, L1ResultsLarge_2__5, L1ResultsLarge_2__4, 
         L1ResultsLarge_2__3, L1ResultsLarge_2__2, L1ResultsLarge_2__1, 
         L1ResultsLarge_2__0, L1ResultsLarge_3__16, L1ResultsLarge_3__15, 
         L1ResultsLarge_3__14, L1ResultsLarge_3__13, L1ResultsLarge_3__12, 
         L1ResultsLarge_3__11, L1ResultsLarge_3__10, L1ResultsLarge_3__9, 
         L1ResultsLarge_3__8, L1ResultsLarge_3__7, L1ResultsLarge_3__6, 
         L1ResultsLarge_3__5, L1ResultsLarge_3__4, L1ResultsLarge_3__3, 
         L1ResultsLarge_3__2, L1ResultsLarge_3__1, L1ResultsLarge_3__0, 
         L1ResultsLarge_4__16, L1ResultsLarge_4__15, L1ResultsLarge_4__14, 
         L1ResultsLarge_4__13, L1ResultsLarge_4__12, L1ResultsLarge_4__11, 
         L1ResultsLarge_4__10, L1ResultsLarge_4__9, L1ResultsLarge_4__8, 
         L1ResultsLarge_4__7, L1ResultsLarge_4__6, L1ResultsLarge_4__5, 
         L1ResultsLarge_4__4, L1ResultsLarge_4__3, L1ResultsLarge_4__2, 
         L1ResultsLarge_4__1, L1ResultsLarge_4__0, L1ResultsLarge_5__16, 
         L1ResultsLarge_5__15, L1ResultsLarge_5__14, L1ResultsLarge_5__13, 
         L1ResultsLarge_5__12, L1ResultsLarge_5__11, L1ResultsLarge_5__10, 
         L1ResultsLarge_5__9, L1ResultsLarge_5__8, L1ResultsLarge_5__7, 
         L1ResultsLarge_5__6, L1ResultsLarge_5__5, L1ResultsLarge_5__4, 
         L1ResultsLarge_5__3, L1ResultsLarge_5__2, L1ResultsLarge_5__1, 
         L1ResultsLarge_5__0, L1ResultsLarge_6__16, L1ResultsLarge_6__15, 
         L1ResultsLarge_6__14, L1ResultsLarge_6__13, L1ResultsLarge_6__12, 
         L1ResultsLarge_6__11, L1ResultsLarge_6__10, L1ResultsLarge_6__9, 
         L1ResultsLarge_6__8, L1ResultsLarge_6__7, L1ResultsLarge_6__6, 
         L1ResultsLarge_6__5, L1ResultsLarge_6__4, L1ResultsLarge_6__3, 
         L1ResultsLarge_6__2, L1ResultsLarge_6__1, L1ResultsLarge_6__0, 
         L1ResultsLarge_7__16, L1ResultsLarge_7__15, L1ResultsLarge_7__14, 
         L1ResultsLarge_7__13, L1ResultsLarge_7__12, L1ResultsLarge_7__11, 
         L1ResultsLarge_7__10, L1ResultsLarge_7__9, L1ResultsLarge_7__8, 
         L1ResultsLarge_7__7, L1ResultsLarge_7__6, L1ResultsLarge_7__5, 
         L1ResultsLarge_7__4, L1ResultsLarge_7__3, L1ResultsLarge_7__2, 
         L1ResultsLarge_7__1, L1ResultsLarge_7__0, L1ResultsLarge_8__16, 
         L1ResultsLarge_8__15, L1ResultsLarge_8__14, L1ResultsLarge_8__13, 
         L1ResultsLarge_8__12, L1ResultsLarge_8__11, L1ResultsLarge_8__10, 
         L1ResultsLarge_8__9, L1ResultsLarge_8__8, L1ResultsLarge_8__7, 
         L1ResultsLarge_8__6, L1ResultsLarge_8__5, L1ResultsLarge_8__4, 
         L1ResultsLarge_8__3, L1ResultsLarge_8__2, L1ResultsLarge_8__1, 
         L1ResultsLarge_8__0, L1ResultsLarge_9__16, L1ResultsLarge_9__15, 
         L1ResultsLarge_9__14, L1ResultsLarge_9__13, L1ResultsLarge_9__12, 
         L1ResultsLarge_9__11, L1ResultsLarge_9__10, L1ResultsLarge_9__9, 
         L1ResultsLarge_9__8, L1ResultsLarge_9__7, L1ResultsLarge_9__6, 
         L1ResultsLarge_9__5, L1ResultsLarge_9__4, L1ResultsLarge_9__3, 
         L1ResultsLarge_9__2, L1ResultsLarge_9__1, L1ResultsLarge_9__0, 
         L1ResultsLarge_10__16, L1ResultsLarge_10__15, L1ResultsLarge_10__14, 
         L1ResultsLarge_10__13, L1ResultsLarge_10__12, L1ResultsLarge_10__11, 
         L1ResultsLarge_10__10, L1ResultsLarge_10__9, L1ResultsLarge_10__8, 
         L1ResultsLarge_10__7, L1ResultsLarge_10__6, L1ResultsLarge_10__5, 
         L1ResultsLarge_10__4, L1ResultsLarge_10__3, L1ResultsLarge_10__2, 
         L1ResultsLarge_10__1, L1ResultsLarge_10__0, L1ResultsLarge_11__16, 
         L1ResultsLarge_11__15, L1ResultsLarge_11__14, L1ResultsLarge_11__13, 
         L1ResultsLarge_11__12, L1ResultsLarge_11__11, L1ResultsLarge_11__10, 
         L1ResultsLarge_11__9, L1ResultsLarge_11__8, L1ResultsLarge_11__7, 
         L1ResultsLarge_11__6, L1ResultsLarge_11__5, L1ResultsLarge_11__4, 
         L1ResultsLarge_11__3, L1ResultsLarge_11__2, L1ResultsLarge_11__1, 
         L1ResultsLarge_11__0, L2ResultsLarge_0__16, L2ResultsLarge_0__15, 
         L2ResultsLarge_0__14, L2ResultsLarge_0__13, L2ResultsLarge_0__12, 
         L2ResultsLarge_0__11, L2ResultsLarge_0__10, L2ResultsLarge_0__9, 
         L2ResultsLarge_0__8, L2ResultsLarge_0__7, L2ResultsLarge_0__6, 
         L2ResultsLarge_0__5, L2ResultsLarge_0__4, L2ResultsLarge_0__3, 
         L2ResultsLarge_0__2, L2ResultsLarge_0__1, L2ResultsLarge_0__0, 
         L2ResultsLarge_1__16, L2ResultsLarge_1__15, L2ResultsLarge_1__14, 
         L2ResultsLarge_1__13, L2ResultsLarge_1__12, L2ResultsLarge_1__11, 
         L2ResultsLarge_1__10, L2ResultsLarge_1__9, L2ResultsLarge_1__8, 
         L2ResultsLarge_1__7, L2ResultsLarge_1__6, L2ResultsLarge_1__5, 
         L2ResultsLarge_1__4, L2ResultsLarge_1__3, L2ResultsLarge_1__2, 
         L2ResultsLarge_1__1, L2ResultsLarge_1__0, L2ResultsLarge_2__16, 
         L2ResultsLarge_2__15, L2ResultsLarge_2__14, L2ResultsLarge_2__13, 
         L2ResultsLarge_2__12, L2ResultsLarge_2__11, L2ResultsLarge_2__10, 
         L2ResultsLarge_2__9, L2ResultsLarge_2__8, L2ResultsLarge_2__7, 
         L2ResultsLarge_2__6, L2ResultsLarge_2__5, L2ResultsLarge_2__4, 
         L2ResultsLarge_2__3, L2ResultsLarge_2__2, L2ResultsLarge_2__1, 
         L2ResultsLarge_2__0, L2ResultsLarge_3__16, L2ResultsLarge_3__15, 
         L2ResultsLarge_3__14, L2ResultsLarge_3__13, L2ResultsLarge_3__12, 
         L2ResultsLarge_3__11, L2ResultsLarge_3__10, L2ResultsLarge_3__9, 
         L2ResultsLarge_3__8, L2ResultsLarge_3__7, L2ResultsLarge_3__6, 
         L2ResultsLarge_3__5, L2ResultsLarge_3__4, L2ResultsLarge_3__3, 
         L2ResultsLarge_3__2, L2ResultsLarge_3__1, L2ResultsLarge_3__0, 
         L2ResultsLarge_4__16, L2ResultsLarge_4__15, L2ResultsLarge_4__14, 
         L2ResultsLarge_4__13, L2ResultsLarge_4__12, L2ResultsLarge_4__11, 
         L2ResultsLarge_4__10, L2ResultsLarge_4__9, L2ResultsLarge_4__8, 
         L2ResultsLarge_4__7, L2ResultsLarge_4__6, L2ResultsLarge_4__5, 
         L2ResultsLarge_4__4, L2ResultsLarge_4__3, L2ResultsLarge_4__2, 
         L2ResultsLarge_4__1, L2ResultsLarge_4__0, L2ResultsLarge_5__16, 
         L2ResultsLarge_5__15, L2ResultsLarge_5__14, L2ResultsLarge_5__13, 
         L2ResultsLarge_5__12, L2ResultsLarge_5__11, L2ResultsLarge_5__10, 
         L2ResultsLarge_5__9, L2ResultsLarge_5__8, L2ResultsLarge_5__7, 
         L2ResultsLarge_5__6, L2ResultsLarge_5__5, L2ResultsLarge_5__4, 
         L2ResultsLarge_5__3, L2ResultsLarge_5__2, L2ResultsLarge_5__1, 
         L2ResultsLarge_5__0, L3ResultsLarge_0__16, L3ResultsLarge_0__15, 
         L3ResultsLarge_0__14, L3ResultsLarge_0__13, L3ResultsLarge_0__12, 
         L3ResultsLarge_0__11, L3ResultsLarge_0__10, L3ResultsLarge_0__9, 
         L3ResultsLarge_0__8, L3ResultsLarge_0__7, L3ResultsLarge_0__6, 
         L3ResultsLarge_0__5, L3ResultsLarge_0__4, L3ResultsLarge_0__3, 
         L3ResultsLarge_0__2, L3ResultsLarge_0__1, L3ResultsLarge_0__0, 
         L3ResultsLarge_1__16, L3ResultsLarge_1__15, L3ResultsLarge_1__14, 
         L3ResultsLarge_1__13, L3ResultsLarge_1__12, L3ResultsLarge_1__11, 
         L3ResultsLarge_1__10, L3ResultsLarge_1__9, L3ResultsLarge_1__8, 
         L3ResultsLarge_1__7, L3ResultsLarge_1__6, L3ResultsLarge_1__5, 
         L3ResultsLarge_1__4, L3ResultsLarge_1__3, L3ResultsLarge_1__2, 
         L3ResultsLarge_1__1, L3ResultsLarge_1__0, L3ResultsLarge_2__16, 
         L3ResultsLarge_2__15, L3ResultsLarge_2__14, L3ResultsLarge_2__13, 
         L3ResultsLarge_2__12, L3ResultsLarge_2__11, L3ResultsLarge_2__10, 
         L3ResultsLarge_2__9, L3ResultsLarge_2__8, L3ResultsLarge_2__7, 
         L3ResultsLarge_2__6, L3ResultsLarge_2__5, L3ResultsLarge_2__4, 
         L3ResultsLarge_2__3, L3ResultsLarge_2__2, L3ResultsLarge_2__1, 
         L3ResultsLarge_2__0, L4ResultsLarge_0__16, L4ResultsLarge_0__15, 
         L4ResultsLarge_0__14, L4ResultsLarge_0__13, L4ResultsLarge_0__12, 
         L4ResultsLarge_0__11, L4ResultsLarge_0__10, L4ResultsLarge_0__9, 
         L4ResultsLarge_0__8, L4ResultsLarge_0__7, L4ResultsLarge_0__6, 
         L4ResultsLarge_0__5, L4ResultsLarge_0__4, L4ResultsLarge_0__3, 
         L4ResultsLarge_0__2, L4ResultsLarge_0__1, L4ResultsLarge_0__0, 
         L5FirstOperands_1__16, L5FirstOperands_1__15, L5FirstOperands_1__14, 
         L5FirstOperands_1__13, L5FirstOperands_1__12, L5FirstOperands_1__11, 
         L5FirstOperands_1__10, L5FirstOperands_1__9, L5FirstOperands_1__8, 
         L5FirstOperands_1__7, L5FirstOperands_1__6, L5FirstOperands_1__5, 
         L5FirstOperands_1__4, L5FirstOperands_1__3, L5FirstOperands_1__2, 
         L5FirstOperands_1__1, L5FirstOperands_1__0, 
         L1_0_L2_0_G1_MINI_ALU_OperationResult_15, 
         L1_0_L2_0_G1_MINI_ALU_OperationResult_14, 
         L1_0_L2_0_G1_MINI_ALU_OperationResult_13, 
         L1_0_L2_0_G1_MINI_ALU_OperationResult_12, 
         L1_0_L2_0_G1_MINI_ALU_OperationResult_11, 
         L1_0_L2_0_G1_MINI_ALU_OperationResult_10, 
         L1_0_L2_0_G1_MINI_ALU_OperationResult_9, 
         L1_0_L2_0_G1_MINI_ALU_OperationResult_8, 
         L1_0_L2_0_G1_MINI_ALU_OperationResult_7, 
         L1_0_L2_0_G1_MINI_ALU_OperationResult_6, 
         L1_0_L2_0_G1_MINI_ALU_OperationResult_5, 
         L1_0_L2_0_G1_MINI_ALU_OperationResult_4, 
         L1_0_L2_0_G1_MINI_ALU_OperationResult_3, 
         L1_0_L2_0_G1_MINI_ALU_OperationResult_2, 
         L1_0_L2_0_G1_MINI_ALU_OperationResult_1, 
         L1_0_L2_0_G1_MINI_ALU_OperationResult_0, 
         L1_0_L2_0_G1_MINI_ALU_BoothXORCheck, 
         L1_0_L2_0_G1_MINI_ALU_BoothOperand_16, 
         L1_0_L2_0_G1_MINI_ALU_BoothOperand_15, 
         L1_0_L2_0_G1_MINI_ALU_BoothOperand_14, 
         L1_0_L2_0_G1_MINI_ALU_BoothOperand_13, 
         L1_0_L2_0_G1_MINI_ALU_BoothOperand_12, 
         L1_0_L2_0_G1_MINI_ALU_BoothOperand_11, 
         L1_0_L2_0_G1_MINI_ALU_BoothOperand_10, 
         L1_0_L2_0_G1_MINI_ALU_BoothOperand_9, L1_0_L2_0_G1_MINI_ALU_BoothP_16, 
         L1_0_L2_0_G1_MINI_ALU_BoothP_15, L1_0_L2_0_G1_MINI_ALU_BoothP_14, 
         L1_0_L2_0_G1_MINI_ALU_BoothP_13, L1_0_L2_0_G1_MINI_ALU_BoothP_12, 
         L1_0_L2_0_G1_MINI_ALU_BoothP_11, L1_0_L2_0_G1_MINI_ALU_BoothP_10, 
         L1_0_L2_0_G1_MINI_ALU_BoothP_9, L1_0_L2_0_G1_MINI_ALU_BoothP_8, 
         L1_0_L2_0_G1_MINI_ALU_BoothP_7, L1_0_L2_0_G1_MINI_ALU_BoothP_6, 
         L1_0_L2_0_G1_MINI_ALU_BoothP_5, L1_0_L2_0_G1_MINI_ALU_BoothP_4, 
         L1_0_L2_0_G1_MINI_ALU_BoothP_3, L1_0_L2_0_G1_MINI_ALU_BoothP_2, 
         L1_0_L2_0_G1_MINI_ALU_BoothP_1, L1_0_L2_0_G1_MINI_ALU_BoothP_0, 
         L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_15, 
         L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_14, 
         L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_13, 
         L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_12, 
         L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_11, 
         L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_10, 
         L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_9, 
         L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_8, 
         L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_7, 
         L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_6, 
         L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_5, 
         L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_4, 
         L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_3, 
         L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_2, 
         L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_1, 
         L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_0, 
         L1_0_L2_1_G1_MINI_ALU_OperationResult_15, 
         L1_0_L2_1_G1_MINI_ALU_OperationResult_14, 
         L1_0_L2_1_G1_MINI_ALU_OperationResult_13, 
         L1_0_L2_1_G1_MINI_ALU_OperationResult_12, 
         L1_0_L2_1_G1_MINI_ALU_OperationResult_11, 
         L1_0_L2_1_G1_MINI_ALU_OperationResult_10, 
         L1_0_L2_1_G1_MINI_ALU_OperationResult_9, 
         L1_0_L2_1_G1_MINI_ALU_OperationResult_8, 
         L1_0_L2_1_G1_MINI_ALU_OperationResult_7, 
         L1_0_L2_1_G1_MINI_ALU_OperationResult_6, 
         L1_0_L2_1_G1_MINI_ALU_OperationResult_5, 
         L1_0_L2_1_G1_MINI_ALU_OperationResult_4, 
         L1_0_L2_1_G1_MINI_ALU_OperationResult_3, 
         L1_0_L2_1_G1_MINI_ALU_OperationResult_2, 
         L1_0_L2_1_G1_MINI_ALU_OperationResult_1, 
         L1_0_L2_1_G1_MINI_ALU_OperationResult_0, 
         L1_0_L2_1_G1_MINI_ALU_BoothXORCheck, 
         L1_0_L2_1_G1_MINI_ALU_BoothOperand_16, 
         L1_0_L2_1_G1_MINI_ALU_BoothOperand_15, 
         L1_0_L2_1_G1_MINI_ALU_BoothOperand_14, 
         L1_0_L2_1_G1_MINI_ALU_BoothOperand_13, 
         L1_0_L2_1_G1_MINI_ALU_BoothOperand_12, 
         L1_0_L2_1_G1_MINI_ALU_BoothOperand_11, 
         L1_0_L2_1_G1_MINI_ALU_BoothOperand_10, 
         L1_0_L2_1_G1_MINI_ALU_BoothOperand_9, L1_0_L2_1_G1_MINI_ALU_BoothP_16, 
         L1_0_L2_1_G1_MINI_ALU_BoothP_15, L1_0_L2_1_G1_MINI_ALU_BoothP_14, 
         L1_0_L2_1_G1_MINI_ALU_BoothP_13, L1_0_L2_1_G1_MINI_ALU_BoothP_12, 
         L1_0_L2_1_G1_MINI_ALU_BoothP_11, L1_0_L2_1_G1_MINI_ALU_BoothP_10, 
         L1_0_L2_1_G1_MINI_ALU_BoothP_9, L1_0_L2_1_G1_MINI_ALU_BoothP_8, 
         L1_0_L2_1_G1_MINI_ALU_BoothP_7, L1_0_L2_1_G1_MINI_ALU_BoothP_6, 
         L1_0_L2_1_G1_MINI_ALU_BoothP_5, L1_0_L2_1_G1_MINI_ALU_BoothP_4, 
         L1_0_L2_1_G1_MINI_ALU_BoothP_3, L1_0_L2_1_G1_MINI_ALU_BoothP_2, 
         L1_0_L2_1_G1_MINI_ALU_BoothP_1, L1_0_L2_1_G1_MINI_ALU_BoothP_0, 
         L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_15, 
         L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_14, 
         L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_13, 
         L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_12, 
         L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_11, 
         L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_10, 
         L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_9, 
         L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_8, 
         L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_7, 
         L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_6, 
         L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_5, 
         L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_4, 
         L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_3, 
         L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_2, 
         L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_1, 
         L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_0, 
         L1_0_L2_2_G1_MINI_ALU_OperationResult_15, 
         L1_0_L2_2_G1_MINI_ALU_OperationResult_14, 
         L1_0_L2_2_G1_MINI_ALU_OperationResult_13, 
         L1_0_L2_2_G1_MINI_ALU_OperationResult_12, 
         L1_0_L2_2_G1_MINI_ALU_OperationResult_11, 
         L1_0_L2_2_G1_MINI_ALU_OperationResult_10, 
         L1_0_L2_2_G1_MINI_ALU_OperationResult_9, 
         L1_0_L2_2_G1_MINI_ALU_OperationResult_8, 
         L1_0_L2_2_G1_MINI_ALU_OperationResult_7, 
         L1_0_L2_2_G1_MINI_ALU_OperationResult_6, 
         L1_0_L2_2_G1_MINI_ALU_OperationResult_5, 
         L1_0_L2_2_G1_MINI_ALU_OperationResult_4, 
         L1_0_L2_2_G1_MINI_ALU_OperationResult_3, 
         L1_0_L2_2_G1_MINI_ALU_OperationResult_2, 
         L1_0_L2_2_G1_MINI_ALU_OperationResult_1, 
         L1_0_L2_2_G1_MINI_ALU_OperationResult_0, 
         L1_0_L2_2_G1_MINI_ALU_BoothXORCheck, 
         L1_0_L2_2_G1_MINI_ALU_BoothOperand_16, 
         L1_0_L2_2_G1_MINI_ALU_BoothOperand_15, 
         L1_0_L2_2_G1_MINI_ALU_BoothOperand_14, 
         L1_0_L2_2_G1_MINI_ALU_BoothOperand_13, 
         L1_0_L2_2_G1_MINI_ALU_BoothOperand_12, 
         L1_0_L2_2_G1_MINI_ALU_BoothOperand_11, 
         L1_0_L2_2_G1_MINI_ALU_BoothOperand_10, 
         L1_0_L2_2_G1_MINI_ALU_BoothOperand_9, L1_0_L2_2_G1_MINI_ALU_BoothP_16, 
         L1_0_L2_2_G1_MINI_ALU_BoothP_15, L1_0_L2_2_G1_MINI_ALU_BoothP_14, 
         L1_0_L2_2_G1_MINI_ALU_BoothP_13, L1_0_L2_2_G1_MINI_ALU_BoothP_12, 
         L1_0_L2_2_G1_MINI_ALU_BoothP_11, L1_0_L2_2_G1_MINI_ALU_BoothP_10, 
         L1_0_L2_2_G1_MINI_ALU_BoothP_9, L1_0_L2_2_G1_MINI_ALU_BoothP_8, 
         L1_0_L2_2_G1_MINI_ALU_BoothP_7, L1_0_L2_2_G1_MINI_ALU_BoothP_6, 
         L1_0_L2_2_G1_MINI_ALU_BoothP_5, L1_0_L2_2_G1_MINI_ALU_BoothP_4, 
         L1_0_L2_2_G1_MINI_ALU_BoothP_3, L1_0_L2_2_G1_MINI_ALU_BoothP_2, 
         L1_0_L2_2_G1_MINI_ALU_BoothP_1, L1_0_L2_2_G1_MINI_ALU_BoothP_0, 
         L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_15, 
         L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_14, 
         L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_13, 
         L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_12, 
         L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_11, 
         L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_10, 
         L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_9, 
         L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_8, 
         L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_7, 
         L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_6, 
         L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_5, 
         L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_4, 
         L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_3, 
         L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_2, 
         L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_1, 
         L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_0, 
         L1_0_L2_3_G1_MINI_ALU_OperationResult_15, 
         L1_0_L2_3_G1_MINI_ALU_OperationResult_14, 
         L1_0_L2_3_G1_MINI_ALU_OperationResult_13, 
         L1_0_L2_3_G1_MINI_ALU_OperationResult_12, 
         L1_0_L2_3_G1_MINI_ALU_OperationResult_11, 
         L1_0_L2_3_G1_MINI_ALU_OperationResult_10, 
         L1_0_L2_3_G1_MINI_ALU_OperationResult_9, 
         L1_0_L2_3_G1_MINI_ALU_OperationResult_8, 
         L1_0_L2_3_G1_MINI_ALU_OperationResult_7, 
         L1_0_L2_3_G1_MINI_ALU_OperationResult_6, 
         L1_0_L2_3_G1_MINI_ALU_OperationResult_5, 
         L1_0_L2_3_G1_MINI_ALU_OperationResult_4, 
         L1_0_L2_3_G1_MINI_ALU_OperationResult_3, 
         L1_0_L2_3_G1_MINI_ALU_OperationResult_2, 
         L1_0_L2_3_G1_MINI_ALU_OperationResult_1, 
         L1_0_L2_3_G1_MINI_ALU_OperationResult_0, 
         L1_0_L2_3_G1_MINI_ALU_BoothXORCheck, 
         L1_0_L2_3_G1_MINI_ALU_BoothOperand_16, 
         L1_0_L2_3_G1_MINI_ALU_BoothOperand_15, 
         L1_0_L2_3_G1_MINI_ALU_BoothOperand_14, 
         L1_0_L2_3_G1_MINI_ALU_BoothOperand_13, 
         L1_0_L2_3_G1_MINI_ALU_BoothOperand_12, 
         L1_0_L2_3_G1_MINI_ALU_BoothOperand_11, 
         L1_0_L2_3_G1_MINI_ALU_BoothOperand_10, 
         L1_0_L2_3_G1_MINI_ALU_BoothOperand_9, L1_0_L2_3_G1_MINI_ALU_BoothP_16, 
         L1_0_L2_3_G1_MINI_ALU_BoothP_15, L1_0_L2_3_G1_MINI_ALU_BoothP_14, 
         L1_0_L2_3_G1_MINI_ALU_BoothP_13, L1_0_L2_3_G1_MINI_ALU_BoothP_12, 
         L1_0_L2_3_G1_MINI_ALU_BoothP_11, L1_0_L2_3_G1_MINI_ALU_BoothP_10, 
         L1_0_L2_3_G1_MINI_ALU_BoothP_9, L1_0_L2_3_G1_MINI_ALU_BoothP_8, 
         L1_0_L2_3_G1_MINI_ALU_BoothP_7, L1_0_L2_3_G1_MINI_ALU_BoothP_6, 
         L1_0_L2_3_G1_MINI_ALU_BoothP_5, L1_0_L2_3_G1_MINI_ALU_BoothP_4, 
         L1_0_L2_3_G1_MINI_ALU_BoothP_3, L1_0_L2_3_G1_MINI_ALU_BoothP_2, 
         L1_0_L2_3_G1_MINI_ALU_BoothP_1, L1_0_L2_3_G1_MINI_ALU_BoothP_0, 
         L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_15, 
         L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_14, 
         L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_13, 
         L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_12, 
         L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_11, 
         L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_10, 
         L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_9, 
         L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_8, 
         L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_7, 
         L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_6, 
         L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_5, 
         L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_4, 
         L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_3, 
         L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_2, 
         L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_1, 
         L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_0, 
         L1_0_L2_4_G1_MINI_ALU_OperationResult_15, 
         L1_0_L2_4_G1_MINI_ALU_OperationResult_14, 
         L1_0_L2_4_G1_MINI_ALU_OperationResult_13, 
         L1_0_L2_4_G1_MINI_ALU_OperationResult_12, 
         L1_0_L2_4_G1_MINI_ALU_OperationResult_11, 
         L1_0_L2_4_G1_MINI_ALU_OperationResult_10, 
         L1_0_L2_4_G1_MINI_ALU_OperationResult_9, 
         L1_0_L2_4_G1_MINI_ALU_OperationResult_8, 
         L1_0_L2_4_G1_MINI_ALU_OperationResult_7, 
         L1_0_L2_4_G1_MINI_ALU_OperationResult_6, 
         L1_0_L2_4_G1_MINI_ALU_OperationResult_5, 
         L1_0_L2_4_G1_MINI_ALU_OperationResult_4, 
         L1_0_L2_4_G1_MINI_ALU_OperationResult_3, 
         L1_0_L2_4_G1_MINI_ALU_OperationResult_2, 
         L1_0_L2_4_G1_MINI_ALU_OperationResult_1, 
         L1_0_L2_4_G1_MINI_ALU_OperationResult_0, 
         L1_0_L2_4_G1_MINI_ALU_BoothXORCheck, 
         L1_0_L2_4_G1_MINI_ALU_BoothOperand_16, 
         L1_0_L2_4_G1_MINI_ALU_BoothOperand_15, 
         L1_0_L2_4_G1_MINI_ALU_BoothOperand_14, 
         L1_0_L2_4_G1_MINI_ALU_BoothOperand_13, 
         L1_0_L2_4_G1_MINI_ALU_BoothOperand_12, 
         L1_0_L2_4_G1_MINI_ALU_BoothOperand_11, 
         L1_0_L2_4_G1_MINI_ALU_BoothOperand_10, 
         L1_0_L2_4_G1_MINI_ALU_BoothOperand_9, L1_0_L2_4_G1_MINI_ALU_BoothP_16, 
         L1_0_L2_4_G1_MINI_ALU_BoothP_15, L1_0_L2_4_G1_MINI_ALU_BoothP_14, 
         L1_0_L2_4_G1_MINI_ALU_BoothP_13, L1_0_L2_4_G1_MINI_ALU_BoothP_12, 
         L1_0_L2_4_G1_MINI_ALU_BoothP_11, L1_0_L2_4_G1_MINI_ALU_BoothP_10, 
         L1_0_L2_4_G1_MINI_ALU_BoothP_9, L1_0_L2_4_G1_MINI_ALU_BoothP_8, 
         L1_0_L2_4_G1_MINI_ALU_BoothP_7, L1_0_L2_4_G1_MINI_ALU_BoothP_6, 
         L1_0_L2_4_G1_MINI_ALU_BoothP_5, L1_0_L2_4_G1_MINI_ALU_BoothP_4, 
         L1_0_L2_4_G1_MINI_ALU_BoothP_3, L1_0_L2_4_G1_MINI_ALU_BoothP_2, 
         L1_0_L2_4_G1_MINI_ALU_BoothP_1, L1_0_L2_4_G1_MINI_ALU_BoothP_0, 
         L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_15, 
         L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_14, 
         L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_13, 
         L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_12, 
         L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_11, 
         L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_10, 
         L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_9, 
         L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_8, 
         L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_7, 
         L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_6, 
         L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_5, 
         L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_4, 
         L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_3, 
         L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_2, 
         L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_1, 
         L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_0, 
         L1_1_L2_0_G1_MINI_ALU_OperationResult_15, 
         L1_1_L2_0_G1_MINI_ALU_OperationResult_14, 
         L1_1_L2_0_G1_MINI_ALU_OperationResult_13, 
         L1_1_L2_0_G1_MINI_ALU_OperationResult_12, 
         L1_1_L2_0_G1_MINI_ALU_OperationResult_11, 
         L1_1_L2_0_G1_MINI_ALU_OperationResult_10, 
         L1_1_L2_0_G1_MINI_ALU_OperationResult_9, 
         L1_1_L2_0_G1_MINI_ALU_OperationResult_8, 
         L1_1_L2_0_G1_MINI_ALU_OperationResult_7, 
         L1_1_L2_0_G1_MINI_ALU_OperationResult_6, 
         L1_1_L2_0_G1_MINI_ALU_OperationResult_5, 
         L1_1_L2_0_G1_MINI_ALU_OperationResult_4, 
         L1_1_L2_0_G1_MINI_ALU_OperationResult_3, 
         L1_1_L2_0_G1_MINI_ALU_OperationResult_2, 
         L1_1_L2_0_G1_MINI_ALU_OperationResult_1, 
         L1_1_L2_0_G1_MINI_ALU_OperationResult_0, 
         L1_1_L2_0_G1_MINI_ALU_BoothXORCheck, 
         L1_1_L2_0_G1_MINI_ALU_BoothOperand_16, 
         L1_1_L2_0_G1_MINI_ALU_BoothOperand_15, 
         L1_1_L2_0_G1_MINI_ALU_BoothOperand_14, 
         L1_1_L2_0_G1_MINI_ALU_BoothOperand_13, 
         L1_1_L2_0_G1_MINI_ALU_BoothOperand_12, 
         L1_1_L2_0_G1_MINI_ALU_BoothOperand_11, 
         L1_1_L2_0_G1_MINI_ALU_BoothOperand_10, 
         L1_1_L2_0_G1_MINI_ALU_BoothOperand_9, L1_1_L2_0_G1_MINI_ALU_BoothP_16, 
         L1_1_L2_0_G1_MINI_ALU_BoothP_15, L1_1_L2_0_G1_MINI_ALU_BoothP_14, 
         L1_1_L2_0_G1_MINI_ALU_BoothP_13, L1_1_L2_0_G1_MINI_ALU_BoothP_12, 
         L1_1_L2_0_G1_MINI_ALU_BoothP_11, L1_1_L2_0_G1_MINI_ALU_BoothP_10, 
         L1_1_L2_0_G1_MINI_ALU_BoothP_9, L1_1_L2_0_G1_MINI_ALU_BoothP_8, 
         L1_1_L2_0_G1_MINI_ALU_BoothP_7, L1_1_L2_0_G1_MINI_ALU_BoothP_6, 
         L1_1_L2_0_G1_MINI_ALU_BoothP_5, L1_1_L2_0_G1_MINI_ALU_BoothP_4, 
         L1_1_L2_0_G1_MINI_ALU_BoothP_3, L1_1_L2_0_G1_MINI_ALU_BoothP_2, 
         L1_1_L2_0_G1_MINI_ALU_BoothP_1, L1_1_L2_0_G1_MINI_ALU_BoothP_0, 
         L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_15, 
         L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_14, 
         L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_13, 
         L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_12, 
         L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_11, 
         L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_10, 
         L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_9, 
         L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_8, 
         L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_7, 
         L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_6, 
         L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_5, 
         L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_4, 
         L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_3, 
         L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_2, 
         L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_1, 
         L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_0, 
         L1_1_L2_1_G1_MINI_ALU_OperationResult_15, 
         L1_1_L2_1_G1_MINI_ALU_OperationResult_14, 
         L1_1_L2_1_G1_MINI_ALU_OperationResult_13, 
         L1_1_L2_1_G1_MINI_ALU_OperationResult_12, 
         L1_1_L2_1_G1_MINI_ALU_OperationResult_11, 
         L1_1_L2_1_G1_MINI_ALU_OperationResult_10, 
         L1_1_L2_1_G1_MINI_ALU_OperationResult_9, 
         L1_1_L2_1_G1_MINI_ALU_OperationResult_8, 
         L1_1_L2_1_G1_MINI_ALU_OperationResult_7, 
         L1_1_L2_1_G1_MINI_ALU_OperationResult_6, 
         L1_1_L2_1_G1_MINI_ALU_OperationResult_5, 
         L1_1_L2_1_G1_MINI_ALU_OperationResult_4, 
         L1_1_L2_1_G1_MINI_ALU_OperationResult_3, 
         L1_1_L2_1_G1_MINI_ALU_OperationResult_2, 
         L1_1_L2_1_G1_MINI_ALU_OperationResult_1, 
         L1_1_L2_1_G1_MINI_ALU_OperationResult_0, 
         L1_1_L2_1_G1_MINI_ALU_BoothXORCheck, 
         L1_1_L2_1_G1_MINI_ALU_BoothOperand_16, 
         L1_1_L2_1_G1_MINI_ALU_BoothOperand_15, 
         L1_1_L2_1_G1_MINI_ALU_BoothOperand_14, 
         L1_1_L2_1_G1_MINI_ALU_BoothOperand_13, 
         L1_1_L2_1_G1_MINI_ALU_BoothOperand_12, 
         L1_1_L2_1_G1_MINI_ALU_BoothOperand_11, 
         L1_1_L2_1_G1_MINI_ALU_BoothOperand_10, 
         L1_1_L2_1_G1_MINI_ALU_BoothOperand_9, L1_1_L2_1_G1_MINI_ALU_BoothP_16, 
         L1_1_L2_1_G1_MINI_ALU_BoothP_15, L1_1_L2_1_G1_MINI_ALU_BoothP_14, 
         L1_1_L2_1_G1_MINI_ALU_BoothP_13, L1_1_L2_1_G1_MINI_ALU_BoothP_12, 
         L1_1_L2_1_G1_MINI_ALU_BoothP_11, L1_1_L2_1_G1_MINI_ALU_BoothP_10, 
         L1_1_L2_1_G1_MINI_ALU_BoothP_9, L1_1_L2_1_G1_MINI_ALU_BoothP_8, 
         L1_1_L2_1_G1_MINI_ALU_BoothP_7, L1_1_L2_1_G1_MINI_ALU_BoothP_6, 
         L1_1_L2_1_G1_MINI_ALU_BoothP_5, L1_1_L2_1_G1_MINI_ALU_BoothP_4, 
         L1_1_L2_1_G1_MINI_ALU_BoothP_3, L1_1_L2_1_G1_MINI_ALU_BoothP_2, 
         L1_1_L2_1_G1_MINI_ALU_BoothP_1, L1_1_L2_1_G1_MINI_ALU_BoothP_0, 
         L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_15, 
         L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_14, 
         L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_13, 
         L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_12, 
         L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_11, 
         L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_10, 
         L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_9, 
         L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_8, 
         L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_7, 
         L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_6, 
         L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_5, 
         L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_4, 
         L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_3, 
         L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_2, 
         L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_1, 
         L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_0, 
         L1_1_L2_2_G1_MINI_ALU_OperationResult_15, 
         L1_1_L2_2_G1_MINI_ALU_OperationResult_14, 
         L1_1_L2_2_G1_MINI_ALU_OperationResult_13, 
         L1_1_L2_2_G1_MINI_ALU_OperationResult_12, 
         L1_1_L2_2_G1_MINI_ALU_OperationResult_11, 
         L1_1_L2_2_G1_MINI_ALU_OperationResult_10, 
         L1_1_L2_2_G1_MINI_ALU_OperationResult_9, 
         L1_1_L2_2_G1_MINI_ALU_OperationResult_8, 
         L1_1_L2_2_G1_MINI_ALU_OperationResult_7, 
         L1_1_L2_2_G1_MINI_ALU_OperationResult_6, 
         L1_1_L2_2_G1_MINI_ALU_OperationResult_5, 
         L1_1_L2_2_G1_MINI_ALU_OperationResult_4, 
         L1_1_L2_2_G1_MINI_ALU_OperationResult_3, 
         L1_1_L2_2_G1_MINI_ALU_OperationResult_2, 
         L1_1_L2_2_G1_MINI_ALU_OperationResult_1, 
         L1_1_L2_2_G1_MINI_ALU_OperationResult_0, 
         L1_1_L2_2_G1_MINI_ALU_BoothXORCheck, 
         L1_1_L2_2_G1_MINI_ALU_BoothOperand_16, 
         L1_1_L2_2_G1_MINI_ALU_BoothOperand_15, 
         L1_1_L2_2_G1_MINI_ALU_BoothOperand_14, 
         L1_1_L2_2_G1_MINI_ALU_BoothOperand_13, 
         L1_1_L2_2_G1_MINI_ALU_BoothOperand_12, 
         L1_1_L2_2_G1_MINI_ALU_BoothOperand_11, 
         L1_1_L2_2_G1_MINI_ALU_BoothOperand_10, 
         L1_1_L2_2_G1_MINI_ALU_BoothOperand_9, L1_1_L2_2_G1_MINI_ALU_BoothP_16, 
         L1_1_L2_2_G1_MINI_ALU_BoothP_15, L1_1_L2_2_G1_MINI_ALU_BoothP_14, 
         L1_1_L2_2_G1_MINI_ALU_BoothP_13, L1_1_L2_2_G1_MINI_ALU_BoothP_12, 
         L1_1_L2_2_G1_MINI_ALU_BoothP_11, L1_1_L2_2_G1_MINI_ALU_BoothP_10, 
         L1_1_L2_2_G1_MINI_ALU_BoothP_9, L1_1_L2_2_G1_MINI_ALU_BoothP_8, 
         L1_1_L2_2_G1_MINI_ALU_BoothP_7, L1_1_L2_2_G1_MINI_ALU_BoothP_6, 
         L1_1_L2_2_G1_MINI_ALU_BoothP_5, L1_1_L2_2_G1_MINI_ALU_BoothP_4, 
         L1_1_L2_2_G1_MINI_ALU_BoothP_3, L1_1_L2_2_G1_MINI_ALU_BoothP_2, 
         L1_1_L2_2_G1_MINI_ALU_BoothP_1, L1_1_L2_2_G1_MINI_ALU_BoothP_0, 
         L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_15, 
         L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_14, 
         L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_13, 
         L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_12, 
         L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_11, 
         L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_10, 
         L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_9, 
         L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_8, 
         L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_7, 
         L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_6, 
         L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_5, 
         L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_4, 
         L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_3, 
         L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_2, 
         L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_1, 
         L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_0, 
         L1_1_L2_3_G1_MINI_ALU_OperationResult_15, 
         L1_1_L2_3_G1_MINI_ALU_OperationResult_14, 
         L1_1_L2_3_G1_MINI_ALU_OperationResult_13, 
         L1_1_L2_3_G1_MINI_ALU_OperationResult_12, 
         L1_1_L2_3_G1_MINI_ALU_OperationResult_11, 
         L1_1_L2_3_G1_MINI_ALU_OperationResult_10, 
         L1_1_L2_3_G1_MINI_ALU_OperationResult_9, 
         L1_1_L2_3_G1_MINI_ALU_OperationResult_8, 
         L1_1_L2_3_G1_MINI_ALU_OperationResult_7, 
         L1_1_L2_3_G1_MINI_ALU_OperationResult_6, 
         L1_1_L2_3_G1_MINI_ALU_OperationResult_5, 
         L1_1_L2_3_G1_MINI_ALU_OperationResult_4, 
         L1_1_L2_3_G1_MINI_ALU_OperationResult_3, 
         L1_1_L2_3_G1_MINI_ALU_OperationResult_2, 
         L1_1_L2_3_G1_MINI_ALU_OperationResult_1, 
         L1_1_L2_3_G1_MINI_ALU_OperationResult_0, 
         L1_1_L2_3_G1_MINI_ALU_BoothXORCheck, 
         L1_1_L2_3_G1_MINI_ALU_BoothOperand_16, 
         L1_1_L2_3_G1_MINI_ALU_BoothOperand_15, 
         L1_1_L2_3_G1_MINI_ALU_BoothOperand_14, 
         L1_1_L2_3_G1_MINI_ALU_BoothOperand_13, 
         L1_1_L2_3_G1_MINI_ALU_BoothOperand_12, 
         L1_1_L2_3_G1_MINI_ALU_BoothOperand_11, 
         L1_1_L2_3_G1_MINI_ALU_BoothOperand_10, 
         L1_1_L2_3_G1_MINI_ALU_BoothOperand_9, L1_1_L2_3_G1_MINI_ALU_BoothP_16, 
         L1_1_L2_3_G1_MINI_ALU_BoothP_15, L1_1_L2_3_G1_MINI_ALU_BoothP_14, 
         L1_1_L2_3_G1_MINI_ALU_BoothP_13, L1_1_L2_3_G1_MINI_ALU_BoothP_12, 
         L1_1_L2_3_G1_MINI_ALU_BoothP_11, L1_1_L2_3_G1_MINI_ALU_BoothP_10, 
         L1_1_L2_3_G1_MINI_ALU_BoothP_9, L1_1_L2_3_G1_MINI_ALU_BoothP_8, 
         L1_1_L2_3_G1_MINI_ALU_BoothP_7, L1_1_L2_3_G1_MINI_ALU_BoothP_6, 
         L1_1_L2_3_G1_MINI_ALU_BoothP_5, L1_1_L2_3_G1_MINI_ALU_BoothP_4, 
         L1_1_L2_3_G1_MINI_ALU_BoothP_3, L1_1_L2_3_G1_MINI_ALU_BoothP_2, 
         L1_1_L2_3_G1_MINI_ALU_BoothP_1, L1_1_L2_3_G1_MINI_ALU_BoothP_0, 
         L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_15, 
         L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_14, 
         L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_13, 
         L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_12, 
         L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_11, 
         L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_10, 
         L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_9, 
         L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_8, 
         L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_7, 
         L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_6, 
         L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_5, 
         L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_4, 
         L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_3, 
         L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_2, 
         L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_1, 
         L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_0, 
         L1_1_L2_4_G1_MINI_ALU_OperationResult_15, 
         L1_1_L2_4_G1_MINI_ALU_OperationResult_14, 
         L1_1_L2_4_G1_MINI_ALU_OperationResult_13, 
         L1_1_L2_4_G1_MINI_ALU_OperationResult_12, 
         L1_1_L2_4_G1_MINI_ALU_OperationResult_11, 
         L1_1_L2_4_G1_MINI_ALU_OperationResult_10, 
         L1_1_L2_4_G1_MINI_ALU_OperationResult_9, 
         L1_1_L2_4_G1_MINI_ALU_OperationResult_8, 
         L1_1_L2_4_G1_MINI_ALU_OperationResult_7, 
         L1_1_L2_4_G1_MINI_ALU_OperationResult_6, 
         L1_1_L2_4_G1_MINI_ALU_OperationResult_5, 
         L1_1_L2_4_G1_MINI_ALU_OperationResult_4, 
         L1_1_L2_4_G1_MINI_ALU_OperationResult_3, 
         L1_1_L2_4_G1_MINI_ALU_OperationResult_2, 
         L1_1_L2_4_G1_MINI_ALU_OperationResult_1, 
         L1_1_L2_4_G1_MINI_ALU_OperationResult_0, 
         L1_1_L2_4_G1_MINI_ALU_BoothXORCheck, 
         L1_1_L2_4_G1_MINI_ALU_BoothOperand_16, 
         L1_1_L2_4_G1_MINI_ALU_BoothOperand_15, 
         L1_1_L2_4_G1_MINI_ALU_BoothOperand_14, 
         L1_1_L2_4_G1_MINI_ALU_BoothOperand_13, 
         L1_1_L2_4_G1_MINI_ALU_BoothOperand_12, 
         L1_1_L2_4_G1_MINI_ALU_BoothOperand_11, 
         L1_1_L2_4_G1_MINI_ALU_BoothOperand_10, 
         L1_1_L2_4_G1_MINI_ALU_BoothOperand_9, L1_1_L2_4_G1_MINI_ALU_BoothP_16, 
         L1_1_L2_4_G1_MINI_ALU_BoothP_15, L1_1_L2_4_G1_MINI_ALU_BoothP_14, 
         L1_1_L2_4_G1_MINI_ALU_BoothP_13, L1_1_L2_4_G1_MINI_ALU_BoothP_12, 
         L1_1_L2_4_G1_MINI_ALU_BoothP_11, L1_1_L2_4_G1_MINI_ALU_BoothP_10, 
         L1_1_L2_4_G1_MINI_ALU_BoothP_9, L1_1_L2_4_G1_MINI_ALU_BoothP_8, 
         L1_1_L2_4_G1_MINI_ALU_BoothP_7, L1_1_L2_4_G1_MINI_ALU_BoothP_6, 
         L1_1_L2_4_G1_MINI_ALU_BoothP_5, L1_1_L2_4_G1_MINI_ALU_BoothP_4, 
         L1_1_L2_4_G1_MINI_ALU_BoothP_3, L1_1_L2_4_G1_MINI_ALU_BoothP_2, 
         L1_1_L2_4_G1_MINI_ALU_BoothP_1, L1_1_L2_4_G1_MINI_ALU_BoothP_0, 
         L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_15, 
         L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_14, 
         L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_13, 
         L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_12, 
         L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_11, 
         L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_10, 
         L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_9, 
         L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_8, 
         L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_7, 
         L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_6, 
         L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_5, 
         L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_4, 
         L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_3, 
         L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_2, 
         L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_1, 
         L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_0, 
         L1_2_L2_0_G1_MINI_ALU_OperationResult_15, 
         L1_2_L2_0_G1_MINI_ALU_OperationResult_14, 
         L1_2_L2_0_G1_MINI_ALU_OperationResult_13, 
         L1_2_L2_0_G1_MINI_ALU_OperationResult_12, 
         L1_2_L2_0_G1_MINI_ALU_OperationResult_11, 
         L1_2_L2_0_G1_MINI_ALU_OperationResult_10, 
         L1_2_L2_0_G1_MINI_ALU_OperationResult_9, 
         L1_2_L2_0_G1_MINI_ALU_OperationResult_8, 
         L1_2_L2_0_G1_MINI_ALU_OperationResult_7, 
         L1_2_L2_0_G1_MINI_ALU_OperationResult_6, 
         L1_2_L2_0_G1_MINI_ALU_OperationResult_5, 
         L1_2_L2_0_G1_MINI_ALU_OperationResult_4, 
         L1_2_L2_0_G1_MINI_ALU_OperationResult_3, 
         L1_2_L2_0_G1_MINI_ALU_OperationResult_2, 
         L1_2_L2_0_G1_MINI_ALU_OperationResult_1, 
         L1_2_L2_0_G1_MINI_ALU_OperationResult_0, 
         L1_2_L2_0_G1_MINI_ALU_BoothXORCheck, 
         L1_2_L2_0_G1_MINI_ALU_BoothOperand_16, 
         L1_2_L2_0_G1_MINI_ALU_BoothOperand_15, 
         L1_2_L2_0_G1_MINI_ALU_BoothOperand_14, 
         L1_2_L2_0_G1_MINI_ALU_BoothOperand_13, 
         L1_2_L2_0_G1_MINI_ALU_BoothOperand_12, 
         L1_2_L2_0_G1_MINI_ALU_BoothOperand_11, 
         L1_2_L2_0_G1_MINI_ALU_BoothOperand_10, 
         L1_2_L2_0_G1_MINI_ALU_BoothOperand_9, L1_2_L2_0_G1_MINI_ALU_BoothP_16, 
         L1_2_L2_0_G1_MINI_ALU_BoothP_15, L1_2_L2_0_G1_MINI_ALU_BoothP_14, 
         L1_2_L2_0_G1_MINI_ALU_BoothP_13, L1_2_L2_0_G1_MINI_ALU_BoothP_12, 
         L1_2_L2_0_G1_MINI_ALU_BoothP_11, L1_2_L2_0_G1_MINI_ALU_BoothP_10, 
         L1_2_L2_0_G1_MINI_ALU_BoothP_9, L1_2_L2_0_G1_MINI_ALU_BoothP_8, 
         L1_2_L2_0_G1_MINI_ALU_BoothP_7, L1_2_L2_0_G1_MINI_ALU_BoothP_6, 
         L1_2_L2_0_G1_MINI_ALU_BoothP_5, L1_2_L2_0_G1_MINI_ALU_BoothP_4, 
         L1_2_L2_0_G1_MINI_ALU_BoothP_3, L1_2_L2_0_G1_MINI_ALU_BoothP_2, 
         L1_2_L2_0_G1_MINI_ALU_BoothP_1, L1_2_L2_0_G1_MINI_ALU_BoothP_0, 
         L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_15, 
         L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_14, 
         L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_13, 
         L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_12, 
         L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_11, 
         L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_10, 
         L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_9, 
         L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_8, 
         L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_7, 
         L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_6, 
         L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_5, 
         L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_4, 
         L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_3, 
         L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_2, 
         L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_1, 
         L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_0, 
         L1_2_L2_1_G1_MINI_ALU_OperationResult_15, 
         L1_2_L2_1_G1_MINI_ALU_OperationResult_14, 
         L1_2_L2_1_G1_MINI_ALU_OperationResult_13, 
         L1_2_L2_1_G1_MINI_ALU_OperationResult_12, 
         L1_2_L2_1_G1_MINI_ALU_OperationResult_11, 
         L1_2_L2_1_G1_MINI_ALU_OperationResult_10, 
         L1_2_L2_1_G1_MINI_ALU_OperationResult_9, 
         L1_2_L2_1_G1_MINI_ALU_OperationResult_8, 
         L1_2_L2_1_G1_MINI_ALU_OperationResult_7, 
         L1_2_L2_1_G1_MINI_ALU_OperationResult_6, 
         L1_2_L2_1_G1_MINI_ALU_OperationResult_5, 
         L1_2_L2_1_G1_MINI_ALU_OperationResult_4, 
         L1_2_L2_1_G1_MINI_ALU_OperationResult_3, 
         L1_2_L2_1_G1_MINI_ALU_OperationResult_2, 
         L1_2_L2_1_G1_MINI_ALU_OperationResult_1, 
         L1_2_L2_1_G1_MINI_ALU_OperationResult_0, 
         L1_2_L2_1_G1_MINI_ALU_BoothXORCheck, 
         L1_2_L2_1_G1_MINI_ALU_BoothOperand_16, 
         L1_2_L2_1_G1_MINI_ALU_BoothOperand_15, 
         L1_2_L2_1_G1_MINI_ALU_BoothOperand_14, 
         L1_2_L2_1_G1_MINI_ALU_BoothOperand_13, 
         L1_2_L2_1_G1_MINI_ALU_BoothOperand_12, 
         L1_2_L2_1_G1_MINI_ALU_BoothOperand_11, 
         L1_2_L2_1_G1_MINI_ALU_BoothOperand_10, 
         L1_2_L2_1_G1_MINI_ALU_BoothOperand_9, L1_2_L2_1_G1_MINI_ALU_BoothP_16, 
         L1_2_L2_1_G1_MINI_ALU_BoothP_15, L1_2_L2_1_G1_MINI_ALU_BoothP_14, 
         L1_2_L2_1_G1_MINI_ALU_BoothP_13, L1_2_L2_1_G1_MINI_ALU_BoothP_12, 
         L1_2_L2_1_G1_MINI_ALU_BoothP_11, L1_2_L2_1_G1_MINI_ALU_BoothP_10, 
         L1_2_L2_1_G1_MINI_ALU_BoothP_9, L1_2_L2_1_G1_MINI_ALU_BoothP_8, 
         L1_2_L2_1_G1_MINI_ALU_BoothP_7, L1_2_L2_1_G1_MINI_ALU_BoothP_6, 
         L1_2_L2_1_G1_MINI_ALU_BoothP_5, L1_2_L2_1_G1_MINI_ALU_BoothP_4, 
         L1_2_L2_1_G1_MINI_ALU_BoothP_3, L1_2_L2_1_G1_MINI_ALU_BoothP_2, 
         L1_2_L2_1_G1_MINI_ALU_BoothP_1, L1_2_L2_1_G1_MINI_ALU_BoothP_0, 
         L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_15, 
         L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_14, 
         L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_13, 
         L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_12, 
         L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_11, 
         L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_10, 
         L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_9, 
         L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_8, 
         L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_7, 
         L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_6, 
         L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_5, 
         L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_4, 
         L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_3, 
         L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_2, 
         L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_1, 
         L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_0, 
         L1_2_L2_2_G1_MINI_ALU_BoothXORCheck, 
         L1_2_L2_2_G1_MINI_ALU_BoothOperand_16, 
         L1_2_L2_2_G1_MINI_ALU_BoothOperand_15, 
         L1_2_L2_2_G1_MINI_ALU_BoothOperand_14, 
         L1_2_L2_2_G1_MINI_ALU_BoothOperand_13, 
         L1_2_L2_2_G1_MINI_ALU_BoothOperand_12, 
         L1_2_L2_2_G1_MINI_ALU_BoothOperand_11, 
         L1_2_L2_2_G1_MINI_ALU_BoothOperand_10, 
         L1_2_L2_2_G1_MINI_ALU_BoothOperand_9, L1_2_L2_2_G1_MINI_ALU_BoothP_16, 
         L1_2_L2_2_G1_MINI_ALU_BoothP_15, L1_2_L2_2_G1_MINI_ALU_BoothP_14, 
         L1_2_L2_2_G1_MINI_ALU_BoothP_13, L1_2_L2_2_G1_MINI_ALU_BoothP_12, 
         L1_2_L2_2_G1_MINI_ALU_BoothP_11, L1_2_L2_2_G1_MINI_ALU_BoothP_10, 
         L1_2_L2_2_G1_MINI_ALU_BoothP_9, L1_2_L2_2_G1_MINI_ALU_BoothP_8, 
         L1_2_L2_2_G1_MINI_ALU_BoothP_7, L1_2_L2_2_G1_MINI_ALU_BoothP_6, 
         L1_2_L2_2_G1_MINI_ALU_BoothP_5, L1_2_L2_2_G1_MINI_ALU_BoothP_4, 
         L1_2_L2_2_G1_MINI_ALU_BoothP_3, L1_2_L2_2_G1_MINI_ALU_BoothP_2, 
         L1_2_L2_2_G1_MINI_ALU_BoothP_1, 
         L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_15, 
         L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_14, 
         L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_13, 
         L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_12, 
         L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_11, 
         L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_10, 
         L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_9, 
         L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_8, 
         L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_7, 
         L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_6, 
         L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_5, 
         L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_4, 
         L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_3, 
         L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_2, 
         L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_1, 
         L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_0, 
         L1_2_L2_3_G2_MINI_ALU_BoothXORCheck, 
         L1_2_L2_3_G2_MINI_ALU_BoothOperand_16, 
         L1_2_L2_3_G2_MINI_ALU_BoothOperand_15, 
         L1_2_L2_3_G2_MINI_ALU_BoothOperand_14, 
         L1_2_L2_3_G2_MINI_ALU_BoothOperand_13, 
         L1_2_L2_3_G2_MINI_ALU_BoothOperand_12, 
         L1_2_L2_3_G2_MINI_ALU_BoothOperand_11, 
         L1_2_L2_3_G2_MINI_ALU_BoothOperand_10, 
         L1_2_L2_3_G2_MINI_ALU_BoothOperand_9, L1_2_L2_3_G2_MINI_ALU_BoothP_16, 
         L1_2_L2_3_G2_MINI_ALU_BoothP_15, L1_2_L2_3_G2_MINI_ALU_BoothP_14, 
         L1_2_L2_3_G2_MINI_ALU_BoothP_13, L1_2_L2_3_G2_MINI_ALU_BoothP_12, 
         L1_2_L2_3_G2_MINI_ALU_BoothP_11, L1_2_L2_3_G2_MINI_ALU_BoothP_10, 
         L1_2_L2_3_G2_MINI_ALU_BoothP_9, L1_2_L2_3_G2_MINI_ALU_BoothP_8, 
         L1_2_L2_3_G2_MINI_ALU_BoothP_7, L1_2_L2_3_G2_MINI_ALU_BoothP_6, 
         L1_2_L2_3_G2_MINI_ALU_BoothP_5, L1_2_L2_3_G2_MINI_ALU_BoothP_4, 
         L1_2_L2_3_G2_MINI_ALU_BoothP_3, L1_2_L2_3_G2_MINI_ALU_BoothP_2, 
         L1_2_L2_3_G2_MINI_ALU_BoothP_1, L1_2_L2_3_G2_MINI_ALU_BoothP_0, 
         L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_15, 
         L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_14, 
         L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_13, 
         L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_12, 
         L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_11, 
         L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_10, 
         L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_9, 
         L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_8, 
         L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_7, 
         L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_6, 
         L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_5, 
         L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_4, 
         L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_3, 
         L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_2, 
         L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_1, 
         L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_0, 
         L1_2_L2_4_G2_MINI_ALU_BoothXORCheck, 
         L1_2_L2_4_G2_MINI_ALU_BoothOperand_16, 
         L1_2_L2_4_G2_MINI_ALU_BoothOperand_15, 
         L1_2_L2_4_G2_MINI_ALU_BoothOperand_14, 
         L1_2_L2_4_G2_MINI_ALU_BoothOperand_13, 
         L1_2_L2_4_G2_MINI_ALU_BoothOperand_12, 
         L1_2_L2_4_G2_MINI_ALU_BoothOperand_11, 
         L1_2_L2_4_G2_MINI_ALU_BoothOperand_10, 
         L1_2_L2_4_G2_MINI_ALU_BoothOperand_9, L1_2_L2_4_G2_MINI_ALU_BoothP_16, 
         L1_2_L2_4_G2_MINI_ALU_BoothP_15, L1_2_L2_4_G2_MINI_ALU_BoothP_14, 
         L1_2_L2_4_G2_MINI_ALU_BoothP_13, L1_2_L2_4_G2_MINI_ALU_BoothP_12, 
         L1_2_L2_4_G2_MINI_ALU_BoothP_11, L1_2_L2_4_G2_MINI_ALU_BoothP_10, 
         L1_2_L2_4_G2_MINI_ALU_BoothP_9, L1_2_L2_4_G2_MINI_ALU_BoothP_8, 
         L1_2_L2_4_G2_MINI_ALU_BoothP_7, L1_2_L2_4_G2_MINI_ALU_BoothP_6, 
         L1_2_L2_4_G2_MINI_ALU_BoothP_5, L1_2_L2_4_G2_MINI_ALU_BoothP_4, 
         L1_2_L2_4_G2_MINI_ALU_BoothP_3, L1_2_L2_4_G2_MINI_ALU_BoothP_2, 
         L1_2_L2_4_G2_MINI_ALU_BoothP_1, L1_2_L2_4_G2_MINI_ALU_BoothP_0, 
         L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_15, 
         L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_14, 
         L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_13, 
         L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_12, 
         L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_11, 
         L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_10, 
         L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_9, 
         L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_8, 
         L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_7, 
         L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_6, 
         L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_5, 
         L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_4, 
         L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_3, 
         L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_2, 
         L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_1, 
         L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_0, 
         L1_3_L2_0_G2_MINI_ALU_BoothXORCheck, 
         L1_3_L2_0_G2_MINI_ALU_BoothOperand_16, 
         L1_3_L2_0_G2_MINI_ALU_BoothOperand_15, 
         L1_3_L2_0_G2_MINI_ALU_BoothOperand_14, 
         L1_3_L2_0_G2_MINI_ALU_BoothOperand_13, 
         L1_3_L2_0_G2_MINI_ALU_BoothOperand_12, 
         L1_3_L2_0_G2_MINI_ALU_BoothOperand_11, 
         L1_3_L2_0_G2_MINI_ALU_BoothOperand_10, 
         L1_3_L2_0_G2_MINI_ALU_BoothOperand_9, L1_3_L2_0_G2_MINI_ALU_BoothP_16, 
         L1_3_L2_0_G2_MINI_ALU_BoothP_15, L1_3_L2_0_G2_MINI_ALU_BoothP_14, 
         L1_3_L2_0_G2_MINI_ALU_BoothP_13, L1_3_L2_0_G2_MINI_ALU_BoothP_12, 
         L1_3_L2_0_G2_MINI_ALU_BoothP_11, L1_3_L2_0_G2_MINI_ALU_BoothP_10, 
         L1_3_L2_0_G2_MINI_ALU_BoothP_9, L1_3_L2_0_G2_MINI_ALU_BoothP_8, 
         L1_3_L2_0_G2_MINI_ALU_BoothP_7, L1_3_L2_0_G2_MINI_ALU_BoothP_6, 
         L1_3_L2_0_G2_MINI_ALU_BoothP_5, L1_3_L2_0_G2_MINI_ALU_BoothP_4, 
         L1_3_L2_0_G2_MINI_ALU_BoothP_3, L1_3_L2_0_G2_MINI_ALU_BoothP_2, 
         L1_3_L2_0_G2_MINI_ALU_BoothP_1, L1_3_L2_0_G2_MINI_ALU_BoothP_0, 
         L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_15, 
         L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_14, 
         L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_13, 
         L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_12, 
         L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_11, 
         L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_10, 
         L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_9, 
         L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_8, 
         L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_7, 
         L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_6, 
         L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_5, 
         L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_4, 
         L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_3, 
         L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_2, 
         L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_1, 
         L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_0, 
         L1_3_L2_1_G2_MINI_ALU_BoothXORCheck, 
         L1_3_L2_1_G2_MINI_ALU_BoothOperand_16, 
         L1_3_L2_1_G2_MINI_ALU_BoothOperand_15, 
         L1_3_L2_1_G2_MINI_ALU_BoothOperand_14, 
         L1_3_L2_1_G2_MINI_ALU_BoothOperand_13, 
         L1_3_L2_1_G2_MINI_ALU_BoothOperand_12, 
         L1_3_L2_1_G2_MINI_ALU_BoothOperand_11, 
         L1_3_L2_1_G2_MINI_ALU_BoothOperand_10, 
         L1_3_L2_1_G2_MINI_ALU_BoothOperand_9, L1_3_L2_1_G2_MINI_ALU_BoothP_16, 
         L1_3_L2_1_G2_MINI_ALU_BoothP_15, L1_3_L2_1_G2_MINI_ALU_BoothP_14, 
         L1_3_L2_1_G2_MINI_ALU_BoothP_13, L1_3_L2_1_G2_MINI_ALU_BoothP_12, 
         L1_3_L2_1_G2_MINI_ALU_BoothP_11, L1_3_L2_1_G2_MINI_ALU_BoothP_10, 
         L1_3_L2_1_G2_MINI_ALU_BoothP_9, L1_3_L2_1_G2_MINI_ALU_BoothP_8, 
         L1_3_L2_1_G2_MINI_ALU_BoothP_7, L1_3_L2_1_G2_MINI_ALU_BoothP_6, 
         L1_3_L2_1_G2_MINI_ALU_BoothP_5, L1_3_L2_1_G2_MINI_ALU_BoothP_4, 
         L1_3_L2_1_G2_MINI_ALU_BoothP_3, L1_3_L2_1_G2_MINI_ALU_BoothP_2, 
         L1_3_L2_1_G2_MINI_ALU_BoothP_1, L1_3_L2_1_G2_MINI_ALU_BoothP_0, 
         L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_15, 
         L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_14, 
         L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_13, 
         L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_12, 
         L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_11, 
         L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_10, 
         L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_9, 
         L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_8, 
         L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_7, 
         L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_6, 
         L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_5, 
         L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_4, 
         L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_3, 
         L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_2, 
         L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_1, 
         L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_0, 
         L1_3_L2_2_G2_MINI_ALU_BoothXORCheck, 
         L1_3_L2_2_G2_MINI_ALU_BoothOperand_16, 
         L1_3_L2_2_G2_MINI_ALU_BoothOperand_15, 
         L1_3_L2_2_G2_MINI_ALU_BoothOperand_14, 
         L1_3_L2_2_G2_MINI_ALU_BoothOperand_13, 
         L1_3_L2_2_G2_MINI_ALU_BoothOperand_12, 
         L1_3_L2_2_G2_MINI_ALU_BoothOperand_11, 
         L1_3_L2_2_G2_MINI_ALU_BoothOperand_10, 
         L1_3_L2_2_G2_MINI_ALU_BoothOperand_9, L1_3_L2_2_G2_MINI_ALU_BoothP_16, 
         L1_3_L2_2_G2_MINI_ALU_BoothP_15, L1_3_L2_2_G2_MINI_ALU_BoothP_14, 
         L1_3_L2_2_G2_MINI_ALU_BoothP_13, L1_3_L2_2_G2_MINI_ALU_BoothP_12, 
         L1_3_L2_2_G2_MINI_ALU_BoothP_11, L1_3_L2_2_G2_MINI_ALU_BoothP_10, 
         L1_3_L2_2_G2_MINI_ALU_BoothP_9, L1_3_L2_2_G2_MINI_ALU_BoothP_8, 
         L1_3_L2_2_G2_MINI_ALU_BoothP_7, L1_3_L2_2_G2_MINI_ALU_BoothP_6, 
         L1_3_L2_2_G2_MINI_ALU_BoothP_5, L1_3_L2_2_G2_MINI_ALU_BoothP_4, 
         L1_3_L2_2_G2_MINI_ALU_BoothP_3, L1_3_L2_2_G2_MINI_ALU_BoothP_2, 
         L1_3_L2_2_G2_MINI_ALU_BoothP_1, L1_3_L2_2_G2_MINI_ALU_BoothP_0, 
         L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_15, 
         L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_14, 
         L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_13, 
         L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_12, 
         L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_11, 
         L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_10, 
         L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_9, 
         L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_8, 
         L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_7, 
         L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_6, 
         L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_5, 
         L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_4, 
         L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_3, 
         L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_2, 
         L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_1, 
         L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_0, 
         L1_3_L2_3_G2_MINI_ALU_BoothXORCheck, 
         L1_3_L2_3_G2_MINI_ALU_BoothOperand_16, 
         L1_3_L2_3_G2_MINI_ALU_BoothOperand_15, 
         L1_3_L2_3_G2_MINI_ALU_BoothOperand_14, 
         L1_3_L2_3_G2_MINI_ALU_BoothOperand_13, 
         L1_3_L2_3_G2_MINI_ALU_BoothOperand_12, 
         L1_3_L2_3_G2_MINI_ALU_BoothOperand_11, 
         L1_3_L2_3_G2_MINI_ALU_BoothOperand_10, 
         L1_3_L2_3_G2_MINI_ALU_BoothOperand_9, L1_3_L2_3_G2_MINI_ALU_BoothP_16, 
         L1_3_L2_3_G2_MINI_ALU_BoothP_15, L1_3_L2_3_G2_MINI_ALU_BoothP_14, 
         L1_3_L2_3_G2_MINI_ALU_BoothP_13, L1_3_L2_3_G2_MINI_ALU_BoothP_12, 
         L1_3_L2_3_G2_MINI_ALU_BoothP_11, L1_3_L2_3_G2_MINI_ALU_BoothP_10, 
         L1_3_L2_3_G2_MINI_ALU_BoothP_9, L1_3_L2_3_G2_MINI_ALU_BoothP_8, 
         L1_3_L2_3_G2_MINI_ALU_BoothP_7, L1_3_L2_3_G2_MINI_ALU_BoothP_6, 
         L1_3_L2_3_G2_MINI_ALU_BoothP_5, L1_3_L2_3_G2_MINI_ALU_BoothP_4, 
         L1_3_L2_3_G2_MINI_ALU_BoothP_3, L1_3_L2_3_G2_MINI_ALU_BoothP_2, 
         L1_3_L2_3_G2_MINI_ALU_BoothP_1, L1_3_L2_3_G2_MINI_ALU_BoothP_0, 
         L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_15, 
         L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_14, 
         L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_13, 
         L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_12, 
         L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_11, 
         L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_10, 
         L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_9, 
         L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_8, 
         L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_7, 
         L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_6, 
         L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_5, 
         L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_4, 
         L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_3, 
         L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_2, 
         L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_1, 
         L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_0, 
         L1_3_L2_4_G3_MINI_ALU_BoothXORCheck, 
         L1_3_L2_4_G3_MINI_ALU_BoothOperand_16, 
         L1_3_L2_4_G3_MINI_ALU_BoothOperand_15, 
         L1_3_L2_4_G3_MINI_ALU_BoothOperand_14, 
         L1_3_L2_4_G3_MINI_ALU_BoothOperand_13, 
         L1_3_L2_4_G3_MINI_ALU_BoothOperand_12, 
         L1_3_L2_4_G3_MINI_ALU_BoothOperand_11, 
         L1_3_L2_4_G3_MINI_ALU_BoothOperand_10, 
         L1_3_L2_4_G3_MINI_ALU_BoothOperand_9, L1_3_L2_4_G3_MINI_ALU_BoothP_16, 
         L1_3_L2_4_G3_MINI_ALU_BoothP_15, L1_3_L2_4_G3_MINI_ALU_BoothP_14, 
         L1_3_L2_4_G3_MINI_ALU_BoothP_13, L1_3_L2_4_G3_MINI_ALU_BoothP_12, 
         L1_3_L2_4_G3_MINI_ALU_BoothP_11, L1_3_L2_4_G3_MINI_ALU_BoothP_10, 
         L1_3_L2_4_G3_MINI_ALU_BoothP_9, L1_3_L2_4_G3_MINI_ALU_BoothP_8, 
         L1_3_L2_4_G3_MINI_ALU_BoothP_7, L1_3_L2_4_G3_MINI_ALU_BoothP_6, 
         L1_3_L2_4_G3_MINI_ALU_BoothP_5, L1_3_L2_4_G3_MINI_ALU_BoothP_4, 
         L1_3_L2_4_G3_MINI_ALU_BoothP_3, L1_3_L2_4_G3_MINI_ALU_BoothP_2, 
         L1_3_L2_4_G3_MINI_ALU_BoothP_1, L1_3_L2_4_G3_MINI_ALU_BoothP_0, 
         L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_15, 
         L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_14, 
         L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_13, 
         L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_12, 
         L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_11, 
         L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_10, 
         L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_9, 
         L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_8, 
         L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_7, 
         L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_6, 
         L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_5, 
         L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_4, 
         L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_3, 
         L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_2, 
         L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_1, 
         L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_0, 
         L1_4_L2_0_G3_MINI_ALU_BoothXORCheck, 
         L1_4_L2_0_G3_MINI_ALU_BoothOperand_16, 
         L1_4_L2_0_G3_MINI_ALU_BoothOperand_15, 
         L1_4_L2_0_G3_MINI_ALU_BoothOperand_14, 
         L1_4_L2_0_G3_MINI_ALU_BoothOperand_13, 
         L1_4_L2_0_G3_MINI_ALU_BoothOperand_12, 
         L1_4_L2_0_G3_MINI_ALU_BoothOperand_11, 
         L1_4_L2_0_G3_MINI_ALU_BoothOperand_10, 
         L1_4_L2_0_G3_MINI_ALU_BoothOperand_9, L1_4_L2_0_G3_MINI_ALU_BoothP_16, 
         L1_4_L2_0_G3_MINI_ALU_BoothP_15, L1_4_L2_0_G3_MINI_ALU_BoothP_14, 
         L1_4_L2_0_G3_MINI_ALU_BoothP_13, L1_4_L2_0_G3_MINI_ALU_BoothP_12, 
         L1_4_L2_0_G3_MINI_ALU_BoothP_11, L1_4_L2_0_G3_MINI_ALU_BoothP_10, 
         L1_4_L2_0_G3_MINI_ALU_BoothP_9, L1_4_L2_0_G3_MINI_ALU_BoothP_8, 
         L1_4_L2_0_G3_MINI_ALU_BoothP_7, L1_4_L2_0_G3_MINI_ALU_BoothP_6, 
         L1_4_L2_0_G3_MINI_ALU_BoothP_5, L1_4_L2_0_G3_MINI_ALU_BoothP_4, 
         L1_4_L2_0_G3_MINI_ALU_BoothP_3, L1_4_L2_0_G3_MINI_ALU_BoothP_2, 
         L1_4_L2_0_G3_MINI_ALU_BoothP_1, L1_4_L2_0_G3_MINI_ALU_BoothP_0, 
         L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_15, 
         L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_14, 
         L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_13, 
         L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_12, 
         L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_11, 
         L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_10, 
         L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_9, 
         L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_8, 
         L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_7, 
         L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_6, 
         L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_5, 
         L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_4, 
         L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_3, 
         L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_2, 
         L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_1, 
         L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_0, 
         L1_4_L2_1_G3_MINI_ALU_BoothXORCheck, 
         L1_4_L2_1_G3_MINI_ALU_BoothOperand_16, 
         L1_4_L2_1_G3_MINI_ALU_BoothOperand_15, 
         L1_4_L2_1_G3_MINI_ALU_BoothOperand_14, 
         L1_4_L2_1_G3_MINI_ALU_BoothOperand_13, 
         L1_4_L2_1_G3_MINI_ALU_BoothOperand_12, 
         L1_4_L2_1_G3_MINI_ALU_BoothOperand_11, 
         L1_4_L2_1_G3_MINI_ALU_BoothOperand_10, 
         L1_4_L2_1_G3_MINI_ALU_BoothOperand_9, L1_4_L2_1_G3_MINI_ALU_BoothP_16, 
         L1_4_L2_1_G3_MINI_ALU_BoothP_15, L1_4_L2_1_G3_MINI_ALU_BoothP_14, 
         L1_4_L2_1_G3_MINI_ALU_BoothP_13, L1_4_L2_1_G3_MINI_ALU_BoothP_12, 
         L1_4_L2_1_G3_MINI_ALU_BoothP_11, L1_4_L2_1_G3_MINI_ALU_BoothP_10, 
         L1_4_L2_1_G3_MINI_ALU_BoothP_9, L1_4_L2_1_G3_MINI_ALU_BoothP_8, 
         L1_4_L2_1_G3_MINI_ALU_BoothP_7, L1_4_L2_1_G3_MINI_ALU_BoothP_6, 
         L1_4_L2_1_G3_MINI_ALU_BoothP_5, L1_4_L2_1_G3_MINI_ALU_BoothP_4, 
         L1_4_L2_1_G3_MINI_ALU_BoothP_3, L1_4_L2_1_G3_MINI_ALU_BoothP_2, 
         L1_4_L2_1_G3_MINI_ALU_BoothP_1, L1_4_L2_1_G3_MINI_ALU_BoothP_0, 
         L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_15, 
         L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_14, 
         L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_13, 
         L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_12, 
         L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_11, 
         L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_10, 
         L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_9, 
         L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_8, 
         L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_7, 
         L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_6, 
         L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_5, 
         L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_4, 
         L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_3, 
         L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_2, 
         L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_1, 
         L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_0, 
         L1_4_L2_2_G4_MINI_ALU_BoothXORCheck, 
         L1_4_L2_2_G4_MINI_ALU_BoothOperand_16, 
         L1_4_L2_2_G4_MINI_ALU_BoothOperand_15, 
         L1_4_L2_2_G4_MINI_ALU_BoothOperand_14, 
         L1_4_L2_2_G4_MINI_ALU_BoothOperand_13, 
         L1_4_L2_2_G4_MINI_ALU_BoothOperand_12, 
         L1_4_L2_2_G4_MINI_ALU_BoothOperand_11, 
         L1_4_L2_2_G4_MINI_ALU_BoothOperand_10, 
         L1_4_L2_2_G4_MINI_ALU_BoothOperand_9, L1_4_L2_2_G4_MINI_ALU_BoothP_16, 
         L1_4_L2_2_G4_MINI_ALU_BoothP_15, L1_4_L2_2_G4_MINI_ALU_BoothP_14, 
         L1_4_L2_2_G4_MINI_ALU_BoothP_13, L1_4_L2_2_G4_MINI_ALU_BoothP_12, 
         L1_4_L2_2_G4_MINI_ALU_BoothP_11, L1_4_L2_2_G4_MINI_ALU_BoothP_10, 
         L1_4_L2_2_G4_MINI_ALU_BoothP_9, L1_4_L2_2_G4_MINI_ALU_BoothP_8, 
         L1_4_L2_2_G4_MINI_ALU_BoothP_7, L1_4_L2_2_G4_MINI_ALU_BoothP_6, 
         L1_4_L2_2_G4_MINI_ALU_BoothP_5, L1_4_L2_2_G4_MINI_ALU_BoothP_4, 
         L1_4_L2_2_G4_MINI_ALU_BoothP_3, L1_4_L2_2_G4_MINI_ALU_BoothP_2, 
         L1_4_L2_2_G4_MINI_ALU_BoothP_1, L1_4_L2_2_G4_MINI_ALU_BoothP_0, 
         L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_15, 
         L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_14, 
         L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_13, 
         L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_12, 
         L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_11, 
         L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_10, 
         L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_9, 
         L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_8, 
         L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_7, 
         L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_6, 
         L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_5, 
         L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_4, 
         L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_3, 
         L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_2, 
         L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_1, 
         L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_0, 
         L1_4_L2_3_G5_MINI_ALU_BoothXORCheck, 
         L1_4_L2_3_G5_MINI_ALU_BoothOperand_16, 
         L1_4_L2_3_G5_MINI_ALU_BoothOperand_15, 
         L1_4_L2_3_G5_MINI_ALU_BoothOperand_14, 
         L1_4_L2_3_G5_MINI_ALU_BoothOperand_13, 
         L1_4_L2_3_G5_MINI_ALU_BoothOperand_12, 
         L1_4_L2_3_G5_MINI_ALU_BoothOperand_11, 
         L1_4_L2_3_G5_MINI_ALU_BoothOperand_10, 
         L1_4_L2_3_G5_MINI_ALU_BoothOperand_9, L1_4_L2_3_G5_MINI_ALU_BoothP_16, 
         L1_4_L2_3_G5_MINI_ALU_BoothP_15, L1_4_L2_3_G5_MINI_ALU_BoothP_14, 
         L1_4_L2_3_G5_MINI_ALU_BoothP_13, L1_4_L2_3_G5_MINI_ALU_BoothP_12, 
         L1_4_L2_3_G5_MINI_ALU_BoothP_11, L1_4_L2_3_G5_MINI_ALU_BoothP_10, 
         L1_4_L2_3_G5_MINI_ALU_BoothP_9, L1_4_L2_3_G5_MINI_ALU_BoothP_8, 
         L1_4_L2_3_G5_MINI_ALU_BoothP_7, L1_4_L2_3_G5_MINI_ALU_BoothP_6, 
         L1_4_L2_3_G5_MINI_ALU_BoothP_5, L1_4_L2_3_G5_MINI_ALU_BoothP_4, 
         L1_4_L2_3_G5_MINI_ALU_BoothP_3, L1_4_L2_3_G5_MINI_ALU_BoothP_2, 
         L1_4_L2_3_G5_MINI_ALU_BoothP_1, L1_4_L2_3_G5_MINI_ALU_BoothP_0, 
         L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_15, 
         L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_14, 
         L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_13, 
         L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_12, 
         L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_11, 
         L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_10, 
         L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_9, 
         L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_8, 
         L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_7, 
         L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_6, 
         L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_5, 
         L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_4, 
         L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_3, 
         L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_2, 
         L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_1, 
         L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_0, 
         L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_7, 
         L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_6, 
         L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_5, 
         L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_4, 
         L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_3, 
         L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_2, 
         L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_1, 
         L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_0, 
         L1_4_L2_4_G5_MINI_ALU_OperationResult_15, 
         L1_4_L2_4_G5_MINI_ALU_OperationResult_14, 
         L1_4_L2_4_G5_MINI_ALU_OperationResult_13, 
         L1_4_L2_4_G5_MINI_ALU_OperationResult_12, 
         L1_4_L2_4_G5_MINI_ALU_OperationResult_11, 
         L1_4_L2_4_G5_MINI_ALU_OperationResult_10, 
         L1_4_L2_4_G5_MINI_ALU_OperationResult_9, 
         L1_4_L2_4_G5_MINI_ALU_OperationResult_8, 
         L1_4_L2_4_G5_MINI_ALU_OperationResult_7, 
         L1_4_L2_4_G5_MINI_ALU_OperationResult_6, 
         L1_4_L2_4_G5_MINI_ALU_OperationResult_5, 
         L1_4_L2_4_G5_MINI_ALU_OperationResult_4, 
         L1_4_L2_4_G5_MINI_ALU_OperationResult_3, 
         L1_4_L2_4_G5_MINI_ALU_OperationResult_2, 
         L1_4_L2_4_G5_MINI_ALU_OperationResult_1, 
         L1_4_L2_4_G5_MINI_ALU_OperationResult_0, 
         L1_4_L2_4_G5_MINI_ALU_BoothXORCheck, 
         L1_4_L2_4_G5_MINI_ALU_BoothOperand_16, 
         L1_4_L2_4_G5_MINI_ALU_BoothOperand_15, 
         L1_4_L2_4_G5_MINI_ALU_BoothOperand_14, 
         L1_4_L2_4_G5_MINI_ALU_BoothOperand_13, 
         L1_4_L2_4_G5_MINI_ALU_BoothOperand_12, 
         L1_4_L2_4_G5_MINI_ALU_BoothOperand_11, 
         L1_4_L2_4_G5_MINI_ALU_BoothOperand_10, 
         L1_4_L2_4_G5_MINI_ALU_BoothOperand_9, L1_4_L2_4_G5_MINI_ALU_BoothP_16, 
         L1_4_L2_4_G5_MINI_ALU_BoothP_15, L1_4_L2_4_G5_MINI_ALU_BoothP_14, 
         L1_4_L2_4_G5_MINI_ALU_BoothP_13, L1_4_L2_4_G5_MINI_ALU_BoothP_12, 
         L1_4_L2_4_G5_MINI_ALU_BoothP_11, L1_4_L2_4_G5_MINI_ALU_BoothP_10, 
         L1_4_L2_4_G5_MINI_ALU_BoothP_9, L1_4_L2_4_G5_MINI_ALU_BoothP_8, 
         L1_4_L2_4_G5_MINI_ALU_BoothP_7, L1_4_L2_4_G5_MINI_ALU_BoothP_6, 
         L1_4_L2_4_G5_MINI_ALU_BoothP_5, L1_4_L2_4_G5_MINI_ALU_BoothP_4, 
         L1_4_L2_4_G5_MINI_ALU_BoothP_3, L1_4_L2_4_G5_MINI_ALU_BoothP_2, 
         L1_4_L2_4_G5_MINI_ALU_BoothP_1, L1_4_L2_4_G5_MINI_ALU_BoothP_0, 
         L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_15, 
         L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_14, 
         L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_13, 
         L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_12, 
         L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_11, 
         L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_10, 
         L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_9, 
         L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_8, 
         L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_7, 
         L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_6, 
         L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_5, 
         L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_4, 
         L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_3, 
         L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_2, 
         L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_1, 
         L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_0, L1FirstOperands_12__16, nx22, 
         CounterOut_0, NOT__145383, nx1032, NOT_CounterOut_0, nx1036, 
         CounterOut_3, CounterOut_2, CounterOut_1, nx1046, nx1058, nx1066, 
         nx2853, nx2865, nx2869, nx2873, nx3230, nx3233, nx3235, nx3239, nx3241, 
         nx3244, nx3246, nx3270, nx3272, nx3274, nx3276, nx3278, nx3280, nx3282, 
         nx3284, nx3286, nx3292;
    wire [903:0] \$dummy ;




    booth_adder_17 L1_0_L2_0_G1_MINI_ALU_BOOTH_ADDER (.AdderFirstOperand ({
                   L1FirstOperands_12__16,L1FirstOperands_0__15,
                   L1FirstOperands_0__14,L1FirstOperands_0__13,
                   L1FirstOperands_0__12,L1FirstOperands_0__11,
                   L1FirstOperands_0__10,L1FirstOperands_0__9,
                   L1FirstOperands_0__8,L1FirstOperands_0__7,
                   L1FirstOperands_0__6,L1FirstOperands_0__5,
                   L1FirstOperands_0__4,L1FirstOperands_0__3,
                   L1FirstOperands_0__2,L1FirstOperands_0__1,
                   L1FirstOperands_0__0}), .AdderSecondOperand ({
                   L1FirstOperands_12__16,
                   L1_0_L2_0_G1_MINI_ALU_OperationResult_15,
                   L1_0_L2_0_G1_MINI_ALU_OperationResult_14,
                   L1_0_L2_0_G1_MINI_ALU_OperationResult_13,
                   L1_0_L2_0_G1_MINI_ALU_OperationResult_12,
                   L1_0_L2_0_G1_MINI_ALU_OperationResult_11,
                   L1_0_L2_0_G1_MINI_ALU_OperationResult_10,
                   L1_0_L2_0_G1_MINI_ALU_OperationResult_9,
                   L1_0_L2_0_G1_MINI_ALU_OperationResult_8,
                   L1_0_L2_0_G1_MINI_ALU_OperationResult_7,
                   L1_0_L2_0_G1_MINI_ALU_OperationResult_6,
                   L1_0_L2_0_G1_MINI_ALU_OperationResult_5,
                   L1_0_L2_0_G1_MINI_ALU_OperationResult_4,
                   L1_0_L2_0_G1_MINI_ALU_OperationResult_3,
                   L1_0_L2_0_G1_MINI_ALU_OperationResult_2,
                   L1_0_L2_0_G1_MINI_ALU_OperationResult_1,
                   L1_0_L2_0_G1_MINI_ALU_OperationResult_0}), .BoothOperand ({
                   L1_0_L2_0_G1_MINI_ALU_BoothOperand_16,
                   L1_0_L2_0_G1_MINI_ALU_BoothOperand_15,
                   L1_0_L2_0_G1_MINI_ALU_BoothOperand_14,
                   L1_0_L2_0_G1_MINI_ALU_BoothOperand_13,
                   L1_0_L2_0_G1_MINI_ALU_BoothOperand_12,
                   L1_0_L2_0_G1_MINI_ALU_BoothOperand_11,
                   L1_0_L2_0_G1_MINI_ALU_BoothOperand_10,
                   L1_0_L2_0_G1_MINI_ALU_BoothOperand_9,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16}), .BoothP ({
                   L1_0_L2_0_G1_MINI_ALU_BoothP_16,
                   L1_0_L2_0_G1_MINI_ALU_BoothP_15,
                   L1_0_L2_0_G1_MINI_ALU_BoothP_14,
                   L1_0_L2_0_G1_MINI_ALU_BoothP_13,
                   L1_0_L2_0_G1_MINI_ALU_BoothP_12,
                   L1_0_L2_0_G1_MINI_ALU_BoothP_11,
                   L1_0_L2_0_G1_MINI_ALU_BoothP_10,
                   L1_0_L2_0_G1_MINI_ALU_BoothP_9,L1_0_L2_0_G1_MINI_ALU_BoothP_8
                   ,L1_0_L2_0_G1_MINI_ALU_BoothP_7,
                   L1_0_L2_0_G1_MINI_ALU_BoothP_6,L1_0_L2_0_G1_MINI_ALU_BoothP_5
                   ,L1_0_L2_0_G1_MINI_ALU_BoothP_4,
                   L1_0_L2_0_G1_MINI_ALU_BoothP_3,L1_0_L2_0_G1_MINI_ALU_BoothP_2
                   ,L1_0_L2_0_G1_MINI_ALU_BoothP_1,
                   L1_0_L2_0_G1_MINI_ALU_BoothP_0}), .SelOperand (nx3282), .Operation (
                   L1_0_L2_0_G1_MINI_ALU_BoothXORCheck), .AdderResult ({
                   L1ResultsLarge_0__16,L1ResultsLarge_0__15,
                   L1ResultsLarge_0__14,L1ResultsLarge_0__13,
                   L1ResultsLarge_0__12,L1ResultsLarge_0__11,
                   L1ResultsLarge_0__10,L1ResultsLarge_0__9,L1ResultsLarge_0__8,
                   L1ResultsLarge_0__7,L1ResultsLarge_0__6,L1ResultsLarge_0__5,
                   L1ResultsLarge_0__4,L1ResultsLarge_0__3,L1ResultsLarge_0__2,
                   L1ResultsLarge_0__1,L1ResultsLarge_0__0}), .AdderBoothResult (
                   {\$dummy [0],L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_15,
                   L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_14,
                   L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_13,
                   L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_12,
                   L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_11,
                   L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_10,
                   L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_9,
                   L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_8,
                   L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_7,
                   L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_6,
                   L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_5,
                   L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_4,
                   L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_3,
                   L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_2,
                   L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_1,
                   L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_0})) ;
    booth_unit_17 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT (.CLK (CLK), .RST (RST), .Start (
                  Start), .Instr (Instr), .LoopingAndResultNotReady (nx3272), .Filter (
                  {FilterDin_0__0__7,FilterDin_0__0__6,FilterDin_0__0__5,
                  FilterDin_0__0__4,FilterDin_0__0__3,FilterDin_0__0__2,
                  FilterDin_0__0__1,FilterDin_0__0__0}), .Window ({
                  WindowDin_0__0__7,WindowDin_0__0__6,WindowDin_0__0__5,
                  WindowDin_0__0__4,WindowDin_0__0__3,WindowDin_0__0__2,
                  WindowDin_0__0__1,WindowDin_0__0__0}), .AdderBoothResult ({
                  L1FirstOperands_12__16,
                  L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_15,
                  L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_14,
                  L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_13,
                  L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_12,
                  L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_11,
                  L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_10,
                  L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_9,
                  L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_8,
                  L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_7,
                  L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_6,
                  L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_5,
                  L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_4,
                  L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_3,
                  L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_2,
                  L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_1,
                  L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_0}), .BoothXORCheck (
                  L1_0_L2_0_G1_MINI_ALU_BoothXORCheck), .BoothResult ({
                  \$dummy [1],\$dummy [2],\$dummy [3],\$dummy [4],\$dummy [5],
                  \$dummy [6],\$dummy [7],\$dummy [8]}), .BoothAddingOperand ({
                  L1_0_L2_0_G1_MINI_ALU_BoothOperand_16,
                  L1_0_L2_0_G1_MINI_ALU_BoothOperand_15,
                  L1_0_L2_0_G1_MINI_ALU_BoothOperand_14,
                  L1_0_L2_0_G1_MINI_ALU_BoothOperand_13,
                  L1_0_L2_0_G1_MINI_ALU_BoothOperand_12,
                  L1_0_L2_0_G1_MINI_ALU_BoothOperand_11,
                  L1_0_L2_0_G1_MINI_ALU_BoothOperand_10,
                  L1_0_L2_0_G1_MINI_ALU_BoothOperand_9,\$dummy [9],\$dummy [10],
                  \$dummy [11],\$dummy [12],\$dummy [13],\$dummy [14],
                  \$dummy [15],\$dummy [16],\$dummy [17]}), .BoothP ({
                  L1_0_L2_0_G1_MINI_ALU_BoothP_16,
                  L1_0_L2_0_G1_MINI_ALU_BoothP_15,
                  L1_0_L2_0_G1_MINI_ALU_BoothP_14,
                  L1_0_L2_0_G1_MINI_ALU_BoothP_13,
                  L1_0_L2_0_G1_MINI_ALU_BoothP_12,
                  L1_0_L2_0_G1_MINI_ALU_BoothP_11,
                  L1_0_L2_0_G1_MINI_ALU_BoothP_10,L1_0_L2_0_G1_MINI_ALU_BoothP_9
                  ,L1_0_L2_0_G1_MINI_ALU_BoothP_8,L1_0_L2_0_G1_MINI_ALU_BoothP_7
                  ,L1_0_L2_0_G1_MINI_ALU_BoothP_6,L1_0_L2_0_G1_MINI_ALU_BoothP_5
                  ,L1_0_L2_0_G1_MINI_ALU_BoothP_4,L1_0_L2_0_G1_MINI_ALU_BoothP_3
                  ,L1_0_L2_0_G1_MINI_ALU_BoothP_2,L1_0_L2_0_G1_MINI_ALU_BoothP_1
                  ,L1_0_L2_0_G1_MINI_ALU_BoothP_0}), .LargeWindowShifted ({
                  \$dummy [18],\$dummy [19],\$dummy [20],\$dummy [21],
                  \$dummy [22],\$dummy [23],\$dummy [24],\$dummy [25],
                  \$dummy [26],\$dummy [27],\$dummy [28],\$dummy [29],
                  \$dummy [30],\$dummy [31],\$dummy [32],\$dummy [33],
                  \$dummy [34]})) ;
    booth_adder_17 L1_0_L2_1_G1_MINI_ALU_BOOTH_ADDER (.AdderFirstOperand ({
                   L1FirstOperands_12__16,L1FirstOperands_0__15,
                   L1FirstOperands_0__14,L1FirstOperands_0__13,
                   L1FirstOperands_0__12,L1FirstOperands_0__11,
                   L1FirstOperands_0__10,L1FirstOperands_0__9,
                   L1FirstOperands_0__8,L1FirstOperands_0__7,
                   L1FirstOperands_0__6,L1FirstOperands_0__5,
                   L1FirstOperands_0__4,L1FirstOperands_0__3,
                   L1FirstOperands_0__2,L1FirstOperands_0__1,
                   L1FirstOperands_0__0}), .AdderSecondOperand ({
                   L1FirstOperands_12__16,
                   L1_0_L2_1_G1_MINI_ALU_OperationResult_15,
                   L1_0_L2_1_G1_MINI_ALU_OperationResult_14,
                   L1_0_L2_1_G1_MINI_ALU_OperationResult_13,
                   L1_0_L2_1_G1_MINI_ALU_OperationResult_12,
                   L1_0_L2_1_G1_MINI_ALU_OperationResult_11,
                   L1_0_L2_1_G1_MINI_ALU_OperationResult_10,
                   L1_0_L2_1_G1_MINI_ALU_OperationResult_9,
                   L1_0_L2_1_G1_MINI_ALU_OperationResult_8,
                   L1_0_L2_1_G1_MINI_ALU_OperationResult_7,
                   L1_0_L2_1_G1_MINI_ALU_OperationResult_6,
                   L1_0_L2_1_G1_MINI_ALU_OperationResult_5,
                   L1_0_L2_1_G1_MINI_ALU_OperationResult_4,
                   L1_0_L2_1_G1_MINI_ALU_OperationResult_3,
                   L1_0_L2_1_G1_MINI_ALU_OperationResult_2,
                   L1_0_L2_1_G1_MINI_ALU_OperationResult_1,
                   L1_0_L2_1_G1_MINI_ALU_OperationResult_0}), .BoothOperand ({
                   L1_0_L2_1_G1_MINI_ALU_BoothOperand_16,
                   L1_0_L2_1_G1_MINI_ALU_BoothOperand_15,
                   L1_0_L2_1_G1_MINI_ALU_BoothOperand_14,
                   L1_0_L2_1_G1_MINI_ALU_BoothOperand_13,
                   L1_0_L2_1_G1_MINI_ALU_BoothOperand_12,
                   L1_0_L2_1_G1_MINI_ALU_BoothOperand_11,
                   L1_0_L2_1_G1_MINI_ALU_BoothOperand_10,
                   L1_0_L2_1_G1_MINI_ALU_BoothOperand_9,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16}), .BoothP ({
                   L1_0_L2_1_G1_MINI_ALU_BoothP_16,
                   L1_0_L2_1_G1_MINI_ALU_BoothP_15,
                   L1_0_L2_1_G1_MINI_ALU_BoothP_14,
                   L1_0_L2_1_G1_MINI_ALU_BoothP_13,
                   L1_0_L2_1_G1_MINI_ALU_BoothP_12,
                   L1_0_L2_1_G1_MINI_ALU_BoothP_11,
                   L1_0_L2_1_G1_MINI_ALU_BoothP_10,
                   L1_0_L2_1_G1_MINI_ALU_BoothP_9,L1_0_L2_1_G1_MINI_ALU_BoothP_8
                   ,L1_0_L2_1_G1_MINI_ALU_BoothP_7,
                   L1_0_L2_1_G1_MINI_ALU_BoothP_6,L1_0_L2_1_G1_MINI_ALU_BoothP_5
                   ,L1_0_L2_1_G1_MINI_ALU_BoothP_4,
                   L1_0_L2_1_G1_MINI_ALU_BoothP_3,L1_0_L2_1_G1_MINI_ALU_BoothP_2
                   ,L1_0_L2_1_G1_MINI_ALU_BoothP_1,
                   L1_0_L2_1_G1_MINI_ALU_BoothP_0}), .SelOperand (nx3282), .Operation (
                   L1_0_L2_1_G1_MINI_ALU_BoothXORCheck), .AdderResult ({
                   L1ResultsLarge_1__16,L1ResultsLarge_1__15,
                   L1ResultsLarge_1__14,L1ResultsLarge_1__13,
                   L1ResultsLarge_1__12,L1ResultsLarge_1__11,
                   L1ResultsLarge_1__10,L1ResultsLarge_1__9,L1ResultsLarge_1__8,
                   L1ResultsLarge_1__7,L1ResultsLarge_1__6,L1ResultsLarge_1__5,
                   L1ResultsLarge_1__4,L1ResultsLarge_1__3,L1ResultsLarge_1__2,
                   L1ResultsLarge_1__1,L1ResultsLarge_1__0}), .AdderBoothResult (
                   {\$dummy [35],L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_15,
                   L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_14,
                   L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_13,
                   L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_12,
                   L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_11,
                   L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_10,
                   L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_9,
                   L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_8,
                   L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_7,
                   L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_6,
                   L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_5,
                   L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_4,
                   L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_3,
                   L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_2,
                   L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_1,
                   L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_0})) ;
    booth_unit_17 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT (.CLK (CLK), .RST (RST), .Start (
                  Start), .Instr (Instr), .LoopingAndResultNotReady (nx3272), .Filter (
                  {FilterDin_0__1__7,FilterDin_0__1__6,FilterDin_0__1__5,
                  FilterDin_0__1__4,FilterDin_0__1__3,FilterDin_0__1__2,
                  FilterDin_0__1__1,FilterDin_0__1__0}), .Window ({
                  WindowDin_0__1__7,WindowDin_0__1__6,WindowDin_0__1__5,
                  WindowDin_0__1__4,WindowDin_0__1__3,WindowDin_0__1__2,
                  WindowDin_0__1__1,WindowDin_0__1__0}), .AdderBoothResult ({
                  L1FirstOperands_12__16,
                  L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_15,
                  L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_14,
                  L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_13,
                  L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_12,
                  L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_11,
                  L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_10,
                  L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_9,
                  L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_8,
                  L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_7,
                  L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_6,
                  L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_5,
                  L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_4,
                  L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_3,
                  L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_2,
                  L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_1,
                  L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_0}), .BoothXORCheck (
                  L1_0_L2_1_G1_MINI_ALU_BoothXORCheck), .BoothResult ({
                  \$dummy [36],\$dummy [37],\$dummy [38],\$dummy [39],
                  \$dummy [40],\$dummy [41],\$dummy [42],\$dummy [43]}), .BoothAddingOperand (
                  {L1_0_L2_1_G1_MINI_ALU_BoothOperand_16,
                  L1_0_L2_1_G1_MINI_ALU_BoothOperand_15,
                  L1_0_L2_1_G1_MINI_ALU_BoothOperand_14,
                  L1_0_L2_1_G1_MINI_ALU_BoothOperand_13,
                  L1_0_L2_1_G1_MINI_ALU_BoothOperand_12,
                  L1_0_L2_1_G1_MINI_ALU_BoothOperand_11,
                  L1_0_L2_1_G1_MINI_ALU_BoothOperand_10,
                  L1_0_L2_1_G1_MINI_ALU_BoothOperand_9,\$dummy [44],\$dummy [45]
                  ,\$dummy [46],\$dummy [47],\$dummy [48],\$dummy [49],
                  \$dummy [50],\$dummy [51],\$dummy [52]}), .BoothP ({
                  L1_0_L2_1_G1_MINI_ALU_BoothP_16,
                  L1_0_L2_1_G1_MINI_ALU_BoothP_15,
                  L1_0_L2_1_G1_MINI_ALU_BoothP_14,
                  L1_0_L2_1_G1_MINI_ALU_BoothP_13,
                  L1_0_L2_1_G1_MINI_ALU_BoothP_12,
                  L1_0_L2_1_G1_MINI_ALU_BoothP_11,
                  L1_0_L2_1_G1_MINI_ALU_BoothP_10,L1_0_L2_1_G1_MINI_ALU_BoothP_9
                  ,L1_0_L2_1_G1_MINI_ALU_BoothP_8,L1_0_L2_1_G1_MINI_ALU_BoothP_7
                  ,L1_0_L2_1_G1_MINI_ALU_BoothP_6,L1_0_L2_1_G1_MINI_ALU_BoothP_5
                  ,L1_0_L2_1_G1_MINI_ALU_BoothP_4,L1_0_L2_1_G1_MINI_ALU_BoothP_3
                  ,L1_0_L2_1_G1_MINI_ALU_BoothP_2,L1_0_L2_1_G1_MINI_ALU_BoothP_1
                  ,L1_0_L2_1_G1_MINI_ALU_BoothP_0}), .LargeWindowShifted ({
                  \$dummy [53],\$dummy [54],\$dummy [55],\$dummy [56],
                  \$dummy [57],\$dummy [58],\$dummy [59],\$dummy [60],
                  \$dummy [61],\$dummy [62],\$dummy [63],\$dummy [64],
                  \$dummy [65],\$dummy [66],\$dummy [67],\$dummy [68],
                  \$dummy [69]})) ;
    booth_adder_17 L1_0_L2_2_G1_MINI_ALU_BOOTH_ADDER (.AdderFirstOperand ({
                   L1FirstOperands_12__16,L1FirstOperands_2__15,
                   L1FirstOperands_2__14,L1FirstOperands_2__13,
                   L1FirstOperands_2__12,L1FirstOperands_2__11,
                   L1FirstOperands_2__10,L1FirstOperands_2__9,
                   L1FirstOperands_2__8,L1FirstOperands_2__7,
                   L1FirstOperands_2__6,L1FirstOperands_2__5,
                   L1FirstOperands_2__4,L1FirstOperands_2__3,
                   L1FirstOperands_2__2,L1FirstOperands_2__1,
                   L1FirstOperands_2__0}), .AdderSecondOperand ({
                   L1FirstOperands_12__16,
                   L1_0_L2_2_G1_MINI_ALU_OperationResult_15,
                   L1_0_L2_2_G1_MINI_ALU_OperationResult_14,
                   L1_0_L2_2_G1_MINI_ALU_OperationResult_13,
                   L1_0_L2_2_G1_MINI_ALU_OperationResult_12,
                   L1_0_L2_2_G1_MINI_ALU_OperationResult_11,
                   L1_0_L2_2_G1_MINI_ALU_OperationResult_10,
                   L1_0_L2_2_G1_MINI_ALU_OperationResult_9,
                   L1_0_L2_2_G1_MINI_ALU_OperationResult_8,
                   L1_0_L2_2_G1_MINI_ALU_OperationResult_7,
                   L1_0_L2_2_G1_MINI_ALU_OperationResult_6,
                   L1_0_L2_2_G1_MINI_ALU_OperationResult_5,
                   L1_0_L2_2_G1_MINI_ALU_OperationResult_4,
                   L1_0_L2_2_G1_MINI_ALU_OperationResult_3,
                   L1_0_L2_2_G1_MINI_ALU_OperationResult_2,
                   L1_0_L2_2_G1_MINI_ALU_OperationResult_1,
                   L1_0_L2_2_G1_MINI_ALU_OperationResult_0}), .BoothOperand ({
                   L1_0_L2_2_G1_MINI_ALU_BoothOperand_16,
                   L1_0_L2_2_G1_MINI_ALU_BoothOperand_15,
                   L1_0_L2_2_G1_MINI_ALU_BoothOperand_14,
                   L1_0_L2_2_G1_MINI_ALU_BoothOperand_13,
                   L1_0_L2_2_G1_MINI_ALU_BoothOperand_12,
                   L1_0_L2_2_G1_MINI_ALU_BoothOperand_11,
                   L1_0_L2_2_G1_MINI_ALU_BoothOperand_10,
                   L1_0_L2_2_G1_MINI_ALU_BoothOperand_9,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16}), .BoothP ({
                   L1_0_L2_2_G1_MINI_ALU_BoothP_16,
                   L1_0_L2_2_G1_MINI_ALU_BoothP_15,
                   L1_0_L2_2_G1_MINI_ALU_BoothP_14,
                   L1_0_L2_2_G1_MINI_ALU_BoothP_13,
                   L1_0_L2_2_G1_MINI_ALU_BoothP_12,
                   L1_0_L2_2_G1_MINI_ALU_BoothP_11,
                   L1_0_L2_2_G1_MINI_ALU_BoothP_10,
                   L1_0_L2_2_G1_MINI_ALU_BoothP_9,L1_0_L2_2_G1_MINI_ALU_BoothP_8
                   ,L1_0_L2_2_G1_MINI_ALU_BoothP_7,
                   L1_0_L2_2_G1_MINI_ALU_BoothP_6,L1_0_L2_2_G1_MINI_ALU_BoothP_5
                   ,L1_0_L2_2_G1_MINI_ALU_BoothP_4,
                   L1_0_L2_2_G1_MINI_ALU_BoothP_3,L1_0_L2_2_G1_MINI_ALU_BoothP_2
                   ,L1_0_L2_2_G1_MINI_ALU_BoothP_1,
                   L1_0_L2_2_G1_MINI_ALU_BoothP_0}), .SelOperand (nx3280), .Operation (
                   L1_0_L2_2_G1_MINI_ALU_BoothXORCheck), .AdderResult ({
                   L1ResultsLarge_2__16,L1ResultsLarge_2__15,
                   L1ResultsLarge_2__14,L1ResultsLarge_2__13,
                   L1ResultsLarge_2__12,L1ResultsLarge_2__11,
                   L1ResultsLarge_2__10,L1ResultsLarge_2__9,L1ResultsLarge_2__8,
                   L1ResultsLarge_2__7,L1ResultsLarge_2__6,L1ResultsLarge_2__5,
                   L1ResultsLarge_2__4,L1ResultsLarge_2__3,L1ResultsLarge_2__2,
                   L1ResultsLarge_2__1,L1ResultsLarge_2__0}), .AdderBoothResult (
                   {\$dummy [70],L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_15,
                   L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_14,
                   L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_13,
                   L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_12,
                   L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_11,
                   L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_10,
                   L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_9,
                   L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_8,
                   L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_7,
                   L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_6,
                   L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_5,
                   L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_4,
                   L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_3,
                   L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_2,
                   L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_1,
                   L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_0})) ;
    booth_unit_17 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT (.CLK (CLK), .RST (RST), .Start (
                  Start), .Instr (Instr), .LoopingAndResultNotReady (nx3272), .Filter (
                  {FilterDin_0__2__7,FilterDin_0__2__6,FilterDin_0__2__5,
                  FilterDin_0__2__4,FilterDin_0__2__3,FilterDin_0__2__2,
                  FilterDin_0__2__1,FilterDin_0__2__0}), .Window ({
                  WindowDin_0__2__7,WindowDin_0__2__6,WindowDin_0__2__5,
                  WindowDin_0__2__4,WindowDin_0__2__3,WindowDin_0__2__2,
                  WindowDin_0__2__1,WindowDin_0__2__0}), .AdderBoothResult ({
                  L1FirstOperands_12__16,
                  L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_15,
                  L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_14,
                  L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_13,
                  L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_12,
                  L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_11,
                  L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_10,
                  L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_9,
                  L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_8,
                  L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_7,
                  L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_6,
                  L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_5,
                  L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_4,
                  L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_3,
                  L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_2,
                  L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_1,
                  L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_0}), .BoothXORCheck (
                  L1_0_L2_2_G1_MINI_ALU_BoothXORCheck), .BoothResult ({
                  \$dummy [71],\$dummy [72],\$dummy [73],\$dummy [74],
                  \$dummy [75],\$dummy [76],\$dummy [77],\$dummy [78]}), .BoothAddingOperand (
                  {L1_0_L2_2_G1_MINI_ALU_BoothOperand_16,
                  L1_0_L2_2_G1_MINI_ALU_BoothOperand_15,
                  L1_0_L2_2_G1_MINI_ALU_BoothOperand_14,
                  L1_0_L2_2_G1_MINI_ALU_BoothOperand_13,
                  L1_0_L2_2_G1_MINI_ALU_BoothOperand_12,
                  L1_0_L2_2_G1_MINI_ALU_BoothOperand_11,
                  L1_0_L2_2_G1_MINI_ALU_BoothOperand_10,
                  L1_0_L2_2_G1_MINI_ALU_BoothOperand_9,\$dummy [79],\$dummy [80]
                  ,\$dummy [81],\$dummy [82],\$dummy [83],\$dummy [84],
                  \$dummy [85],\$dummy [86],\$dummy [87]}), .BoothP ({
                  L1_0_L2_2_G1_MINI_ALU_BoothP_16,
                  L1_0_L2_2_G1_MINI_ALU_BoothP_15,
                  L1_0_L2_2_G1_MINI_ALU_BoothP_14,
                  L1_0_L2_2_G1_MINI_ALU_BoothP_13,
                  L1_0_L2_2_G1_MINI_ALU_BoothP_12,
                  L1_0_L2_2_G1_MINI_ALU_BoothP_11,
                  L1_0_L2_2_G1_MINI_ALU_BoothP_10,L1_0_L2_2_G1_MINI_ALU_BoothP_9
                  ,L1_0_L2_2_G1_MINI_ALU_BoothP_8,L1_0_L2_2_G1_MINI_ALU_BoothP_7
                  ,L1_0_L2_2_G1_MINI_ALU_BoothP_6,L1_0_L2_2_G1_MINI_ALU_BoothP_5
                  ,L1_0_L2_2_G1_MINI_ALU_BoothP_4,L1_0_L2_2_G1_MINI_ALU_BoothP_3
                  ,L1_0_L2_2_G1_MINI_ALU_BoothP_2,L1_0_L2_2_G1_MINI_ALU_BoothP_1
                  ,L1_0_L2_2_G1_MINI_ALU_BoothP_0}), .LargeWindowShifted ({
                  \$dummy [88],\$dummy [89],\$dummy [90],\$dummy [91],
                  \$dummy [92],\$dummy [93],\$dummy [94],\$dummy [95],
                  \$dummy [96],\$dummy [97],\$dummy [98],\$dummy [99],
                  \$dummy [100],\$dummy [101],\$dummy [102],\$dummy [103],
                  \$dummy [104]})) ;
    booth_adder_17 L1_0_L2_3_G1_MINI_ALU_BOOTH_ADDER (.AdderFirstOperand ({
                   L1FirstOperands_12__16,L1FirstOperands_3__15,
                   L1FirstOperands_3__14,L1FirstOperands_3__13,
                   L1FirstOperands_3__12,L1FirstOperands_3__11,
                   L1FirstOperands_3__10,L1FirstOperands_3__9,
                   L1FirstOperands_3__8,L1FirstOperands_3__7,
                   L1FirstOperands_3__6,L1FirstOperands_3__5,
                   L1FirstOperands_3__4,L1FirstOperands_3__3,
                   L1FirstOperands_3__2,L1FirstOperands_3__1,
                   L1FirstOperands_3__0}), .AdderSecondOperand ({
                   L1FirstOperands_12__16,
                   L1_0_L2_3_G1_MINI_ALU_OperationResult_15,
                   L1_0_L2_3_G1_MINI_ALU_OperationResult_14,
                   L1_0_L2_3_G1_MINI_ALU_OperationResult_13,
                   L1_0_L2_3_G1_MINI_ALU_OperationResult_12,
                   L1_0_L2_3_G1_MINI_ALU_OperationResult_11,
                   L1_0_L2_3_G1_MINI_ALU_OperationResult_10,
                   L1_0_L2_3_G1_MINI_ALU_OperationResult_9,
                   L1_0_L2_3_G1_MINI_ALU_OperationResult_8,
                   L1_0_L2_3_G1_MINI_ALU_OperationResult_7,
                   L1_0_L2_3_G1_MINI_ALU_OperationResult_6,
                   L1_0_L2_3_G1_MINI_ALU_OperationResult_5,
                   L1_0_L2_3_G1_MINI_ALU_OperationResult_4,
                   L1_0_L2_3_G1_MINI_ALU_OperationResult_3,
                   L1_0_L2_3_G1_MINI_ALU_OperationResult_2,
                   L1_0_L2_3_G1_MINI_ALU_OperationResult_1,
                   L1_0_L2_3_G1_MINI_ALU_OperationResult_0}), .BoothOperand ({
                   L1_0_L2_3_G1_MINI_ALU_BoothOperand_16,
                   L1_0_L2_3_G1_MINI_ALU_BoothOperand_15,
                   L1_0_L2_3_G1_MINI_ALU_BoothOperand_14,
                   L1_0_L2_3_G1_MINI_ALU_BoothOperand_13,
                   L1_0_L2_3_G1_MINI_ALU_BoothOperand_12,
                   L1_0_L2_3_G1_MINI_ALU_BoothOperand_11,
                   L1_0_L2_3_G1_MINI_ALU_BoothOperand_10,
                   L1_0_L2_3_G1_MINI_ALU_BoothOperand_9,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16}), .BoothP ({
                   L1_0_L2_3_G1_MINI_ALU_BoothP_16,
                   L1_0_L2_3_G1_MINI_ALU_BoothP_15,
                   L1_0_L2_3_G1_MINI_ALU_BoothP_14,
                   L1_0_L2_3_G1_MINI_ALU_BoothP_13,
                   L1_0_L2_3_G1_MINI_ALU_BoothP_12,
                   L1_0_L2_3_G1_MINI_ALU_BoothP_11,
                   L1_0_L2_3_G1_MINI_ALU_BoothP_10,
                   L1_0_L2_3_G1_MINI_ALU_BoothP_9,L1_0_L2_3_G1_MINI_ALU_BoothP_8
                   ,L1_0_L2_3_G1_MINI_ALU_BoothP_7,
                   L1_0_L2_3_G1_MINI_ALU_BoothP_6,L1_0_L2_3_G1_MINI_ALU_BoothP_5
                   ,L1_0_L2_3_G1_MINI_ALU_BoothP_4,
                   L1_0_L2_3_G1_MINI_ALU_BoothP_3,L1_0_L2_3_G1_MINI_ALU_BoothP_2
                   ,L1_0_L2_3_G1_MINI_ALU_BoothP_1,
                   L1_0_L2_3_G1_MINI_ALU_BoothP_0}), .SelOperand (nx3280), .Operation (
                   L1_0_L2_3_G1_MINI_ALU_BoothXORCheck), .AdderResult ({
                   L1ResultsLarge_3__16,L1ResultsLarge_3__15,
                   L1ResultsLarge_3__14,L1ResultsLarge_3__13,
                   L1ResultsLarge_3__12,L1ResultsLarge_3__11,
                   L1ResultsLarge_3__10,L1ResultsLarge_3__9,L1ResultsLarge_3__8,
                   L1ResultsLarge_3__7,L1ResultsLarge_3__6,L1ResultsLarge_3__5,
                   L1ResultsLarge_3__4,L1ResultsLarge_3__3,L1ResultsLarge_3__2,
                   L1ResultsLarge_3__1,L1ResultsLarge_3__0}), .AdderBoothResult (
                   {\$dummy [105],L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_15,
                   L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_14,
                   L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_13,
                   L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_12,
                   L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_11,
                   L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_10,
                   L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_9,
                   L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_8,
                   L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_7,
                   L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_6,
                   L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_5,
                   L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_4,
                   L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_3,
                   L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_2,
                   L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_1,
                   L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_0})) ;
    booth_unit_17 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT (.CLK (CLK), .RST (RST), .Start (
                  Start), .Instr (Instr), .LoopingAndResultNotReady (nx3272), .Filter (
                  {FilterDin_0__3__7,FilterDin_0__3__6,FilterDin_0__3__5,
                  FilterDin_0__3__4,FilterDin_0__3__3,FilterDin_0__3__2,
                  FilterDin_0__3__1,FilterDin_0__3__0}), .Window ({
                  WindowDin_0__3__7,WindowDin_0__3__6,WindowDin_0__3__5,
                  WindowDin_0__3__4,WindowDin_0__3__3,WindowDin_0__3__2,
                  WindowDin_0__3__1,WindowDin_0__3__0}), .AdderBoothResult ({
                  L1FirstOperands_12__16,
                  L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_15,
                  L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_14,
                  L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_13,
                  L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_12,
                  L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_11,
                  L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_10,
                  L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_9,
                  L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_8,
                  L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_7,
                  L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_6,
                  L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_5,
                  L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_4,
                  L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_3,
                  L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_2,
                  L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_1,
                  L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_0}), .BoothXORCheck (
                  L1_0_L2_3_G1_MINI_ALU_BoothXORCheck), .BoothResult ({
                  \$dummy [106],\$dummy [107],\$dummy [108],\$dummy [109],
                  \$dummy [110],\$dummy [111],\$dummy [112],\$dummy [113]}), .BoothAddingOperand (
                  {L1_0_L2_3_G1_MINI_ALU_BoothOperand_16,
                  L1_0_L2_3_G1_MINI_ALU_BoothOperand_15,
                  L1_0_L2_3_G1_MINI_ALU_BoothOperand_14,
                  L1_0_L2_3_G1_MINI_ALU_BoothOperand_13,
                  L1_0_L2_3_G1_MINI_ALU_BoothOperand_12,
                  L1_0_L2_3_G1_MINI_ALU_BoothOperand_11,
                  L1_0_L2_3_G1_MINI_ALU_BoothOperand_10,
                  L1_0_L2_3_G1_MINI_ALU_BoothOperand_9,\$dummy [114],
                  \$dummy [115],\$dummy [116],\$dummy [117],\$dummy [118],
                  \$dummy [119],\$dummy [120],\$dummy [121],\$dummy [122]}), .BoothP (
                  {L1_0_L2_3_G1_MINI_ALU_BoothP_16,
                  L1_0_L2_3_G1_MINI_ALU_BoothP_15,
                  L1_0_L2_3_G1_MINI_ALU_BoothP_14,
                  L1_0_L2_3_G1_MINI_ALU_BoothP_13,
                  L1_0_L2_3_G1_MINI_ALU_BoothP_12,
                  L1_0_L2_3_G1_MINI_ALU_BoothP_11,
                  L1_0_L2_3_G1_MINI_ALU_BoothP_10,L1_0_L2_3_G1_MINI_ALU_BoothP_9
                  ,L1_0_L2_3_G1_MINI_ALU_BoothP_8,L1_0_L2_3_G1_MINI_ALU_BoothP_7
                  ,L1_0_L2_3_G1_MINI_ALU_BoothP_6,L1_0_L2_3_G1_MINI_ALU_BoothP_5
                  ,L1_0_L2_3_G1_MINI_ALU_BoothP_4,L1_0_L2_3_G1_MINI_ALU_BoothP_3
                  ,L1_0_L2_3_G1_MINI_ALU_BoothP_2,L1_0_L2_3_G1_MINI_ALU_BoothP_1
                  ,L1_0_L2_3_G1_MINI_ALU_BoothP_0}), .LargeWindowShifted ({
                  \$dummy [123],\$dummy [124],\$dummy [125],\$dummy [126],
                  \$dummy [127],\$dummy [128],\$dummy [129],\$dummy [130],
                  \$dummy [131],\$dummy [132],\$dummy [133],\$dummy [134],
                  \$dummy [135],\$dummy [136],\$dummy [137],\$dummy [138],
                  \$dummy [139]})) ;
    booth_adder_17 L1_0_L2_4_G1_MINI_ALU_BOOTH_ADDER (.AdderFirstOperand ({
                   L1FirstOperands_12__16,L1FirstOperands_4__15,
                   L1FirstOperands_4__14,L1FirstOperands_4__13,
                   L1FirstOperands_4__12,L1FirstOperands_4__11,
                   L1FirstOperands_4__10,L1FirstOperands_4__9,
                   L1FirstOperands_4__8,L1FirstOperands_4__7,
                   L1FirstOperands_4__6,L1FirstOperands_4__5,
                   L1FirstOperands_4__4,L1FirstOperands_4__3,
                   L1FirstOperands_4__2,L1FirstOperands_4__1,
                   L1FirstOperands_4__0}), .AdderSecondOperand ({
                   L1FirstOperands_12__16,
                   L1_0_L2_4_G1_MINI_ALU_OperationResult_15,
                   L1_0_L2_4_G1_MINI_ALU_OperationResult_14,
                   L1_0_L2_4_G1_MINI_ALU_OperationResult_13,
                   L1_0_L2_4_G1_MINI_ALU_OperationResult_12,
                   L1_0_L2_4_G1_MINI_ALU_OperationResult_11,
                   L1_0_L2_4_G1_MINI_ALU_OperationResult_10,
                   L1_0_L2_4_G1_MINI_ALU_OperationResult_9,
                   L1_0_L2_4_G1_MINI_ALU_OperationResult_8,
                   L1_0_L2_4_G1_MINI_ALU_OperationResult_7,
                   L1_0_L2_4_G1_MINI_ALU_OperationResult_6,
                   L1_0_L2_4_G1_MINI_ALU_OperationResult_5,
                   L1_0_L2_4_G1_MINI_ALU_OperationResult_4,
                   L1_0_L2_4_G1_MINI_ALU_OperationResult_3,
                   L1_0_L2_4_G1_MINI_ALU_OperationResult_2,
                   L1_0_L2_4_G1_MINI_ALU_OperationResult_1,
                   L1_0_L2_4_G1_MINI_ALU_OperationResult_0}), .BoothOperand ({
                   L1_0_L2_4_G1_MINI_ALU_BoothOperand_16,
                   L1_0_L2_4_G1_MINI_ALU_BoothOperand_15,
                   L1_0_L2_4_G1_MINI_ALU_BoothOperand_14,
                   L1_0_L2_4_G1_MINI_ALU_BoothOperand_13,
                   L1_0_L2_4_G1_MINI_ALU_BoothOperand_12,
                   L1_0_L2_4_G1_MINI_ALU_BoothOperand_11,
                   L1_0_L2_4_G1_MINI_ALU_BoothOperand_10,
                   L1_0_L2_4_G1_MINI_ALU_BoothOperand_9,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16}), .BoothP ({
                   L1_0_L2_4_G1_MINI_ALU_BoothP_16,
                   L1_0_L2_4_G1_MINI_ALU_BoothP_15,
                   L1_0_L2_4_G1_MINI_ALU_BoothP_14,
                   L1_0_L2_4_G1_MINI_ALU_BoothP_13,
                   L1_0_L2_4_G1_MINI_ALU_BoothP_12,
                   L1_0_L2_4_G1_MINI_ALU_BoothP_11,
                   L1_0_L2_4_G1_MINI_ALU_BoothP_10,
                   L1_0_L2_4_G1_MINI_ALU_BoothP_9,L1_0_L2_4_G1_MINI_ALU_BoothP_8
                   ,L1_0_L2_4_G1_MINI_ALU_BoothP_7,
                   L1_0_L2_4_G1_MINI_ALU_BoothP_6,L1_0_L2_4_G1_MINI_ALU_BoothP_5
                   ,L1_0_L2_4_G1_MINI_ALU_BoothP_4,
                   L1_0_L2_4_G1_MINI_ALU_BoothP_3,L1_0_L2_4_G1_MINI_ALU_BoothP_2
                   ,L1_0_L2_4_G1_MINI_ALU_BoothP_1,
                   L1_0_L2_4_G1_MINI_ALU_BoothP_0}), .SelOperand (nx3280), .Operation (
                   L1_0_L2_4_G1_MINI_ALU_BoothXORCheck), .AdderResult ({
                   L1ResultsLarge_4__16,L1ResultsLarge_4__15,
                   L1ResultsLarge_4__14,L1ResultsLarge_4__13,
                   L1ResultsLarge_4__12,L1ResultsLarge_4__11,
                   L1ResultsLarge_4__10,L1ResultsLarge_4__9,L1ResultsLarge_4__8,
                   L1ResultsLarge_4__7,L1ResultsLarge_4__6,L1ResultsLarge_4__5,
                   L1ResultsLarge_4__4,L1ResultsLarge_4__3,L1ResultsLarge_4__2,
                   L1ResultsLarge_4__1,L1ResultsLarge_4__0}), .AdderBoothResult (
                   {\$dummy [140],L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_15,
                   L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_14,
                   L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_13,
                   L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_12,
                   L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_11,
                   L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_10,
                   L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_9,
                   L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_8,
                   L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_7,
                   L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_6,
                   L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_5,
                   L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_4,
                   L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_3,
                   L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_2,
                   L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_1,
                   L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_0})) ;
    booth_unit_17 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT (.CLK (CLK), .RST (RST), .Start (
                  Start), .Instr (Instr), .LoopingAndResultNotReady (nx3272), .Filter (
                  {FilterDin_0__4__7,FilterDin_0__4__6,FilterDin_0__4__5,
                  FilterDin_0__4__4,FilterDin_0__4__3,FilterDin_0__4__2,
                  FilterDin_0__4__1,FilterDin_0__4__0}), .Window ({
                  WindowDin_0__4__7,WindowDin_0__4__6,WindowDin_0__4__5,
                  WindowDin_0__4__4,WindowDin_0__4__3,WindowDin_0__4__2,
                  WindowDin_0__4__1,WindowDin_0__4__0}), .AdderBoothResult ({
                  L1FirstOperands_12__16,
                  L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_15,
                  L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_14,
                  L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_13,
                  L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_12,
                  L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_11,
                  L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_10,
                  L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_9,
                  L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_8,
                  L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_7,
                  L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_6,
                  L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_5,
                  L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_4,
                  L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_3,
                  L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_2,
                  L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_1,
                  L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_0}), .BoothXORCheck (
                  L1_0_L2_4_G1_MINI_ALU_BoothXORCheck), .BoothResult ({
                  \$dummy [141],\$dummy [142],\$dummy [143],\$dummy [144],
                  \$dummy [145],\$dummy [146],\$dummy [147],\$dummy [148]}), .BoothAddingOperand (
                  {L1_0_L2_4_G1_MINI_ALU_BoothOperand_16,
                  L1_0_L2_4_G1_MINI_ALU_BoothOperand_15,
                  L1_0_L2_4_G1_MINI_ALU_BoothOperand_14,
                  L1_0_L2_4_G1_MINI_ALU_BoothOperand_13,
                  L1_0_L2_4_G1_MINI_ALU_BoothOperand_12,
                  L1_0_L2_4_G1_MINI_ALU_BoothOperand_11,
                  L1_0_L2_4_G1_MINI_ALU_BoothOperand_10,
                  L1_0_L2_4_G1_MINI_ALU_BoothOperand_9,\$dummy [149],
                  \$dummy [150],\$dummy [151],\$dummy [152],\$dummy [153],
                  \$dummy [154],\$dummy [155],\$dummy [156],\$dummy [157]}), .BoothP (
                  {L1_0_L2_4_G1_MINI_ALU_BoothP_16,
                  L1_0_L2_4_G1_MINI_ALU_BoothP_15,
                  L1_0_L2_4_G1_MINI_ALU_BoothP_14,
                  L1_0_L2_4_G1_MINI_ALU_BoothP_13,
                  L1_0_L2_4_G1_MINI_ALU_BoothP_12,
                  L1_0_L2_4_G1_MINI_ALU_BoothP_11,
                  L1_0_L2_4_G1_MINI_ALU_BoothP_10,L1_0_L2_4_G1_MINI_ALU_BoothP_9
                  ,L1_0_L2_4_G1_MINI_ALU_BoothP_8,L1_0_L2_4_G1_MINI_ALU_BoothP_7
                  ,L1_0_L2_4_G1_MINI_ALU_BoothP_6,L1_0_L2_4_G1_MINI_ALU_BoothP_5
                  ,L1_0_L2_4_G1_MINI_ALU_BoothP_4,L1_0_L2_4_G1_MINI_ALU_BoothP_3
                  ,L1_0_L2_4_G1_MINI_ALU_BoothP_2,L1_0_L2_4_G1_MINI_ALU_BoothP_1
                  ,L1_0_L2_4_G1_MINI_ALU_BoothP_0}), .LargeWindowShifted ({
                  \$dummy [158],\$dummy [159],\$dummy [160],\$dummy [161],
                  \$dummy [162],\$dummy [163],\$dummy [164],\$dummy [165],
                  \$dummy [166],\$dummy [167],\$dummy [168],\$dummy [169],
                  \$dummy [170],\$dummy [171],\$dummy [172],\$dummy [173],
                  \$dummy [174]})) ;
    booth_adder_17 L1_1_L2_0_G1_MINI_ALU_BOOTH_ADDER (.AdderFirstOperand ({
                   L1FirstOperands_12__16,L1FirstOperands_2__15,
                   L1FirstOperands_2__14,L1FirstOperands_2__13,
                   L1FirstOperands_2__12,L1FirstOperands_2__11,
                   L1FirstOperands_2__10,L1FirstOperands_2__9,
                   L1FirstOperands_2__8,L1FirstOperands_2__7,
                   L1FirstOperands_2__6,L1FirstOperands_2__5,
                   L1FirstOperands_2__4,L1FirstOperands_2__3,
                   L1FirstOperands_2__2,L1FirstOperands_2__1,
                   L1FirstOperands_2__0}), .AdderSecondOperand ({
                   L1FirstOperands_12__16,
                   L1_1_L2_0_G1_MINI_ALU_OperationResult_15,
                   L1_1_L2_0_G1_MINI_ALU_OperationResult_14,
                   L1_1_L2_0_G1_MINI_ALU_OperationResult_13,
                   L1_1_L2_0_G1_MINI_ALU_OperationResult_12,
                   L1_1_L2_0_G1_MINI_ALU_OperationResult_11,
                   L1_1_L2_0_G1_MINI_ALU_OperationResult_10,
                   L1_1_L2_0_G1_MINI_ALU_OperationResult_9,
                   L1_1_L2_0_G1_MINI_ALU_OperationResult_8,
                   L1_1_L2_0_G1_MINI_ALU_OperationResult_7,
                   L1_1_L2_0_G1_MINI_ALU_OperationResult_6,
                   L1_1_L2_0_G1_MINI_ALU_OperationResult_5,
                   L1_1_L2_0_G1_MINI_ALU_OperationResult_4,
                   L1_1_L2_0_G1_MINI_ALU_OperationResult_3,
                   L1_1_L2_0_G1_MINI_ALU_OperationResult_2,
                   L1_1_L2_0_G1_MINI_ALU_OperationResult_1,
                   L1_1_L2_0_G1_MINI_ALU_OperationResult_0}), .BoothOperand ({
                   L1_1_L2_0_G1_MINI_ALU_BoothOperand_16,
                   L1_1_L2_0_G1_MINI_ALU_BoothOperand_15,
                   L1_1_L2_0_G1_MINI_ALU_BoothOperand_14,
                   L1_1_L2_0_G1_MINI_ALU_BoothOperand_13,
                   L1_1_L2_0_G1_MINI_ALU_BoothOperand_12,
                   L1_1_L2_0_G1_MINI_ALU_BoothOperand_11,
                   L1_1_L2_0_G1_MINI_ALU_BoothOperand_10,
                   L1_1_L2_0_G1_MINI_ALU_BoothOperand_9,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16}), .BoothP ({
                   L1_1_L2_0_G1_MINI_ALU_BoothP_16,
                   L1_1_L2_0_G1_MINI_ALU_BoothP_15,
                   L1_1_L2_0_G1_MINI_ALU_BoothP_14,
                   L1_1_L2_0_G1_MINI_ALU_BoothP_13,
                   L1_1_L2_0_G1_MINI_ALU_BoothP_12,
                   L1_1_L2_0_G1_MINI_ALU_BoothP_11,
                   L1_1_L2_0_G1_MINI_ALU_BoothP_10,
                   L1_1_L2_0_G1_MINI_ALU_BoothP_9,L1_1_L2_0_G1_MINI_ALU_BoothP_8
                   ,L1_1_L2_0_G1_MINI_ALU_BoothP_7,
                   L1_1_L2_0_G1_MINI_ALU_BoothP_6,L1_1_L2_0_G1_MINI_ALU_BoothP_5
                   ,L1_1_L2_0_G1_MINI_ALU_BoothP_4,
                   L1_1_L2_0_G1_MINI_ALU_BoothP_3,L1_1_L2_0_G1_MINI_ALU_BoothP_2
                   ,L1_1_L2_0_G1_MINI_ALU_BoothP_1,
                   L1_1_L2_0_G1_MINI_ALU_BoothP_0}), .SelOperand (nx3280), .Operation (
                   L1_1_L2_0_G1_MINI_ALU_BoothXORCheck), .AdderResult ({
                   L1ResultsLarge_5__16,L1ResultsLarge_5__15,
                   L1ResultsLarge_5__14,L1ResultsLarge_5__13,
                   L1ResultsLarge_5__12,L1ResultsLarge_5__11,
                   L1ResultsLarge_5__10,L1ResultsLarge_5__9,L1ResultsLarge_5__8,
                   L1ResultsLarge_5__7,L1ResultsLarge_5__6,L1ResultsLarge_5__5,
                   L1ResultsLarge_5__4,L1ResultsLarge_5__3,L1ResultsLarge_5__2,
                   L1ResultsLarge_5__1,L1ResultsLarge_5__0}), .AdderBoothResult (
                   {\$dummy [175],L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_15,
                   L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_14,
                   L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_13,
                   L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_12,
                   L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_11,
                   L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_10,
                   L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_9,
                   L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_8,
                   L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_7,
                   L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_6,
                   L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_5,
                   L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_4,
                   L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_3,
                   L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_2,
                   L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_1,
                   L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_0})) ;
    booth_unit_17 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT (.CLK (CLK), .RST (RST), .Start (
                  Start), .Instr (Instr), .LoopingAndResultNotReady (nx3272), .Filter (
                  {FilterDin_1__0__7,FilterDin_1__0__6,FilterDin_1__0__5,
                  FilterDin_1__0__4,FilterDin_1__0__3,FilterDin_1__0__2,
                  FilterDin_1__0__1,FilterDin_1__0__0}), .Window ({
                  WindowDin_1__0__7,WindowDin_1__0__6,WindowDin_1__0__5,
                  WindowDin_1__0__4,WindowDin_1__0__3,WindowDin_1__0__2,
                  WindowDin_1__0__1,WindowDin_1__0__0}), .AdderBoothResult ({
                  L1FirstOperands_12__16,
                  L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_15,
                  L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_14,
                  L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_13,
                  L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_12,
                  L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_11,
                  L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_10,
                  L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_9,
                  L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_8,
                  L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_7,
                  L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_6,
                  L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_5,
                  L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_4,
                  L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_3,
                  L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_2,
                  L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_1,
                  L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_0}), .BoothXORCheck (
                  L1_1_L2_0_G1_MINI_ALU_BoothXORCheck), .BoothResult ({
                  \$dummy [176],\$dummy [177],\$dummy [178],\$dummy [179],
                  \$dummy [180],\$dummy [181],\$dummy [182],\$dummy [183]}), .BoothAddingOperand (
                  {L1_1_L2_0_G1_MINI_ALU_BoothOperand_16,
                  L1_1_L2_0_G1_MINI_ALU_BoothOperand_15,
                  L1_1_L2_0_G1_MINI_ALU_BoothOperand_14,
                  L1_1_L2_0_G1_MINI_ALU_BoothOperand_13,
                  L1_1_L2_0_G1_MINI_ALU_BoothOperand_12,
                  L1_1_L2_0_G1_MINI_ALU_BoothOperand_11,
                  L1_1_L2_0_G1_MINI_ALU_BoothOperand_10,
                  L1_1_L2_0_G1_MINI_ALU_BoothOperand_9,\$dummy [184],
                  \$dummy [185],\$dummy [186],\$dummy [187],\$dummy [188],
                  \$dummy [189],\$dummy [190],\$dummy [191],\$dummy [192]}), .BoothP (
                  {L1_1_L2_0_G1_MINI_ALU_BoothP_16,
                  L1_1_L2_0_G1_MINI_ALU_BoothP_15,
                  L1_1_L2_0_G1_MINI_ALU_BoothP_14,
                  L1_1_L2_0_G1_MINI_ALU_BoothP_13,
                  L1_1_L2_0_G1_MINI_ALU_BoothP_12,
                  L1_1_L2_0_G1_MINI_ALU_BoothP_11,
                  L1_1_L2_0_G1_MINI_ALU_BoothP_10,L1_1_L2_0_G1_MINI_ALU_BoothP_9
                  ,L1_1_L2_0_G1_MINI_ALU_BoothP_8,L1_1_L2_0_G1_MINI_ALU_BoothP_7
                  ,L1_1_L2_0_G1_MINI_ALU_BoothP_6,L1_1_L2_0_G1_MINI_ALU_BoothP_5
                  ,L1_1_L2_0_G1_MINI_ALU_BoothP_4,L1_1_L2_0_G1_MINI_ALU_BoothP_3
                  ,L1_1_L2_0_G1_MINI_ALU_BoothP_2,L1_1_L2_0_G1_MINI_ALU_BoothP_1
                  ,L1_1_L2_0_G1_MINI_ALU_BoothP_0}), .LargeWindowShifted ({
                  \$dummy [193],\$dummy [194],\$dummy [195],\$dummy [196],
                  \$dummy [197],\$dummy [198],\$dummy [199],\$dummy [200],
                  \$dummy [201],\$dummy [202],\$dummy [203],\$dummy [204],
                  \$dummy [205],\$dummy [206],\$dummy [207],\$dummy [208],
                  \$dummy [209]})) ;
    booth_adder_17 L1_1_L2_1_G1_MINI_ALU_BOOTH_ADDER (.AdderFirstOperand ({
                   L1FirstOperands_12__16,L1FirstOperands_6__15,
                   L1FirstOperands_6__14,L1FirstOperands_6__13,
                   L1FirstOperands_6__12,L1FirstOperands_6__11,
                   L1FirstOperands_6__10,L1FirstOperands_6__9,
                   L1FirstOperands_6__8,L1FirstOperands_6__7,
                   L1FirstOperands_6__6,L1FirstOperands_6__5,
                   L1FirstOperands_6__4,L1FirstOperands_6__3,
                   L1FirstOperands_6__2,L1FirstOperands_6__1,
                   L1FirstOperands_6__0}), .AdderSecondOperand ({
                   L1FirstOperands_12__16,
                   L1_1_L2_1_G1_MINI_ALU_OperationResult_15,
                   L1_1_L2_1_G1_MINI_ALU_OperationResult_14,
                   L1_1_L2_1_G1_MINI_ALU_OperationResult_13,
                   L1_1_L2_1_G1_MINI_ALU_OperationResult_12,
                   L1_1_L2_1_G1_MINI_ALU_OperationResult_11,
                   L1_1_L2_1_G1_MINI_ALU_OperationResult_10,
                   L1_1_L2_1_G1_MINI_ALU_OperationResult_9,
                   L1_1_L2_1_G1_MINI_ALU_OperationResult_8,
                   L1_1_L2_1_G1_MINI_ALU_OperationResult_7,
                   L1_1_L2_1_G1_MINI_ALU_OperationResult_6,
                   L1_1_L2_1_G1_MINI_ALU_OperationResult_5,
                   L1_1_L2_1_G1_MINI_ALU_OperationResult_4,
                   L1_1_L2_1_G1_MINI_ALU_OperationResult_3,
                   L1_1_L2_1_G1_MINI_ALU_OperationResult_2,
                   L1_1_L2_1_G1_MINI_ALU_OperationResult_1,
                   L1_1_L2_1_G1_MINI_ALU_OperationResult_0}), .BoothOperand ({
                   L1_1_L2_1_G1_MINI_ALU_BoothOperand_16,
                   L1_1_L2_1_G1_MINI_ALU_BoothOperand_15,
                   L1_1_L2_1_G1_MINI_ALU_BoothOperand_14,
                   L1_1_L2_1_G1_MINI_ALU_BoothOperand_13,
                   L1_1_L2_1_G1_MINI_ALU_BoothOperand_12,
                   L1_1_L2_1_G1_MINI_ALU_BoothOperand_11,
                   L1_1_L2_1_G1_MINI_ALU_BoothOperand_10,
                   L1_1_L2_1_G1_MINI_ALU_BoothOperand_9,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16}), .BoothP ({
                   L1_1_L2_1_G1_MINI_ALU_BoothP_16,
                   L1_1_L2_1_G1_MINI_ALU_BoothP_15,
                   L1_1_L2_1_G1_MINI_ALU_BoothP_14,
                   L1_1_L2_1_G1_MINI_ALU_BoothP_13,
                   L1_1_L2_1_G1_MINI_ALU_BoothP_12,
                   L1_1_L2_1_G1_MINI_ALU_BoothP_11,
                   L1_1_L2_1_G1_MINI_ALU_BoothP_10,
                   L1_1_L2_1_G1_MINI_ALU_BoothP_9,L1_1_L2_1_G1_MINI_ALU_BoothP_8
                   ,L1_1_L2_1_G1_MINI_ALU_BoothP_7,
                   L1_1_L2_1_G1_MINI_ALU_BoothP_6,L1_1_L2_1_G1_MINI_ALU_BoothP_5
                   ,L1_1_L2_1_G1_MINI_ALU_BoothP_4,
                   L1_1_L2_1_G1_MINI_ALU_BoothP_3,L1_1_L2_1_G1_MINI_ALU_BoothP_2
                   ,L1_1_L2_1_G1_MINI_ALU_BoothP_1,
                   L1_1_L2_1_G1_MINI_ALU_BoothP_0}), .SelOperand (nx3280), .Operation (
                   L1_1_L2_1_G1_MINI_ALU_BoothXORCheck), .AdderResult ({
                   L1ResultsLarge_6__16,L1ResultsLarge_6__15,
                   L1ResultsLarge_6__14,L1ResultsLarge_6__13,
                   L1ResultsLarge_6__12,L1ResultsLarge_6__11,
                   L1ResultsLarge_6__10,L1ResultsLarge_6__9,L1ResultsLarge_6__8,
                   L1ResultsLarge_6__7,L1ResultsLarge_6__6,L1ResultsLarge_6__5,
                   L1ResultsLarge_6__4,L1ResultsLarge_6__3,L1ResultsLarge_6__2,
                   L1ResultsLarge_6__1,L1ResultsLarge_6__0}), .AdderBoothResult (
                   {\$dummy [210],L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_15,
                   L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_14,
                   L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_13,
                   L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_12,
                   L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_11,
                   L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_10,
                   L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_9,
                   L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_8,
                   L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_7,
                   L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_6,
                   L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_5,
                   L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_4,
                   L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_3,
                   L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_2,
                   L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_1,
                   L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_0})) ;
    booth_unit_17 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT (.CLK (CLK), .RST (RST), .Start (
                  Start), .Instr (Instr), .LoopingAndResultNotReady (nx3272), .Filter (
                  {FilterDin_1__1__7,FilterDin_1__1__6,FilterDin_1__1__5,
                  FilterDin_1__1__4,FilterDin_1__1__3,FilterDin_1__1__2,
                  FilterDin_1__1__1,FilterDin_1__1__0}), .Window ({
                  WindowDin_1__1__7,WindowDin_1__1__6,WindowDin_1__1__5,
                  WindowDin_1__1__4,WindowDin_1__1__3,WindowDin_1__1__2,
                  WindowDin_1__1__1,WindowDin_1__1__0}), .AdderBoothResult ({
                  L1FirstOperands_12__16,
                  L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_15,
                  L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_14,
                  L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_13,
                  L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_12,
                  L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_11,
                  L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_10,
                  L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_9,
                  L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_8,
                  L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_7,
                  L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_6,
                  L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_5,
                  L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_4,
                  L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_3,
                  L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_2,
                  L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_1,
                  L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_0}), .BoothXORCheck (
                  L1_1_L2_1_G1_MINI_ALU_BoothXORCheck), .BoothResult ({
                  \$dummy [211],\$dummy [212],\$dummy [213],\$dummy [214],
                  \$dummy [215],\$dummy [216],\$dummy [217],\$dummy [218]}), .BoothAddingOperand (
                  {L1_1_L2_1_G1_MINI_ALU_BoothOperand_16,
                  L1_1_L2_1_G1_MINI_ALU_BoothOperand_15,
                  L1_1_L2_1_G1_MINI_ALU_BoothOperand_14,
                  L1_1_L2_1_G1_MINI_ALU_BoothOperand_13,
                  L1_1_L2_1_G1_MINI_ALU_BoothOperand_12,
                  L1_1_L2_1_G1_MINI_ALU_BoothOperand_11,
                  L1_1_L2_1_G1_MINI_ALU_BoothOperand_10,
                  L1_1_L2_1_G1_MINI_ALU_BoothOperand_9,\$dummy [219],
                  \$dummy [220],\$dummy [221],\$dummy [222],\$dummy [223],
                  \$dummy [224],\$dummy [225],\$dummy [226],\$dummy [227]}), .BoothP (
                  {L1_1_L2_1_G1_MINI_ALU_BoothP_16,
                  L1_1_L2_1_G1_MINI_ALU_BoothP_15,
                  L1_1_L2_1_G1_MINI_ALU_BoothP_14,
                  L1_1_L2_1_G1_MINI_ALU_BoothP_13,
                  L1_1_L2_1_G1_MINI_ALU_BoothP_12,
                  L1_1_L2_1_G1_MINI_ALU_BoothP_11,
                  L1_1_L2_1_G1_MINI_ALU_BoothP_10,L1_1_L2_1_G1_MINI_ALU_BoothP_9
                  ,L1_1_L2_1_G1_MINI_ALU_BoothP_8,L1_1_L2_1_G1_MINI_ALU_BoothP_7
                  ,L1_1_L2_1_G1_MINI_ALU_BoothP_6,L1_1_L2_1_G1_MINI_ALU_BoothP_5
                  ,L1_1_L2_1_G1_MINI_ALU_BoothP_4,L1_1_L2_1_G1_MINI_ALU_BoothP_3
                  ,L1_1_L2_1_G1_MINI_ALU_BoothP_2,L1_1_L2_1_G1_MINI_ALU_BoothP_1
                  ,L1_1_L2_1_G1_MINI_ALU_BoothP_0}), .LargeWindowShifted ({
                  \$dummy [228],\$dummy [229],\$dummy [230],\$dummy [231],
                  \$dummy [232],\$dummy [233],\$dummy [234],\$dummy [235],
                  \$dummy [236],\$dummy [237],\$dummy [238],\$dummy [239],
                  \$dummy [240],\$dummy [241],\$dummy [242],\$dummy [243],
                  \$dummy [244]})) ;
    booth_adder_17 L1_1_L2_2_G1_MINI_ALU_BOOTH_ADDER (.AdderFirstOperand ({
                   L1FirstOperands_12__16,L1FirstOperands_7__15,
                   L1FirstOperands_7__14,L1FirstOperands_7__13,
                   L1FirstOperands_7__12,L1FirstOperands_7__11,
                   L1FirstOperands_7__10,L1FirstOperands_7__9,
                   L1FirstOperands_7__8,L1FirstOperands_7__7,
                   L1FirstOperands_7__6,L1FirstOperands_7__5,
                   L1FirstOperands_7__4,L1FirstOperands_7__3,
                   L1FirstOperands_7__2,L1FirstOperands_7__1,
                   L1FirstOperands_7__0}), .AdderSecondOperand ({
                   L1FirstOperands_12__16,
                   L1_1_L2_2_G1_MINI_ALU_OperationResult_15,
                   L1_1_L2_2_G1_MINI_ALU_OperationResult_14,
                   L1_1_L2_2_G1_MINI_ALU_OperationResult_13,
                   L1_1_L2_2_G1_MINI_ALU_OperationResult_12,
                   L1_1_L2_2_G1_MINI_ALU_OperationResult_11,
                   L1_1_L2_2_G1_MINI_ALU_OperationResult_10,
                   L1_1_L2_2_G1_MINI_ALU_OperationResult_9,
                   L1_1_L2_2_G1_MINI_ALU_OperationResult_8,
                   L1_1_L2_2_G1_MINI_ALU_OperationResult_7,
                   L1_1_L2_2_G1_MINI_ALU_OperationResult_6,
                   L1_1_L2_2_G1_MINI_ALU_OperationResult_5,
                   L1_1_L2_2_G1_MINI_ALU_OperationResult_4,
                   L1_1_L2_2_G1_MINI_ALU_OperationResult_3,
                   L1_1_L2_2_G1_MINI_ALU_OperationResult_2,
                   L1_1_L2_2_G1_MINI_ALU_OperationResult_1,
                   L1_1_L2_2_G1_MINI_ALU_OperationResult_0}), .BoothOperand ({
                   L1_1_L2_2_G1_MINI_ALU_BoothOperand_16,
                   L1_1_L2_2_G1_MINI_ALU_BoothOperand_15,
                   L1_1_L2_2_G1_MINI_ALU_BoothOperand_14,
                   L1_1_L2_2_G1_MINI_ALU_BoothOperand_13,
                   L1_1_L2_2_G1_MINI_ALU_BoothOperand_12,
                   L1_1_L2_2_G1_MINI_ALU_BoothOperand_11,
                   L1_1_L2_2_G1_MINI_ALU_BoothOperand_10,
                   L1_1_L2_2_G1_MINI_ALU_BoothOperand_9,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16}), .BoothP ({
                   L1_1_L2_2_G1_MINI_ALU_BoothP_16,
                   L1_1_L2_2_G1_MINI_ALU_BoothP_15,
                   L1_1_L2_2_G1_MINI_ALU_BoothP_14,
                   L1_1_L2_2_G1_MINI_ALU_BoothP_13,
                   L1_1_L2_2_G1_MINI_ALU_BoothP_12,
                   L1_1_L2_2_G1_MINI_ALU_BoothP_11,
                   L1_1_L2_2_G1_MINI_ALU_BoothP_10,
                   L1_1_L2_2_G1_MINI_ALU_BoothP_9,L1_1_L2_2_G1_MINI_ALU_BoothP_8
                   ,L1_1_L2_2_G1_MINI_ALU_BoothP_7,
                   L1_1_L2_2_G1_MINI_ALU_BoothP_6,L1_1_L2_2_G1_MINI_ALU_BoothP_5
                   ,L1_1_L2_2_G1_MINI_ALU_BoothP_4,
                   L1_1_L2_2_G1_MINI_ALU_BoothP_3,L1_1_L2_2_G1_MINI_ALU_BoothP_2
                   ,L1_1_L2_2_G1_MINI_ALU_BoothP_1,
                   L1_1_L2_2_G1_MINI_ALU_BoothP_0}), .SelOperand (nx3280), .Operation (
                   L1_1_L2_2_G1_MINI_ALU_BoothXORCheck), .AdderResult ({
                   L1ResultsLarge_7__16,L1ResultsLarge_7__15,
                   L1ResultsLarge_7__14,L1ResultsLarge_7__13,
                   L1ResultsLarge_7__12,L1ResultsLarge_7__11,
                   L1ResultsLarge_7__10,L1ResultsLarge_7__9,L1ResultsLarge_7__8,
                   L1ResultsLarge_7__7,L1ResultsLarge_7__6,L1ResultsLarge_7__5,
                   L1ResultsLarge_7__4,L1ResultsLarge_7__3,L1ResultsLarge_7__2,
                   L1ResultsLarge_7__1,L1ResultsLarge_7__0}), .AdderBoothResult (
                   {\$dummy [245],L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_15,
                   L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_14,
                   L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_13,
                   L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_12,
                   L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_11,
                   L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_10,
                   L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_9,
                   L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_8,
                   L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_7,
                   L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_6,
                   L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_5,
                   L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_4,
                   L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_3,
                   L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_2,
                   L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_1,
                   L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_0})) ;
    booth_unit_17 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT (.CLK (CLK), .RST (RST), .Start (
                  Start), .Instr (Instr), .LoopingAndResultNotReady (nx3274), .Filter (
                  {FilterDin_1__2__7,FilterDin_1__2__6,FilterDin_1__2__5,
                  FilterDin_1__2__4,FilterDin_1__2__3,FilterDin_1__2__2,
                  FilterDin_1__2__1,FilterDin_1__2__0}), .Window ({
                  WindowDin_1__2__7,WindowDin_1__2__6,WindowDin_1__2__5,
                  WindowDin_1__2__4,WindowDin_1__2__3,WindowDin_1__2__2,
                  WindowDin_1__2__1,WindowDin_1__2__0}), .AdderBoothResult ({
                  L1FirstOperands_12__16,
                  L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_15,
                  L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_14,
                  L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_13,
                  L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_12,
                  L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_11,
                  L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_10,
                  L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_9,
                  L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_8,
                  L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_7,
                  L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_6,
                  L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_5,
                  L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_4,
                  L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_3,
                  L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_2,
                  L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_1,
                  L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_0}), .BoothXORCheck (
                  L1_1_L2_2_G1_MINI_ALU_BoothXORCheck), .BoothResult ({
                  \$dummy [246],\$dummy [247],\$dummy [248],\$dummy [249],
                  \$dummy [250],\$dummy [251],\$dummy [252],\$dummy [253]}), .BoothAddingOperand (
                  {L1_1_L2_2_G1_MINI_ALU_BoothOperand_16,
                  L1_1_L2_2_G1_MINI_ALU_BoothOperand_15,
                  L1_1_L2_2_G1_MINI_ALU_BoothOperand_14,
                  L1_1_L2_2_G1_MINI_ALU_BoothOperand_13,
                  L1_1_L2_2_G1_MINI_ALU_BoothOperand_12,
                  L1_1_L2_2_G1_MINI_ALU_BoothOperand_11,
                  L1_1_L2_2_G1_MINI_ALU_BoothOperand_10,
                  L1_1_L2_2_G1_MINI_ALU_BoothOperand_9,\$dummy [254],
                  \$dummy [255],\$dummy [256],\$dummy [257],\$dummy [258],
                  \$dummy [259],\$dummy [260],\$dummy [261],\$dummy [262]}), .BoothP (
                  {L1_1_L2_2_G1_MINI_ALU_BoothP_16,
                  L1_1_L2_2_G1_MINI_ALU_BoothP_15,
                  L1_1_L2_2_G1_MINI_ALU_BoothP_14,
                  L1_1_L2_2_G1_MINI_ALU_BoothP_13,
                  L1_1_L2_2_G1_MINI_ALU_BoothP_12,
                  L1_1_L2_2_G1_MINI_ALU_BoothP_11,
                  L1_1_L2_2_G1_MINI_ALU_BoothP_10,L1_1_L2_2_G1_MINI_ALU_BoothP_9
                  ,L1_1_L2_2_G1_MINI_ALU_BoothP_8,L1_1_L2_2_G1_MINI_ALU_BoothP_7
                  ,L1_1_L2_2_G1_MINI_ALU_BoothP_6,L1_1_L2_2_G1_MINI_ALU_BoothP_5
                  ,L1_1_L2_2_G1_MINI_ALU_BoothP_4,L1_1_L2_2_G1_MINI_ALU_BoothP_3
                  ,L1_1_L2_2_G1_MINI_ALU_BoothP_2,L1_1_L2_2_G1_MINI_ALU_BoothP_1
                  ,L1_1_L2_2_G1_MINI_ALU_BoothP_0}), .LargeWindowShifted ({
                  \$dummy [263],\$dummy [264],\$dummy [265],\$dummy [266],
                  \$dummy [267],\$dummy [268],\$dummy [269],\$dummy [270],
                  \$dummy [271],\$dummy [272],\$dummy [273],\$dummy [274],
                  \$dummy [275],\$dummy [276],\$dummy [277],\$dummy [278],
                  \$dummy [279]})) ;
    booth_adder_17 L1_1_L2_3_G1_MINI_ALU_BOOTH_ADDER (.AdderFirstOperand ({
                   L1FirstOperands_12__16,L1FirstOperands_8__15,
                   L1FirstOperands_8__14,L1FirstOperands_8__13,
                   L1FirstOperands_8__12,L1FirstOperands_8__11,
                   L1FirstOperands_8__10,L1FirstOperands_8__9,
                   L1FirstOperands_8__8,L1FirstOperands_8__7,
                   L1FirstOperands_8__6,L1FirstOperands_8__5,
                   L1FirstOperands_8__4,L1FirstOperands_8__3,
                   L1FirstOperands_8__2,L1FirstOperands_8__1,
                   L1FirstOperands_8__0}), .AdderSecondOperand ({
                   L1FirstOperands_12__16,
                   L1_1_L2_3_G1_MINI_ALU_OperationResult_15,
                   L1_1_L2_3_G1_MINI_ALU_OperationResult_14,
                   L1_1_L2_3_G1_MINI_ALU_OperationResult_13,
                   L1_1_L2_3_G1_MINI_ALU_OperationResult_12,
                   L1_1_L2_3_G1_MINI_ALU_OperationResult_11,
                   L1_1_L2_3_G1_MINI_ALU_OperationResult_10,
                   L1_1_L2_3_G1_MINI_ALU_OperationResult_9,
                   L1_1_L2_3_G1_MINI_ALU_OperationResult_8,
                   L1_1_L2_3_G1_MINI_ALU_OperationResult_7,
                   L1_1_L2_3_G1_MINI_ALU_OperationResult_6,
                   L1_1_L2_3_G1_MINI_ALU_OperationResult_5,
                   L1_1_L2_3_G1_MINI_ALU_OperationResult_4,
                   L1_1_L2_3_G1_MINI_ALU_OperationResult_3,
                   L1_1_L2_3_G1_MINI_ALU_OperationResult_2,
                   L1_1_L2_3_G1_MINI_ALU_OperationResult_1,
                   L1_1_L2_3_G1_MINI_ALU_OperationResult_0}), .BoothOperand ({
                   L1_1_L2_3_G1_MINI_ALU_BoothOperand_16,
                   L1_1_L2_3_G1_MINI_ALU_BoothOperand_15,
                   L1_1_L2_3_G1_MINI_ALU_BoothOperand_14,
                   L1_1_L2_3_G1_MINI_ALU_BoothOperand_13,
                   L1_1_L2_3_G1_MINI_ALU_BoothOperand_12,
                   L1_1_L2_3_G1_MINI_ALU_BoothOperand_11,
                   L1_1_L2_3_G1_MINI_ALU_BoothOperand_10,
                   L1_1_L2_3_G1_MINI_ALU_BoothOperand_9,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16}), .BoothP ({
                   L1_1_L2_3_G1_MINI_ALU_BoothP_16,
                   L1_1_L2_3_G1_MINI_ALU_BoothP_15,
                   L1_1_L2_3_G1_MINI_ALU_BoothP_14,
                   L1_1_L2_3_G1_MINI_ALU_BoothP_13,
                   L1_1_L2_3_G1_MINI_ALU_BoothP_12,
                   L1_1_L2_3_G1_MINI_ALU_BoothP_11,
                   L1_1_L2_3_G1_MINI_ALU_BoothP_10,
                   L1_1_L2_3_G1_MINI_ALU_BoothP_9,L1_1_L2_3_G1_MINI_ALU_BoothP_8
                   ,L1_1_L2_3_G1_MINI_ALU_BoothP_7,
                   L1_1_L2_3_G1_MINI_ALU_BoothP_6,L1_1_L2_3_G1_MINI_ALU_BoothP_5
                   ,L1_1_L2_3_G1_MINI_ALU_BoothP_4,
                   L1_1_L2_3_G1_MINI_ALU_BoothP_3,L1_1_L2_3_G1_MINI_ALU_BoothP_2
                   ,L1_1_L2_3_G1_MINI_ALU_BoothP_1,
                   L1_1_L2_3_G1_MINI_ALU_BoothP_0}), .SelOperand (nx3282), .Operation (
                   L1_1_L2_3_G1_MINI_ALU_BoothXORCheck), .AdderResult ({
                   L1ResultsLarge_8__16,L1ResultsLarge_8__15,
                   L1ResultsLarge_8__14,L1ResultsLarge_8__13,
                   L1ResultsLarge_8__12,L1ResultsLarge_8__11,
                   L1ResultsLarge_8__10,L1ResultsLarge_8__9,L1ResultsLarge_8__8,
                   L1ResultsLarge_8__7,L1ResultsLarge_8__6,L1ResultsLarge_8__5,
                   L1ResultsLarge_8__4,L1ResultsLarge_8__3,L1ResultsLarge_8__2,
                   L1ResultsLarge_8__1,L1ResultsLarge_8__0}), .AdderBoothResult (
                   {\$dummy [280],L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_15,
                   L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_14,
                   L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_13,
                   L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_12,
                   L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_11,
                   L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_10,
                   L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_9,
                   L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_8,
                   L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_7,
                   L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_6,
                   L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_5,
                   L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_4,
                   L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_3,
                   L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_2,
                   L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_1,
                   L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_0})) ;
    booth_unit_17 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT (.CLK (CLK), .RST (RST), .Start (
                  Start), .Instr (Instr), .LoopingAndResultNotReady (nx3274), .Filter (
                  {FilterDin_1__3__7,FilterDin_1__3__6,FilterDin_1__3__5,
                  FilterDin_1__3__4,FilterDin_1__3__3,FilterDin_1__3__2,
                  FilterDin_1__3__1,FilterDin_1__3__0}), .Window ({
                  WindowDin_1__3__7,WindowDin_1__3__6,WindowDin_1__3__5,
                  WindowDin_1__3__4,WindowDin_1__3__3,WindowDin_1__3__2,
                  WindowDin_1__3__1,WindowDin_1__3__0}), .AdderBoothResult ({
                  L1FirstOperands_12__16,
                  L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_15,
                  L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_14,
                  L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_13,
                  L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_12,
                  L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_11,
                  L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_10,
                  L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_9,
                  L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_8,
                  L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_7,
                  L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_6,
                  L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_5,
                  L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_4,
                  L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_3,
                  L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_2,
                  L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_1,
                  L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_0}), .BoothXORCheck (
                  L1_1_L2_3_G1_MINI_ALU_BoothXORCheck), .BoothResult ({
                  \$dummy [281],\$dummy [282],\$dummy [283],\$dummy [284],
                  \$dummy [285],\$dummy [286],\$dummy [287],\$dummy [288]}), .BoothAddingOperand (
                  {L1_1_L2_3_G1_MINI_ALU_BoothOperand_16,
                  L1_1_L2_3_G1_MINI_ALU_BoothOperand_15,
                  L1_1_L2_3_G1_MINI_ALU_BoothOperand_14,
                  L1_1_L2_3_G1_MINI_ALU_BoothOperand_13,
                  L1_1_L2_3_G1_MINI_ALU_BoothOperand_12,
                  L1_1_L2_3_G1_MINI_ALU_BoothOperand_11,
                  L1_1_L2_3_G1_MINI_ALU_BoothOperand_10,
                  L1_1_L2_3_G1_MINI_ALU_BoothOperand_9,\$dummy [289],
                  \$dummy [290],\$dummy [291],\$dummy [292],\$dummy [293],
                  \$dummy [294],\$dummy [295],\$dummy [296],\$dummy [297]}), .BoothP (
                  {L1_1_L2_3_G1_MINI_ALU_BoothP_16,
                  L1_1_L2_3_G1_MINI_ALU_BoothP_15,
                  L1_1_L2_3_G1_MINI_ALU_BoothP_14,
                  L1_1_L2_3_G1_MINI_ALU_BoothP_13,
                  L1_1_L2_3_G1_MINI_ALU_BoothP_12,
                  L1_1_L2_3_G1_MINI_ALU_BoothP_11,
                  L1_1_L2_3_G1_MINI_ALU_BoothP_10,L1_1_L2_3_G1_MINI_ALU_BoothP_9
                  ,L1_1_L2_3_G1_MINI_ALU_BoothP_8,L1_1_L2_3_G1_MINI_ALU_BoothP_7
                  ,L1_1_L2_3_G1_MINI_ALU_BoothP_6,L1_1_L2_3_G1_MINI_ALU_BoothP_5
                  ,L1_1_L2_3_G1_MINI_ALU_BoothP_4,L1_1_L2_3_G1_MINI_ALU_BoothP_3
                  ,L1_1_L2_3_G1_MINI_ALU_BoothP_2,L1_1_L2_3_G1_MINI_ALU_BoothP_1
                  ,L1_1_L2_3_G1_MINI_ALU_BoothP_0}), .LargeWindowShifted ({
                  \$dummy [298],\$dummy [299],\$dummy [300],\$dummy [301],
                  \$dummy [302],\$dummy [303],\$dummy [304],\$dummy [305],
                  \$dummy [306],\$dummy [307],\$dummy [308],\$dummy [309],
                  \$dummy [310],\$dummy [311],\$dummy [312],\$dummy [313],
                  \$dummy [314]})) ;
    booth_adder_17 L1_1_L2_4_G1_MINI_ALU_BOOTH_ADDER (.AdderFirstOperand ({
                   L1FirstOperands_12__16,L1FirstOperands_4__15,
                   L1FirstOperands_4__14,L1FirstOperands_4__13,
                   L1FirstOperands_4__12,L1FirstOperands_4__11,
                   L1FirstOperands_4__10,L1FirstOperands_4__9,
                   L1FirstOperands_4__8,L1FirstOperands_4__7,
                   L1FirstOperands_4__6,L1FirstOperands_4__5,
                   L1FirstOperands_4__4,L1FirstOperands_4__3,
                   L1FirstOperands_4__2,L1FirstOperands_4__1,
                   L1FirstOperands_4__0}), .AdderSecondOperand ({
                   L1FirstOperands_12__16,
                   L1_1_L2_4_G1_MINI_ALU_OperationResult_15,
                   L1_1_L2_4_G1_MINI_ALU_OperationResult_14,
                   L1_1_L2_4_G1_MINI_ALU_OperationResult_13,
                   L1_1_L2_4_G1_MINI_ALU_OperationResult_12,
                   L1_1_L2_4_G1_MINI_ALU_OperationResult_11,
                   L1_1_L2_4_G1_MINI_ALU_OperationResult_10,
                   L1_1_L2_4_G1_MINI_ALU_OperationResult_9,
                   L1_1_L2_4_G1_MINI_ALU_OperationResult_8,
                   L1_1_L2_4_G1_MINI_ALU_OperationResult_7,
                   L1_1_L2_4_G1_MINI_ALU_OperationResult_6,
                   L1_1_L2_4_G1_MINI_ALU_OperationResult_5,
                   L1_1_L2_4_G1_MINI_ALU_OperationResult_4,
                   L1_1_L2_4_G1_MINI_ALU_OperationResult_3,
                   L1_1_L2_4_G1_MINI_ALU_OperationResult_2,
                   L1_1_L2_4_G1_MINI_ALU_OperationResult_1,
                   L1_1_L2_4_G1_MINI_ALU_OperationResult_0}), .BoothOperand ({
                   L1_1_L2_4_G1_MINI_ALU_BoothOperand_16,
                   L1_1_L2_4_G1_MINI_ALU_BoothOperand_15,
                   L1_1_L2_4_G1_MINI_ALU_BoothOperand_14,
                   L1_1_L2_4_G1_MINI_ALU_BoothOperand_13,
                   L1_1_L2_4_G1_MINI_ALU_BoothOperand_12,
                   L1_1_L2_4_G1_MINI_ALU_BoothOperand_11,
                   L1_1_L2_4_G1_MINI_ALU_BoothOperand_10,
                   L1_1_L2_4_G1_MINI_ALU_BoothOperand_9,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16}), .BoothP ({
                   L1_1_L2_4_G1_MINI_ALU_BoothP_16,
                   L1_1_L2_4_G1_MINI_ALU_BoothP_15,
                   L1_1_L2_4_G1_MINI_ALU_BoothP_14,
                   L1_1_L2_4_G1_MINI_ALU_BoothP_13,
                   L1_1_L2_4_G1_MINI_ALU_BoothP_12,
                   L1_1_L2_4_G1_MINI_ALU_BoothP_11,
                   L1_1_L2_4_G1_MINI_ALU_BoothP_10,
                   L1_1_L2_4_G1_MINI_ALU_BoothP_9,L1_1_L2_4_G1_MINI_ALU_BoothP_8
                   ,L1_1_L2_4_G1_MINI_ALU_BoothP_7,
                   L1_1_L2_4_G1_MINI_ALU_BoothP_6,L1_1_L2_4_G1_MINI_ALU_BoothP_5
                   ,L1_1_L2_4_G1_MINI_ALU_BoothP_4,
                   L1_1_L2_4_G1_MINI_ALU_BoothP_3,L1_1_L2_4_G1_MINI_ALU_BoothP_2
                   ,L1_1_L2_4_G1_MINI_ALU_BoothP_1,
                   L1_1_L2_4_G1_MINI_ALU_BoothP_0}), .SelOperand (nx3282), .Operation (
                   L1_1_L2_4_G1_MINI_ALU_BoothXORCheck), .AdderResult ({
                   L1ResultsLarge_9__16,L1ResultsLarge_9__15,
                   L1ResultsLarge_9__14,L1ResultsLarge_9__13,
                   L1ResultsLarge_9__12,L1ResultsLarge_9__11,
                   L1ResultsLarge_9__10,L1ResultsLarge_9__9,L1ResultsLarge_9__8,
                   L1ResultsLarge_9__7,L1ResultsLarge_9__6,L1ResultsLarge_9__5,
                   L1ResultsLarge_9__4,L1ResultsLarge_9__3,L1ResultsLarge_9__2,
                   L1ResultsLarge_9__1,L1ResultsLarge_9__0}), .AdderBoothResult (
                   {\$dummy [315],L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_15,
                   L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_14,
                   L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_13,
                   L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_12,
                   L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_11,
                   L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_10,
                   L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_9,
                   L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_8,
                   L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_7,
                   L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_6,
                   L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_5,
                   L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_4,
                   L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_3,
                   L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_2,
                   L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_1,
                   L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_0})) ;
    booth_unit_17 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT (.CLK (CLK), .RST (RST), .Start (
                  Start), .Instr (Instr), .LoopingAndResultNotReady (nx3274), .Filter (
                  {FilterDin_1__4__7,FilterDin_1__4__6,FilterDin_1__4__5,
                  FilterDin_1__4__4,FilterDin_1__4__3,FilterDin_1__4__2,
                  FilterDin_1__4__1,FilterDin_1__4__0}), .Window ({
                  WindowDin_1__4__7,WindowDin_1__4__6,WindowDin_1__4__5,
                  WindowDin_1__4__4,WindowDin_1__4__3,WindowDin_1__4__2,
                  WindowDin_1__4__1,WindowDin_1__4__0}), .AdderBoothResult ({
                  L1FirstOperands_12__16,
                  L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_15,
                  L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_14,
                  L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_13,
                  L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_12,
                  L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_11,
                  L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_10,
                  L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_9,
                  L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_8,
                  L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_7,
                  L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_6,
                  L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_5,
                  L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_4,
                  L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_3,
                  L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_2,
                  L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_1,
                  L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_0}), .BoothXORCheck (
                  L1_1_L2_4_G1_MINI_ALU_BoothXORCheck), .BoothResult ({
                  \$dummy [316],\$dummy [317],\$dummy [318],\$dummy [319],
                  \$dummy [320],\$dummy [321],\$dummy [322],\$dummy [323]}), .BoothAddingOperand (
                  {L1_1_L2_4_G1_MINI_ALU_BoothOperand_16,
                  L1_1_L2_4_G1_MINI_ALU_BoothOperand_15,
                  L1_1_L2_4_G1_MINI_ALU_BoothOperand_14,
                  L1_1_L2_4_G1_MINI_ALU_BoothOperand_13,
                  L1_1_L2_4_G1_MINI_ALU_BoothOperand_12,
                  L1_1_L2_4_G1_MINI_ALU_BoothOperand_11,
                  L1_1_L2_4_G1_MINI_ALU_BoothOperand_10,
                  L1_1_L2_4_G1_MINI_ALU_BoothOperand_9,\$dummy [324],
                  \$dummy [325],\$dummy [326],\$dummy [327],\$dummy [328],
                  \$dummy [329],\$dummy [330],\$dummy [331],\$dummy [332]}), .BoothP (
                  {L1_1_L2_4_G1_MINI_ALU_BoothP_16,
                  L1_1_L2_4_G1_MINI_ALU_BoothP_15,
                  L1_1_L2_4_G1_MINI_ALU_BoothP_14,
                  L1_1_L2_4_G1_MINI_ALU_BoothP_13,
                  L1_1_L2_4_G1_MINI_ALU_BoothP_12,
                  L1_1_L2_4_G1_MINI_ALU_BoothP_11,
                  L1_1_L2_4_G1_MINI_ALU_BoothP_10,L1_1_L2_4_G1_MINI_ALU_BoothP_9
                  ,L1_1_L2_4_G1_MINI_ALU_BoothP_8,L1_1_L2_4_G1_MINI_ALU_BoothP_7
                  ,L1_1_L2_4_G1_MINI_ALU_BoothP_6,L1_1_L2_4_G1_MINI_ALU_BoothP_5
                  ,L1_1_L2_4_G1_MINI_ALU_BoothP_4,L1_1_L2_4_G1_MINI_ALU_BoothP_3
                  ,L1_1_L2_4_G1_MINI_ALU_BoothP_2,L1_1_L2_4_G1_MINI_ALU_BoothP_1
                  ,L1_1_L2_4_G1_MINI_ALU_BoothP_0}), .LargeWindowShifted ({
                  \$dummy [333],\$dummy [334],\$dummy [335],\$dummy [336],
                  \$dummy [337],\$dummy [338],\$dummy [339],\$dummy [340],
                  \$dummy [341],\$dummy [342],\$dummy [343],\$dummy [344],
                  \$dummy [345],\$dummy [346],\$dummy [347],\$dummy [348],
                  \$dummy [349]})) ;
    booth_adder_17 L1_2_L2_0_G1_MINI_ALU_BOOTH_ADDER (.AdderFirstOperand ({
                   L1FirstOperands_12__16,L1FirstOperands_10__15,
                   L1FirstOperands_10__14,L1FirstOperands_10__13,
                   L1FirstOperands_10__12,L1FirstOperands_10__11,
                   L1FirstOperands_10__10,L1FirstOperands_10__9,
                   L1FirstOperands_10__8,L1FirstOperands_10__7,
                   L1FirstOperands_10__6,L1FirstOperands_10__5,
                   L1FirstOperands_10__4,L1FirstOperands_10__3,
                   L1FirstOperands_10__2,L1FirstOperands_10__1,
                   L1FirstOperands_10__0}), .AdderSecondOperand ({
                   L1FirstOperands_12__16,
                   L1_2_L2_0_G1_MINI_ALU_OperationResult_15,
                   L1_2_L2_0_G1_MINI_ALU_OperationResult_14,
                   L1_2_L2_0_G1_MINI_ALU_OperationResult_13,
                   L1_2_L2_0_G1_MINI_ALU_OperationResult_12,
                   L1_2_L2_0_G1_MINI_ALU_OperationResult_11,
                   L1_2_L2_0_G1_MINI_ALU_OperationResult_10,
                   L1_2_L2_0_G1_MINI_ALU_OperationResult_9,
                   L1_2_L2_0_G1_MINI_ALU_OperationResult_8,
                   L1_2_L2_0_G1_MINI_ALU_OperationResult_7,
                   L1_2_L2_0_G1_MINI_ALU_OperationResult_6,
                   L1_2_L2_0_G1_MINI_ALU_OperationResult_5,
                   L1_2_L2_0_G1_MINI_ALU_OperationResult_4,
                   L1_2_L2_0_G1_MINI_ALU_OperationResult_3,
                   L1_2_L2_0_G1_MINI_ALU_OperationResult_2,
                   L1_2_L2_0_G1_MINI_ALU_OperationResult_1,
                   L1_2_L2_0_G1_MINI_ALU_OperationResult_0}), .BoothOperand ({
                   L1_2_L2_0_G1_MINI_ALU_BoothOperand_16,
                   L1_2_L2_0_G1_MINI_ALU_BoothOperand_15,
                   L1_2_L2_0_G1_MINI_ALU_BoothOperand_14,
                   L1_2_L2_0_G1_MINI_ALU_BoothOperand_13,
                   L1_2_L2_0_G1_MINI_ALU_BoothOperand_12,
                   L1_2_L2_0_G1_MINI_ALU_BoothOperand_11,
                   L1_2_L2_0_G1_MINI_ALU_BoothOperand_10,
                   L1_2_L2_0_G1_MINI_ALU_BoothOperand_9,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16}), .BoothP ({
                   L1_2_L2_0_G1_MINI_ALU_BoothP_16,
                   L1_2_L2_0_G1_MINI_ALU_BoothP_15,
                   L1_2_L2_0_G1_MINI_ALU_BoothP_14,
                   L1_2_L2_0_G1_MINI_ALU_BoothP_13,
                   L1_2_L2_0_G1_MINI_ALU_BoothP_12,
                   L1_2_L2_0_G1_MINI_ALU_BoothP_11,
                   L1_2_L2_0_G1_MINI_ALU_BoothP_10,
                   L1_2_L2_0_G1_MINI_ALU_BoothP_9,L1_2_L2_0_G1_MINI_ALU_BoothP_8
                   ,L1_2_L2_0_G1_MINI_ALU_BoothP_7,
                   L1_2_L2_0_G1_MINI_ALU_BoothP_6,L1_2_L2_0_G1_MINI_ALU_BoothP_5
                   ,L1_2_L2_0_G1_MINI_ALU_BoothP_4,
                   L1_2_L2_0_G1_MINI_ALU_BoothP_3,L1_2_L2_0_G1_MINI_ALU_BoothP_2
                   ,L1_2_L2_0_G1_MINI_ALU_BoothP_1,
                   L1_2_L2_0_G1_MINI_ALU_BoothP_0}), .SelOperand (nx3282), .Operation (
                   L1_2_L2_0_G1_MINI_ALU_BoothXORCheck), .AdderResult ({
                   L1ResultsLarge_10__16,L1ResultsLarge_10__15,
                   L1ResultsLarge_10__14,L1ResultsLarge_10__13,
                   L1ResultsLarge_10__12,L1ResultsLarge_10__11,
                   L1ResultsLarge_10__10,L1ResultsLarge_10__9,
                   L1ResultsLarge_10__8,L1ResultsLarge_10__7,
                   L1ResultsLarge_10__6,L1ResultsLarge_10__5,
                   L1ResultsLarge_10__4,L1ResultsLarge_10__3,
                   L1ResultsLarge_10__2,L1ResultsLarge_10__1,
                   L1ResultsLarge_10__0}), .AdderBoothResult ({\$dummy [350],
                   L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_15,
                   L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_14,
                   L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_13,
                   L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_12,
                   L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_11,
                   L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_10,
                   L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_9,
                   L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_8,
                   L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_7,
                   L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_6,
                   L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_5,
                   L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_4,
                   L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_3,
                   L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_2,
                   L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_1,
                   L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_0})) ;
    booth_unit_17 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT (.CLK (CLK), .RST (RST), .Start (
                  Start), .Instr (Instr), .LoopingAndResultNotReady (nx3274), .Filter (
                  {FilterDin_2__0__7,FilterDin_2__0__6,FilterDin_2__0__5,
                  FilterDin_2__0__4,FilterDin_2__0__3,FilterDin_2__0__2,
                  FilterDin_2__0__1,FilterDin_2__0__0}), .Window ({
                  WindowDin_2__0__7,WindowDin_2__0__6,WindowDin_2__0__5,
                  WindowDin_2__0__4,WindowDin_2__0__3,WindowDin_2__0__2,
                  WindowDin_2__0__1,WindowDin_2__0__0}), .AdderBoothResult ({
                  L1FirstOperands_12__16,
                  L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_15,
                  L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_14,
                  L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_13,
                  L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_12,
                  L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_11,
                  L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_10,
                  L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_9,
                  L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_8,
                  L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_7,
                  L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_6,
                  L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_5,
                  L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_4,
                  L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_3,
                  L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_2,
                  L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_1,
                  L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_0}), .BoothXORCheck (
                  L1_2_L2_0_G1_MINI_ALU_BoothXORCheck), .BoothResult ({
                  \$dummy [351],\$dummy [352],\$dummy [353],\$dummy [354],
                  \$dummy [355],\$dummy [356],\$dummy [357],\$dummy [358]}), .BoothAddingOperand (
                  {L1_2_L2_0_G1_MINI_ALU_BoothOperand_16,
                  L1_2_L2_0_G1_MINI_ALU_BoothOperand_15,
                  L1_2_L2_0_G1_MINI_ALU_BoothOperand_14,
                  L1_2_L2_0_G1_MINI_ALU_BoothOperand_13,
                  L1_2_L2_0_G1_MINI_ALU_BoothOperand_12,
                  L1_2_L2_0_G1_MINI_ALU_BoothOperand_11,
                  L1_2_L2_0_G1_MINI_ALU_BoothOperand_10,
                  L1_2_L2_0_G1_MINI_ALU_BoothOperand_9,\$dummy [359],
                  \$dummy [360],\$dummy [361],\$dummy [362],\$dummy [363],
                  \$dummy [364],\$dummy [365],\$dummy [366],\$dummy [367]}), .BoothP (
                  {L1_2_L2_0_G1_MINI_ALU_BoothP_16,
                  L1_2_L2_0_G1_MINI_ALU_BoothP_15,
                  L1_2_L2_0_G1_MINI_ALU_BoothP_14,
                  L1_2_L2_0_G1_MINI_ALU_BoothP_13,
                  L1_2_L2_0_G1_MINI_ALU_BoothP_12,
                  L1_2_L2_0_G1_MINI_ALU_BoothP_11,
                  L1_2_L2_0_G1_MINI_ALU_BoothP_10,L1_2_L2_0_G1_MINI_ALU_BoothP_9
                  ,L1_2_L2_0_G1_MINI_ALU_BoothP_8,L1_2_L2_0_G1_MINI_ALU_BoothP_7
                  ,L1_2_L2_0_G1_MINI_ALU_BoothP_6,L1_2_L2_0_G1_MINI_ALU_BoothP_5
                  ,L1_2_L2_0_G1_MINI_ALU_BoothP_4,L1_2_L2_0_G1_MINI_ALU_BoothP_3
                  ,L1_2_L2_0_G1_MINI_ALU_BoothP_2,L1_2_L2_0_G1_MINI_ALU_BoothP_1
                  ,L1_2_L2_0_G1_MINI_ALU_BoothP_0}), .LargeWindowShifted ({
                  \$dummy [368],\$dummy [369],\$dummy [370],\$dummy [371],
                  \$dummy [372],\$dummy [373],\$dummy [374],\$dummy [375],
                  \$dummy [376],\$dummy [377],\$dummy [378],\$dummy [379],
                  \$dummy [380],\$dummy [381],\$dummy [382],\$dummy [383],
                  \$dummy [384]})) ;
    booth_adder_17 L1_2_L2_1_G1_MINI_ALU_BOOTH_ADDER (.AdderFirstOperand ({
                   L1FirstOperands_12__16,L1FirstOperands_11__15,
                   L1FirstOperands_11__14,L1FirstOperands_11__13,
                   L1FirstOperands_11__12,L1FirstOperands_11__11,
                   L1FirstOperands_11__10,L1FirstOperands_11__9,
                   L1FirstOperands_11__8,L1FirstOperands_11__7,
                   L1FirstOperands_11__6,L1FirstOperands_11__5,
                   L1FirstOperands_11__4,L1FirstOperands_11__3,
                   L1FirstOperands_11__2,L1FirstOperands_11__1,
                   L1FirstOperands_11__0}), .AdderSecondOperand ({
                   L1FirstOperands_12__16,
                   L1_2_L2_1_G1_MINI_ALU_OperationResult_15,
                   L1_2_L2_1_G1_MINI_ALU_OperationResult_14,
                   L1_2_L2_1_G1_MINI_ALU_OperationResult_13,
                   L1_2_L2_1_G1_MINI_ALU_OperationResult_12,
                   L1_2_L2_1_G1_MINI_ALU_OperationResult_11,
                   L1_2_L2_1_G1_MINI_ALU_OperationResult_10,
                   L1_2_L2_1_G1_MINI_ALU_OperationResult_9,
                   L1_2_L2_1_G1_MINI_ALU_OperationResult_8,
                   L1_2_L2_1_G1_MINI_ALU_OperationResult_7,
                   L1_2_L2_1_G1_MINI_ALU_OperationResult_6,
                   L1_2_L2_1_G1_MINI_ALU_OperationResult_5,
                   L1_2_L2_1_G1_MINI_ALU_OperationResult_4,
                   L1_2_L2_1_G1_MINI_ALU_OperationResult_3,
                   L1_2_L2_1_G1_MINI_ALU_OperationResult_2,
                   L1_2_L2_1_G1_MINI_ALU_OperationResult_1,
                   L1_2_L2_1_G1_MINI_ALU_OperationResult_0}), .BoothOperand ({
                   L1_2_L2_1_G1_MINI_ALU_BoothOperand_16,
                   L1_2_L2_1_G1_MINI_ALU_BoothOperand_15,
                   L1_2_L2_1_G1_MINI_ALU_BoothOperand_14,
                   L1_2_L2_1_G1_MINI_ALU_BoothOperand_13,
                   L1_2_L2_1_G1_MINI_ALU_BoothOperand_12,
                   L1_2_L2_1_G1_MINI_ALU_BoothOperand_11,
                   L1_2_L2_1_G1_MINI_ALU_BoothOperand_10,
                   L1_2_L2_1_G1_MINI_ALU_BoothOperand_9,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16}), .BoothP ({
                   L1_2_L2_1_G1_MINI_ALU_BoothP_16,
                   L1_2_L2_1_G1_MINI_ALU_BoothP_15,
                   L1_2_L2_1_G1_MINI_ALU_BoothP_14,
                   L1_2_L2_1_G1_MINI_ALU_BoothP_13,
                   L1_2_L2_1_G1_MINI_ALU_BoothP_12,
                   L1_2_L2_1_G1_MINI_ALU_BoothP_11,
                   L1_2_L2_1_G1_MINI_ALU_BoothP_10,
                   L1_2_L2_1_G1_MINI_ALU_BoothP_9,L1_2_L2_1_G1_MINI_ALU_BoothP_8
                   ,L1_2_L2_1_G1_MINI_ALU_BoothP_7,
                   L1_2_L2_1_G1_MINI_ALU_BoothP_6,L1_2_L2_1_G1_MINI_ALU_BoothP_5
                   ,L1_2_L2_1_G1_MINI_ALU_BoothP_4,
                   L1_2_L2_1_G1_MINI_ALU_BoothP_3,L1_2_L2_1_G1_MINI_ALU_BoothP_2
                   ,L1_2_L2_1_G1_MINI_ALU_BoothP_1,
                   L1_2_L2_1_G1_MINI_ALU_BoothP_0}), .SelOperand (nx3282), .Operation (
                   L1_2_L2_1_G1_MINI_ALU_BoothXORCheck), .AdderResult ({
                   L1ResultsLarge_11__16,L1ResultsLarge_11__15,
                   L1ResultsLarge_11__14,L1ResultsLarge_11__13,
                   L1ResultsLarge_11__12,L1ResultsLarge_11__11,
                   L1ResultsLarge_11__10,L1ResultsLarge_11__9,
                   L1ResultsLarge_11__8,L1ResultsLarge_11__7,
                   L1ResultsLarge_11__6,L1ResultsLarge_11__5,
                   L1ResultsLarge_11__4,L1ResultsLarge_11__3,
                   L1ResultsLarge_11__2,L1ResultsLarge_11__1,
                   L1ResultsLarge_11__0}), .AdderBoothResult ({\$dummy [385],
                   L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_15,
                   L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_14,
                   L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_13,
                   L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_12,
                   L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_11,
                   L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_10,
                   L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_9,
                   L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_8,
                   L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_7,
                   L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_6,
                   L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_5,
                   L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_4,
                   L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_3,
                   L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_2,
                   L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_1,
                   L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_0})) ;
    booth_unit_17 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT (.CLK (CLK), .RST (RST), .Start (
                  Start), .Instr (Instr), .LoopingAndResultNotReady (nx3274), .Filter (
                  {FilterDin_2__1__7,FilterDin_2__1__6,FilterDin_2__1__5,
                  FilterDin_2__1__4,FilterDin_2__1__3,FilterDin_2__1__2,
                  FilterDin_2__1__1,FilterDin_2__1__0}), .Window ({
                  WindowDin_2__1__7,WindowDin_2__1__6,WindowDin_2__1__5,
                  WindowDin_2__1__4,WindowDin_2__1__3,WindowDin_2__1__2,
                  WindowDin_2__1__1,WindowDin_2__1__0}), .AdderBoothResult ({
                  L1FirstOperands_12__16,
                  L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_15,
                  L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_14,
                  L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_13,
                  L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_12,
                  L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_11,
                  L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_10,
                  L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_9,
                  L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_8,
                  L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_7,
                  L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_6,
                  L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_5,
                  L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_4,
                  L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_3,
                  L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_2,
                  L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_1,
                  L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_0}), .BoothXORCheck (
                  L1_2_L2_1_G1_MINI_ALU_BoothXORCheck), .BoothResult ({
                  \$dummy [386],\$dummy [387],\$dummy [388],\$dummy [389],
                  \$dummy [390],\$dummy [391],\$dummy [392],\$dummy [393]}), .BoothAddingOperand (
                  {L1_2_L2_1_G1_MINI_ALU_BoothOperand_16,
                  L1_2_L2_1_G1_MINI_ALU_BoothOperand_15,
                  L1_2_L2_1_G1_MINI_ALU_BoothOperand_14,
                  L1_2_L2_1_G1_MINI_ALU_BoothOperand_13,
                  L1_2_L2_1_G1_MINI_ALU_BoothOperand_12,
                  L1_2_L2_1_G1_MINI_ALU_BoothOperand_11,
                  L1_2_L2_1_G1_MINI_ALU_BoothOperand_10,
                  L1_2_L2_1_G1_MINI_ALU_BoothOperand_9,\$dummy [394],
                  \$dummy [395],\$dummy [396],\$dummy [397],\$dummy [398],
                  \$dummy [399],\$dummy [400],\$dummy [401],\$dummy [402]}), .BoothP (
                  {L1_2_L2_1_G1_MINI_ALU_BoothP_16,
                  L1_2_L2_1_G1_MINI_ALU_BoothP_15,
                  L1_2_L2_1_G1_MINI_ALU_BoothP_14,
                  L1_2_L2_1_G1_MINI_ALU_BoothP_13,
                  L1_2_L2_1_G1_MINI_ALU_BoothP_12,
                  L1_2_L2_1_G1_MINI_ALU_BoothP_11,
                  L1_2_L2_1_G1_MINI_ALU_BoothP_10,L1_2_L2_1_G1_MINI_ALU_BoothP_9
                  ,L1_2_L2_1_G1_MINI_ALU_BoothP_8,L1_2_L2_1_G1_MINI_ALU_BoothP_7
                  ,L1_2_L2_1_G1_MINI_ALU_BoothP_6,L1_2_L2_1_G1_MINI_ALU_BoothP_5
                  ,L1_2_L2_1_G1_MINI_ALU_BoothP_4,L1_2_L2_1_G1_MINI_ALU_BoothP_3
                  ,L1_2_L2_1_G1_MINI_ALU_BoothP_2,L1_2_L2_1_G1_MINI_ALU_BoothP_1
                  ,L1_2_L2_1_G1_MINI_ALU_BoothP_0}), .LargeWindowShifted ({
                  \$dummy [403],\$dummy [404],\$dummy [405],\$dummy [406],
                  \$dummy [407],\$dummy [408],\$dummy [409],\$dummy [410],
                  \$dummy [411],\$dummy [412],\$dummy [413],\$dummy [414],
                  \$dummy [415],\$dummy [416],\$dummy [417],\$dummy [418],
                  \$dummy [419]})) ;
    booth_adder_17_unfolded12 L1_2_L2_2_G1_MINI_ALU_BOOTH_ADDER (.AdderFirstOperand (
                              {L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16}), .AdderSecondOperand ({
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16}), .BoothOperand ({
                              L1_2_L2_2_G1_MINI_ALU_BoothOperand_16,
                              L1_2_L2_2_G1_MINI_ALU_BoothOperand_15,
                              L1_2_L2_2_G1_MINI_ALU_BoothOperand_14,
                              L1_2_L2_2_G1_MINI_ALU_BoothOperand_13,
                              L1_2_L2_2_G1_MINI_ALU_BoothOperand_12,
                              L1_2_L2_2_G1_MINI_ALU_BoothOperand_11,
                              L1_2_L2_2_G1_MINI_ALU_BoothOperand_10,
                              L1_2_L2_2_G1_MINI_ALU_BoothOperand_9,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16}), .BoothP ({
                              L1_2_L2_2_G1_MINI_ALU_BoothP_16,
                              L1_2_L2_2_G1_MINI_ALU_BoothP_15,
                              L1_2_L2_2_G1_MINI_ALU_BoothP_14,
                              L1_2_L2_2_G1_MINI_ALU_BoothP_13,
                              L1_2_L2_2_G1_MINI_ALU_BoothP_12,
                              L1_2_L2_2_G1_MINI_ALU_BoothP_11,
                              L1_2_L2_2_G1_MINI_ALU_BoothP_10,
                              L1_2_L2_2_G1_MINI_ALU_BoothP_9,
                              L1_2_L2_2_G1_MINI_ALU_BoothP_8,
                              L1_2_L2_2_G1_MINI_ALU_BoothP_7,
                              L1_2_L2_2_G1_MINI_ALU_BoothP_6,
                              L1_2_L2_2_G1_MINI_ALU_BoothP_5,
                              L1_2_L2_2_G1_MINI_ALU_BoothP_4,
                              L1_2_L2_2_G1_MINI_ALU_BoothP_3,
                              L1_2_L2_2_G1_MINI_ALU_BoothP_2,
                              L1_2_L2_2_G1_MINI_ALU_BoothP_1,
                              L1FirstOperands_12__16}), .SelOperand (nx3280), .Operation (
                              L1_2_L2_2_G1_MINI_ALU_BoothXORCheck), .AdderResult (
                              {\$dummy [420],\$dummy [421],\$dummy [422],
                              \$dummy [423],\$dummy [424],\$dummy [425],
                              \$dummy [426],\$dummy [427],\$dummy [428],
                              \$dummy [429],\$dummy [430],\$dummy [431],
                              \$dummy [432],\$dummy [433],\$dummy [434],
                              \$dummy [435],\$dummy [436]}), .AdderBoothResult (
                              {\$dummy [437],
                              L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_15,
                              L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_14,
                              L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_13,
                              L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_12,
                              L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_11,
                              L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_10,
                              L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_9,
                              L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_8,
                              L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_7,
                              L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_6,
                              L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_5,
                              L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_4,
                              L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_3,
                              L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_2,
                              L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_1,
                              L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_0})) ;
    booth_unit_17_unfolded4 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT (.CLK (CLK), .RST (
                            RST), .Start (Start), .Instr (Instr), .LoopingAndResultNotReady (
                            nx3274), .Filter ({FilterDin_2__2__7,
                            FilterDin_2__2__6,FilterDin_2__2__5,
                            FilterDin_2__2__4,FilterDin_2__2__3,
                            FilterDin_2__2__2,FilterDin_2__2__1,
                            FilterDin_2__2__0}), .Window ({WindowDin_2__2__7,
                            WindowDin_2__2__6,WindowDin_2__2__5,
                            WindowDin_2__2__4,WindowDin_2__2__3,
                            WindowDin_2__2__2,WindowDin_2__2__1,
                            WindowDin_2__2__0}), .AdderBoothResult ({
                            L1FirstOperands_12__16,
                            L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_15,
                            L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_14,
                            L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_13,
                            L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_12,
                            L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_11,
                            L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_10,
                            L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_9,
                            L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_8,
                            L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_7,
                            L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_6,
                            L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_5,
                            L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_4,
                            L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_3,
                            L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_2,
                            L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_1,
                            L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_0}), .BoothXORCheck (
                            L1_2_L2_2_G1_MINI_ALU_BoothXORCheck), .BoothResult (
                            {\$dummy [438],\$dummy [439],\$dummy [440],
                            \$dummy [441],\$dummy [442],\$dummy [443],
                            \$dummy [444],\$dummy [445]}), .BoothAddingOperand (
                            {L1_2_L2_2_G1_MINI_ALU_BoothOperand_16,
                            L1_2_L2_2_G1_MINI_ALU_BoothOperand_15,
                            L1_2_L2_2_G1_MINI_ALU_BoothOperand_14,
                            L1_2_L2_2_G1_MINI_ALU_BoothOperand_13,
                            L1_2_L2_2_G1_MINI_ALU_BoothOperand_12,
                            L1_2_L2_2_G1_MINI_ALU_BoothOperand_11,
                            L1_2_L2_2_G1_MINI_ALU_BoothOperand_10,
                            L1_2_L2_2_G1_MINI_ALU_BoothOperand_9,\$dummy [446],
                            \$dummy [447],\$dummy [448],\$dummy [449],
                            \$dummy [450],\$dummy [451],\$dummy [452],
                            \$dummy [453],\$dummy [454]}), .BoothP ({
                            L1_2_L2_2_G1_MINI_ALU_BoothP_16,
                            L1_2_L2_2_G1_MINI_ALU_BoothP_15,
                            L1_2_L2_2_G1_MINI_ALU_BoothP_14,
                            L1_2_L2_2_G1_MINI_ALU_BoothP_13,
                            L1_2_L2_2_G1_MINI_ALU_BoothP_12,
                            L1_2_L2_2_G1_MINI_ALU_BoothP_11,
                            L1_2_L2_2_G1_MINI_ALU_BoothP_10,
                            L1_2_L2_2_G1_MINI_ALU_BoothP_9,
                            L1_2_L2_2_G1_MINI_ALU_BoothP_8,
                            L1_2_L2_2_G1_MINI_ALU_BoothP_7,
                            L1_2_L2_2_G1_MINI_ALU_BoothP_6,
                            L1_2_L2_2_G1_MINI_ALU_BoothP_5,
                            L1_2_L2_2_G1_MINI_ALU_BoothP_4,
                            L1_2_L2_2_G1_MINI_ALU_BoothP_3,
                            L1_2_L2_2_G1_MINI_ALU_BoothP_2,
                            L1_2_L2_2_G1_MINI_ALU_BoothP_1,\$dummy [455]}), .LargeWindowShifted (
                            {\$dummy [456],\$dummy [457],\$dummy [458],
                            \$dummy [459],\$dummy [460],\$dummy [461],
                            \$dummy [462],\$dummy [463],\$dummy [464],
                            \$dummy [465],\$dummy [466],\$dummy [467],
                            \$dummy [468],\$dummy [469],\$dummy [470],
                            \$dummy [471],\$dummy [472]})) ;
    booth_adder_17_unfolded13 L1_2_L2_3_G2_MINI_ALU_BOOTH_ADDER (.AdderFirstOperand (
                              {L1ResultsLarge_0__16,L1ResultsLarge_0__15,
                              L1ResultsLarge_0__14,L1ResultsLarge_0__13,
                              L1ResultsLarge_0__12,L1ResultsLarge_0__11,
                              L1ResultsLarge_0__10,L1ResultsLarge_0__9,
                              L1ResultsLarge_0__8,L1ResultsLarge_0__7,
                              L1ResultsLarge_0__6,L1ResultsLarge_0__5,
                              L1ResultsLarge_0__4,L1ResultsLarge_0__3,
                              L1ResultsLarge_0__2,L1ResultsLarge_0__1,
                              L1ResultsLarge_0__0}), .AdderSecondOperand ({
                              L1ResultsLarge_1__16,L1ResultsLarge_1__15,
                              L1ResultsLarge_1__14,L1ResultsLarge_1__13,
                              L1ResultsLarge_1__12,L1ResultsLarge_1__11,
                              L1ResultsLarge_1__10,L1ResultsLarge_1__9,
                              L1ResultsLarge_1__8,L1ResultsLarge_1__7,
                              L1ResultsLarge_1__6,L1ResultsLarge_1__5,
                              L1ResultsLarge_1__4,L1ResultsLarge_1__3,
                              L1ResultsLarge_1__2,L1ResultsLarge_1__1,
                              L1ResultsLarge_1__0}), .BoothOperand ({
                              L1_2_L2_3_G2_MINI_ALU_BoothOperand_16,
                              L1_2_L2_3_G2_MINI_ALU_BoothOperand_15,
                              L1_2_L2_3_G2_MINI_ALU_BoothOperand_14,
                              L1_2_L2_3_G2_MINI_ALU_BoothOperand_13,
                              L1_2_L2_3_G2_MINI_ALU_BoothOperand_12,
                              L1_2_L2_3_G2_MINI_ALU_BoothOperand_11,
                              L1_2_L2_3_G2_MINI_ALU_BoothOperand_10,
                              L1_2_L2_3_G2_MINI_ALU_BoothOperand_9,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16}), .BoothP ({
                              L1_2_L2_3_G2_MINI_ALU_BoothP_16,
                              L1_2_L2_3_G2_MINI_ALU_BoothP_15,
                              L1_2_L2_3_G2_MINI_ALU_BoothP_14,
                              L1_2_L2_3_G2_MINI_ALU_BoothP_13,
                              L1_2_L2_3_G2_MINI_ALU_BoothP_12,
                              L1_2_L2_3_G2_MINI_ALU_BoothP_11,
                              L1_2_L2_3_G2_MINI_ALU_BoothP_10,
                              L1_2_L2_3_G2_MINI_ALU_BoothP_9,
                              L1_2_L2_3_G2_MINI_ALU_BoothP_8,
                              L1_2_L2_3_G2_MINI_ALU_BoothP_7,
                              L1_2_L2_3_G2_MINI_ALU_BoothP_6,
                              L1_2_L2_3_G2_MINI_ALU_BoothP_5,
                              L1_2_L2_3_G2_MINI_ALU_BoothP_4,
                              L1_2_L2_3_G2_MINI_ALU_BoothP_3,
                              L1_2_L2_3_G2_MINI_ALU_BoothP_2,
                              L1_2_L2_3_G2_MINI_ALU_BoothP_1,
                              L1_2_L2_3_G2_MINI_ALU_BoothP_0}), .SelOperand (
                              nx3284), .Operation (
                              L1_2_L2_3_G2_MINI_ALU_BoothXORCheck), .AdderResult (
                              {L2ResultsLarge_0__16,L2ResultsLarge_0__15,
                              L2ResultsLarge_0__14,L2ResultsLarge_0__13,
                              L2ResultsLarge_0__12,L2ResultsLarge_0__11,
                              L2ResultsLarge_0__10,L2ResultsLarge_0__9,
                              L2ResultsLarge_0__8,L2ResultsLarge_0__7,
                              L2ResultsLarge_0__6,L2ResultsLarge_0__5,
                              L2ResultsLarge_0__4,L2ResultsLarge_0__3,
                              L2ResultsLarge_0__2,L2ResultsLarge_0__1,
                              L2ResultsLarge_0__0}), .AdderBoothResult ({
                              \$dummy [473],
                              L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_15,
                              L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_14,
                              L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_13,
                              L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_12,
                              L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_11,
                              L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_10,
                              L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_9,
                              L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_8,
                              L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_7,
                              L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_6,
                              L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_5,
                              L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_4,
                              L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_3,
                              L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_2,
                              L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_1,
                              L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_0})) ;
    booth_unit_17 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT (.CLK (CLK), .RST (RST), .Start (
                  Start), .Instr (Instr), .LoopingAndResultNotReady (nx3274), .Filter (
                  {FilterDin_2__3__7,FilterDin_2__3__6,FilterDin_2__3__5,
                  FilterDin_2__3__4,FilterDin_2__3__3,FilterDin_2__3__2,
                  FilterDin_2__3__1,FilterDin_2__3__0}), .Window ({
                  WindowDin_2__3__7,WindowDin_2__3__6,WindowDin_2__3__5,
                  WindowDin_2__3__4,WindowDin_2__3__3,WindowDin_2__3__2,
                  WindowDin_2__3__1,WindowDin_2__3__0}), .AdderBoothResult ({
                  L1FirstOperands_12__16,
                  L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_15,
                  L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_14,
                  L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_13,
                  L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_12,
                  L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_11,
                  L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_10,
                  L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_9,
                  L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_8,
                  L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_7,
                  L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_6,
                  L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_5,
                  L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_4,
                  L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_3,
                  L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_2,
                  L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_1,
                  L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_0}), .BoothXORCheck (
                  L1_2_L2_3_G2_MINI_ALU_BoothXORCheck), .BoothResult ({
                  \$dummy [474],\$dummy [475],\$dummy [476],\$dummy [477],
                  \$dummy [478],\$dummy [479],\$dummy [480],\$dummy [481]}), .BoothAddingOperand (
                  {L1_2_L2_3_G2_MINI_ALU_BoothOperand_16,
                  L1_2_L2_3_G2_MINI_ALU_BoothOperand_15,
                  L1_2_L2_3_G2_MINI_ALU_BoothOperand_14,
                  L1_2_L2_3_G2_MINI_ALU_BoothOperand_13,
                  L1_2_L2_3_G2_MINI_ALU_BoothOperand_12,
                  L1_2_L2_3_G2_MINI_ALU_BoothOperand_11,
                  L1_2_L2_3_G2_MINI_ALU_BoothOperand_10,
                  L1_2_L2_3_G2_MINI_ALU_BoothOperand_9,\$dummy [482],
                  \$dummy [483],\$dummy [484],\$dummy [485],\$dummy [486],
                  \$dummy [487],\$dummy [488],\$dummy [489],\$dummy [490]}), .BoothP (
                  {L1_2_L2_3_G2_MINI_ALU_BoothP_16,
                  L1_2_L2_3_G2_MINI_ALU_BoothP_15,
                  L1_2_L2_3_G2_MINI_ALU_BoothP_14,
                  L1_2_L2_3_G2_MINI_ALU_BoothP_13,
                  L1_2_L2_3_G2_MINI_ALU_BoothP_12,
                  L1_2_L2_3_G2_MINI_ALU_BoothP_11,
                  L1_2_L2_3_G2_MINI_ALU_BoothP_10,L1_2_L2_3_G2_MINI_ALU_BoothP_9
                  ,L1_2_L2_3_G2_MINI_ALU_BoothP_8,L1_2_L2_3_G2_MINI_ALU_BoothP_7
                  ,L1_2_L2_3_G2_MINI_ALU_BoothP_6,L1_2_L2_3_G2_MINI_ALU_BoothP_5
                  ,L1_2_L2_3_G2_MINI_ALU_BoothP_4,L1_2_L2_3_G2_MINI_ALU_BoothP_3
                  ,L1_2_L2_3_G2_MINI_ALU_BoothP_2,L1_2_L2_3_G2_MINI_ALU_BoothP_1
                  ,L1_2_L2_3_G2_MINI_ALU_BoothP_0}), .LargeWindowShifted ({
                  \$dummy [491],\$dummy [492],\$dummy [493],\$dummy [494],
                  \$dummy [495],\$dummy [496],\$dummy [497],\$dummy [498],
                  \$dummy [499],\$dummy [500],\$dummy [501],\$dummy [502],
                  \$dummy [503],\$dummy [504],\$dummy [505],\$dummy [506],
                  \$dummy [507]})) ;
    booth_adder_17_unfolded13 L1_2_L2_4_G2_MINI_ALU_BOOTH_ADDER (.AdderFirstOperand (
                              {L1ResultsLarge_2__16,L1ResultsLarge_2__15,
                              L1ResultsLarge_2__14,L1ResultsLarge_2__13,
                              L1ResultsLarge_2__12,L1ResultsLarge_2__11,
                              L1ResultsLarge_2__10,L1ResultsLarge_2__9,
                              L1ResultsLarge_2__8,L1ResultsLarge_2__7,
                              L1ResultsLarge_2__6,L1ResultsLarge_2__5,
                              L1ResultsLarge_2__4,L1ResultsLarge_2__3,
                              L1ResultsLarge_2__2,L1ResultsLarge_2__1,
                              L1ResultsLarge_2__0}), .AdderSecondOperand ({
                              L1ResultsLarge_3__16,L1ResultsLarge_3__15,
                              L1ResultsLarge_3__14,L1ResultsLarge_3__13,
                              L1ResultsLarge_3__12,L1ResultsLarge_3__11,
                              L1ResultsLarge_3__10,L1ResultsLarge_3__9,
                              L1ResultsLarge_3__8,L1ResultsLarge_3__7,
                              L1ResultsLarge_3__6,L1ResultsLarge_3__5,
                              L1ResultsLarge_3__4,L1ResultsLarge_3__3,
                              L1ResultsLarge_3__2,L1ResultsLarge_3__1,
                              L1ResultsLarge_3__0}), .BoothOperand ({
                              L1_2_L2_4_G2_MINI_ALU_BoothOperand_16,
                              L1_2_L2_4_G2_MINI_ALU_BoothOperand_15,
                              L1_2_L2_4_G2_MINI_ALU_BoothOperand_14,
                              L1_2_L2_4_G2_MINI_ALU_BoothOperand_13,
                              L1_2_L2_4_G2_MINI_ALU_BoothOperand_12,
                              L1_2_L2_4_G2_MINI_ALU_BoothOperand_11,
                              L1_2_L2_4_G2_MINI_ALU_BoothOperand_10,
                              L1_2_L2_4_G2_MINI_ALU_BoothOperand_9,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16}), .BoothP ({
                              L1_2_L2_4_G2_MINI_ALU_BoothP_16,
                              L1_2_L2_4_G2_MINI_ALU_BoothP_15,
                              L1_2_L2_4_G2_MINI_ALU_BoothP_14,
                              L1_2_L2_4_G2_MINI_ALU_BoothP_13,
                              L1_2_L2_4_G2_MINI_ALU_BoothP_12,
                              L1_2_L2_4_G2_MINI_ALU_BoothP_11,
                              L1_2_L2_4_G2_MINI_ALU_BoothP_10,
                              L1_2_L2_4_G2_MINI_ALU_BoothP_9,
                              L1_2_L2_4_G2_MINI_ALU_BoothP_8,
                              L1_2_L2_4_G2_MINI_ALU_BoothP_7,
                              L1_2_L2_4_G2_MINI_ALU_BoothP_6,
                              L1_2_L2_4_G2_MINI_ALU_BoothP_5,
                              L1_2_L2_4_G2_MINI_ALU_BoothP_4,
                              L1_2_L2_4_G2_MINI_ALU_BoothP_3,
                              L1_2_L2_4_G2_MINI_ALU_BoothP_2,
                              L1_2_L2_4_G2_MINI_ALU_BoothP_1,
                              L1_2_L2_4_G2_MINI_ALU_BoothP_0}), .SelOperand (
                              nx3284), .Operation (
                              L1_2_L2_4_G2_MINI_ALU_BoothXORCheck), .AdderResult (
                              {L2ResultsLarge_1__16,L2ResultsLarge_1__15,
                              L2ResultsLarge_1__14,L2ResultsLarge_1__13,
                              L2ResultsLarge_1__12,L2ResultsLarge_1__11,
                              L2ResultsLarge_1__10,L2ResultsLarge_1__9,
                              L2ResultsLarge_1__8,L2ResultsLarge_1__7,
                              L2ResultsLarge_1__6,L2ResultsLarge_1__5,
                              L2ResultsLarge_1__4,L2ResultsLarge_1__3,
                              L2ResultsLarge_1__2,L2ResultsLarge_1__1,
                              L2ResultsLarge_1__0}), .AdderBoothResult ({
                              \$dummy [508],
                              L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_15,
                              L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_14,
                              L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_13,
                              L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_12,
                              L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_11,
                              L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_10,
                              L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_9,
                              L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_8,
                              L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_7,
                              L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_6,
                              L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_5,
                              L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_4,
                              L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_3,
                              L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_2,
                              L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_1,
                              L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_0})) ;
    booth_unit_17 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT (.CLK (CLK), .RST (RST), .Start (
                  Start), .Instr (Instr), .LoopingAndResultNotReady (nx3276), .Filter (
                  {FilterDin_2__4__7,FilterDin_2__4__6,FilterDin_2__4__5,
                  FilterDin_2__4__4,FilterDin_2__4__3,FilterDin_2__4__2,
                  FilterDin_2__4__1,FilterDin_2__4__0}), .Window ({
                  WindowDin_2__4__7,WindowDin_2__4__6,WindowDin_2__4__5,
                  WindowDin_2__4__4,WindowDin_2__4__3,WindowDin_2__4__2,
                  WindowDin_2__4__1,WindowDin_2__4__0}), .AdderBoothResult ({
                  L1FirstOperands_12__16,
                  L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_15,
                  L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_14,
                  L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_13,
                  L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_12,
                  L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_11,
                  L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_10,
                  L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_9,
                  L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_8,
                  L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_7,
                  L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_6,
                  L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_5,
                  L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_4,
                  L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_3,
                  L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_2,
                  L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_1,
                  L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_0}), .BoothXORCheck (
                  L1_2_L2_4_G2_MINI_ALU_BoothXORCheck), .BoothResult ({
                  \$dummy [509],\$dummy [510],\$dummy [511],\$dummy [512],
                  \$dummy [513],\$dummy [514],\$dummy [515],\$dummy [516]}), .BoothAddingOperand (
                  {L1_2_L2_4_G2_MINI_ALU_BoothOperand_16,
                  L1_2_L2_4_G2_MINI_ALU_BoothOperand_15,
                  L1_2_L2_4_G2_MINI_ALU_BoothOperand_14,
                  L1_2_L2_4_G2_MINI_ALU_BoothOperand_13,
                  L1_2_L2_4_G2_MINI_ALU_BoothOperand_12,
                  L1_2_L2_4_G2_MINI_ALU_BoothOperand_11,
                  L1_2_L2_4_G2_MINI_ALU_BoothOperand_10,
                  L1_2_L2_4_G2_MINI_ALU_BoothOperand_9,\$dummy [517],
                  \$dummy [518],\$dummy [519],\$dummy [520],\$dummy [521],
                  \$dummy [522],\$dummy [523],\$dummy [524],\$dummy [525]}), .BoothP (
                  {L1_2_L2_4_G2_MINI_ALU_BoothP_16,
                  L1_2_L2_4_G2_MINI_ALU_BoothP_15,
                  L1_2_L2_4_G2_MINI_ALU_BoothP_14,
                  L1_2_L2_4_G2_MINI_ALU_BoothP_13,
                  L1_2_L2_4_G2_MINI_ALU_BoothP_12,
                  L1_2_L2_4_G2_MINI_ALU_BoothP_11,
                  L1_2_L2_4_G2_MINI_ALU_BoothP_10,L1_2_L2_4_G2_MINI_ALU_BoothP_9
                  ,L1_2_L2_4_G2_MINI_ALU_BoothP_8,L1_2_L2_4_G2_MINI_ALU_BoothP_7
                  ,L1_2_L2_4_G2_MINI_ALU_BoothP_6,L1_2_L2_4_G2_MINI_ALU_BoothP_5
                  ,L1_2_L2_4_G2_MINI_ALU_BoothP_4,L1_2_L2_4_G2_MINI_ALU_BoothP_3
                  ,L1_2_L2_4_G2_MINI_ALU_BoothP_2,L1_2_L2_4_G2_MINI_ALU_BoothP_1
                  ,L1_2_L2_4_G2_MINI_ALU_BoothP_0}), .LargeWindowShifted ({
                  \$dummy [526],\$dummy [527],\$dummy [528],\$dummy [529],
                  \$dummy [530],\$dummy [531],\$dummy [532],\$dummy [533],
                  \$dummy [534],\$dummy [535],\$dummy [536],\$dummy [537],
                  \$dummy [538],\$dummy [539],\$dummy [540],\$dummy [541],
                  \$dummy [542]})) ;
    booth_adder_17_unfolded13 L1_3_L2_0_G2_MINI_ALU_BOOTH_ADDER (.AdderFirstOperand (
                              {L1ResultsLarge_4__16,L1ResultsLarge_4__15,
                              L1ResultsLarge_4__14,L1ResultsLarge_4__13,
                              L1ResultsLarge_4__12,L1ResultsLarge_4__11,
                              L1ResultsLarge_4__10,L1ResultsLarge_4__9,
                              L1ResultsLarge_4__8,L1ResultsLarge_4__7,
                              L1ResultsLarge_4__6,L1ResultsLarge_4__5,
                              L1ResultsLarge_4__4,L1ResultsLarge_4__3,
                              L1ResultsLarge_4__2,L1ResultsLarge_4__1,
                              L1ResultsLarge_4__0}), .AdderSecondOperand ({
                              L1ResultsLarge_5__16,L1ResultsLarge_5__15,
                              L1ResultsLarge_5__14,L1ResultsLarge_5__13,
                              L1ResultsLarge_5__12,L1ResultsLarge_5__11,
                              L1ResultsLarge_5__10,L1ResultsLarge_5__9,
                              L1ResultsLarge_5__8,L1ResultsLarge_5__7,
                              L1ResultsLarge_5__6,L1ResultsLarge_5__5,
                              L1ResultsLarge_5__4,L1ResultsLarge_5__3,
                              L1ResultsLarge_5__2,L1ResultsLarge_5__1,
                              L1ResultsLarge_5__0}), .BoothOperand ({
                              L1_3_L2_0_G2_MINI_ALU_BoothOperand_16,
                              L1_3_L2_0_G2_MINI_ALU_BoothOperand_15,
                              L1_3_L2_0_G2_MINI_ALU_BoothOperand_14,
                              L1_3_L2_0_G2_MINI_ALU_BoothOperand_13,
                              L1_3_L2_0_G2_MINI_ALU_BoothOperand_12,
                              L1_3_L2_0_G2_MINI_ALU_BoothOperand_11,
                              L1_3_L2_0_G2_MINI_ALU_BoothOperand_10,
                              L1_3_L2_0_G2_MINI_ALU_BoothOperand_9,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16}), .BoothP ({
                              L1_3_L2_0_G2_MINI_ALU_BoothP_16,
                              L1_3_L2_0_G2_MINI_ALU_BoothP_15,
                              L1_3_L2_0_G2_MINI_ALU_BoothP_14,
                              L1_3_L2_0_G2_MINI_ALU_BoothP_13,
                              L1_3_L2_0_G2_MINI_ALU_BoothP_12,
                              L1_3_L2_0_G2_MINI_ALU_BoothP_11,
                              L1_3_L2_0_G2_MINI_ALU_BoothP_10,
                              L1_3_L2_0_G2_MINI_ALU_BoothP_9,
                              L1_3_L2_0_G2_MINI_ALU_BoothP_8,
                              L1_3_L2_0_G2_MINI_ALU_BoothP_7,
                              L1_3_L2_0_G2_MINI_ALU_BoothP_6,
                              L1_3_L2_0_G2_MINI_ALU_BoothP_5,
                              L1_3_L2_0_G2_MINI_ALU_BoothP_4,
                              L1_3_L2_0_G2_MINI_ALU_BoothP_3,
                              L1_3_L2_0_G2_MINI_ALU_BoothP_2,
                              L1_3_L2_0_G2_MINI_ALU_BoothP_1,
                              L1_3_L2_0_G2_MINI_ALU_BoothP_0}), .SelOperand (
                              nx3284), .Operation (
                              L1_3_L2_0_G2_MINI_ALU_BoothXORCheck), .AdderResult (
                              {L2ResultsLarge_2__16,L2ResultsLarge_2__15,
                              L2ResultsLarge_2__14,L2ResultsLarge_2__13,
                              L2ResultsLarge_2__12,L2ResultsLarge_2__11,
                              L2ResultsLarge_2__10,L2ResultsLarge_2__9,
                              L2ResultsLarge_2__8,L2ResultsLarge_2__7,
                              L2ResultsLarge_2__6,L2ResultsLarge_2__5,
                              L2ResultsLarge_2__4,L2ResultsLarge_2__3,
                              L2ResultsLarge_2__2,L2ResultsLarge_2__1,
                              L2ResultsLarge_2__0}), .AdderBoothResult ({
                              \$dummy [543],
                              L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_15,
                              L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_14,
                              L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_13,
                              L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_12,
                              L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_11,
                              L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_10,
                              L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_9,
                              L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_8,
                              L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_7,
                              L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_6,
                              L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_5,
                              L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_4,
                              L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_3,
                              L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_2,
                              L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_1,
                              L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_0})) ;
    booth_unit_17 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT (.CLK (CLK), .RST (RST), .Start (
                  Start), .Instr (Instr), .LoopingAndResultNotReady (nx3276), .Filter (
                  {FilterDin_3__0__7,FilterDin_3__0__6,FilterDin_3__0__5,
                  FilterDin_3__0__4,FilterDin_3__0__3,FilterDin_3__0__2,
                  FilterDin_3__0__1,FilterDin_3__0__0}), .Window ({
                  WindowDin_3__0__7,WindowDin_3__0__6,WindowDin_3__0__5,
                  WindowDin_3__0__4,WindowDin_3__0__3,WindowDin_3__0__2,
                  WindowDin_3__0__1,WindowDin_3__0__0}), .AdderBoothResult ({
                  L1FirstOperands_12__16,
                  L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_15,
                  L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_14,
                  L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_13,
                  L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_12,
                  L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_11,
                  L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_10,
                  L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_9,
                  L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_8,
                  L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_7,
                  L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_6,
                  L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_5,
                  L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_4,
                  L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_3,
                  L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_2,
                  L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_1,
                  L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_0}), .BoothXORCheck (
                  L1_3_L2_0_G2_MINI_ALU_BoothXORCheck), .BoothResult ({
                  \$dummy [544],\$dummy [545],\$dummy [546],\$dummy [547],
                  \$dummy [548],\$dummy [549],\$dummy [550],\$dummy [551]}), .BoothAddingOperand (
                  {L1_3_L2_0_G2_MINI_ALU_BoothOperand_16,
                  L1_3_L2_0_G2_MINI_ALU_BoothOperand_15,
                  L1_3_L2_0_G2_MINI_ALU_BoothOperand_14,
                  L1_3_L2_0_G2_MINI_ALU_BoothOperand_13,
                  L1_3_L2_0_G2_MINI_ALU_BoothOperand_12,
                  L1_3_L2_0_G2_MINI_ALU_BoothOperand_11,
                  L1_3_L2_0_G2_MINI_ALU_BoothOperand_10,
                  L1_3_L2_0_G2_MINI_ALU_BoothOperand_9,\$dummy [552],
                  \$dummy [553],\$dummy [554],\$dummy [555],\$dummy [556],
                  \$dummy [557],\$dummy [558],\$dummy [559],\$dummy [560]}), .BoothP (
                  {L1_3_L2_0_G2_MINI_ALU_BoothP_16,
                  L1_3_L2_0_G2_MINI_ALU_BoothP_15,
                  L1_3_L2_0_G2_MINI_ALU_BoothP_14,
                  L1_3_L2_0_G2_MINI_ALU_BoothP_13,
                  L1_3_L2_0_G2_MINI_ALU_BoothP_12,
                  L1_3_L2_0_G2_MINI_ALU_BoothP_11,
                  L1_3_L2_0_G2_MINI_ALU_BoothP_10,L1_3_L2_0_G2_MINI_ALU_BoothP_9
                  ,L1_3_L2_0_G2_MINI_ALU_BoothP_8,L1_3_L2_0_G2_MINI_ALU_BoothP_7
                  ,L1_3_L2_0_G2_MINI_ALU_BoothP_6,L1_3_L2_0_G2_MINI_ALU_BoothP_5
                  ,L1_3_L2_0_G2_MINI_ALU_BoothP_4,L1_3_L2_0_G2_MINI_ALU_BoothP_3
                  ,L1_3_L2_0_G2_MINI_ALU_BoothP_2,L1_3_L2_0_G2_MINI_ALU_BoothP_1
                  ,L1_3_L2_0_G2_MINI_ALU_BoothP_0}), .LargeWindowShifted ({
                  \$dummy [561],\$dummy [562],\$dummy [563],\$dummy [564],
                  \$dummy [565],\$dummy [566],\$dummy [567],\$dummy [568],
                  \$dummy [569],\$dummy [570],\$dummy [571],\$dummy [572],
                  \$dummy [573],\$dummy [574],\$dummy [575],\$dummy [576],
                  \$dummy [577]})) ;
    booth_adder_17_unfolded13 L1_3_L2_1_G2_MINI_ALU_BOOTH_ADDER (.AdderFirstOperand (
                              {L1ResultsLarge_6__16,L1ResultsLarge_6__15,
                              L1ResultsLarge_6__14,L1ResultsLarge_6__13,
                              L1ResultsLarge_6__12,L1ResultsLarge_6__11,
                              L1ResultsLarge_6__10,L1ResultsLarge_6__9,
                              L1ResultsLarge_6__8,L1ResultsLarge_6__7,
                              L1ResultsLarge_6__6,L1ResultsLarge_6__5,
                              L1ResultsLarge_6__4,L1ResultsLarge_6__3,
                              L1ResultsLarge_6__2,L1ResultsLarge_6__1,
                              L1ResultsLarge_6__0}), .AdderSecondOperand ({
                              L1ResultsLarge_7__16,L1ResultsLarge_7__15,
                              L1ResultsLarge_7__14,L1ResultsLarge_7__13,
                              L1ResultsLarge_7__12,L1ResultsLarge_7__11,
                              L1ResultsLarge_7__10,L1ResultsLarge_7__9,
                              L1ResultsLarge_7__8,L1ResultsLarge_7__7,
                              L1ResultsLarge_7__6,L1ResultsLarge_7__5,
                              L1ResultsLarge_7__4,L1ResultsLarge_7__3,
                              L1ResultsLarge_7__2,L1ResultsLarge_7__1,
                              L1ResultsLarge_7__0}), .BoothOperand ({
                              L1_3_L2_1_G2_MINI_ALU_BoothOperand_16,
                              L1_3_L2_1_G2_MINI_ALU_BoothOperand_15,
                              L1_3_L2_1_G2_MINI_ALU_BoothOperand_14,
                              L1_3_L2_1_G2_MINI_ALU_BoothOperand_13,
                              L1_3_L2_1_G2_MINI_ALU_BoothOperand_12,
                              L1_3_L2_1_G2_MINI_ALU_BoothOperand_11,
                              L1_3_L2_1_G2_MINI_ALU_BoothOperand_10,
                              L1_3_L2_1_G2_MINI_ALU_BoothOperand_9,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16}), .BoothP ({
                              L1_3_L2_1_G2_MINI_ALU_BoothP_16,
                              L1_3_L2_1_G2_MINI_ALU_BoothP_15,
                              L1_3_L2_1_G2_MINI_ALU_BoothP_14,
                              L1_3_L2_1_G2_MINI_ALU_BoothP_13,
                              L1_3_L2_1_G2_MINI_ALU_BoothP_12,
                              L1_3_L2_1_G2_MINI_ALU_BoothP_11,
                              L1_3_L2_1_G2_MINI_ALU_BoothP_10,
                              L1_3_L2_1_G2_MINI_ALU_BoothP_9,
                              L1_3_L2_1_G2_MINI_ALU_BoothP_8,
                              L1_3_L2_1_G2_MINI_ALU_BoothP_7,
                              L1_3_L2_1_G2_MINI_ALU_BoothP_6,
                              L1_3_L2_1_G2_MINI_ALU_BoothP_5,
                              L1_3_L2_1_G2_MINI_ALU_BoothP_4,
                              L1_3_L2_1_G2_MINI_ALU_BoothP_3,
                              L1_3_L2_1_G2_MINI_ALU_BoothP_2,
                              L1_3_L2_1_G2_MINI_ALU_BoothP_1,
                              L1_3_L2_1_G2_MINI_ALU_BoothP_0}), .SelOperand (
                              nx3282), .Operation (
                              L1_3_L2_1_G2_MINI_ALU_BoothXORCheck), .AdderResult (
                              {L2ResultsLarge_3__16,L2ResultsLarge_3__15,
                              L2ResultsLarge_3__14,L2ResultsLarge_3__13,
                              L2ResultsLarge_3__12,L2ResultsLarge_3__11,
                              L2ResultsLarge_3__10,L2ResultsLarge_3__9,
                              L2ResultsLarge_3__8,L2ResultsLarge_3__7,
                              L2ResultsLarge_3__6,L2ResultsLarge_3__5,
                              L2ResultsLarge_3__4,L2ResultsLarge_3__3,
                              L2ResultsLarge_3__2,L2ResultsLarge_3__1,
                              L2ResultsLarge_3__0}), .AdderBoothResult ({
                              \$dummy [578],
                              L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_15,
                              L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_14,
                              L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_13,
                              L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_12,
                              L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_11,
                              L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_10,
                              L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_9,
                              L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_8,
                              L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_7,
                              L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_6,
                              L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_5,
                              L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_4,
                              L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_3,
                              L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_2,
                              L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_1,
                              L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_0})) ;
    booth_unit_17 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT (.CLK (CLK), .RST (RST), .Start (
                  Start), .Instr (Instr), .LoopingAndResultNotReady (nx3276), .Filter (
                  {FilterDin_3__1__7,FilterDin_3__1__6,FilterDin_3__1__5,
                  FilterDin_3__1__4,FilterDin_3__1__3,FilterDin_3__1__2,
                  FilterDin_3__1__1,FilterDin_3__1__0}), .Window ({
                  WindowDin_3__1__7,WindowDin_3__1__6,WindowDin_3__1__5,
                  WindowDin_3__1__4,WindowDin_3__1__3,WindowDin_3__1__2,
                  WindowDin_3__1__1,WindowDin_3__1__0}), .AdderBoothResult ({
                  L1FirstOperands_12__16,
                  L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_15,
                  L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_14,
                  L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_13,
                  L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_12,
                  L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_11,
                  L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_10,
                  L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_9,
                  L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_8,
                  L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_7,
                  L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_6,
                  L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_5,
                  L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_4,
                  L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_3,
                  L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_2,
                  L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_1,
                  L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_0}), .BoothXORCheck (
                  L1_3_L2_1_G2_MINI_ALU_BoothXORCheck), .BoothResult ({
                  \$dummy [579],\$dummy [580],\$dummy [581],\$dummy [582],
                  \$dummy [583],\$dummy [584],\$dummy [585],\$dummy [586]}), .BoothAddingOperand (
                  {L1_3_L2_1_G2_MINI_ALU_BoothOperand_16,
                  L1_3_L2_1_G2_MINI_ALU_BoothOperand_15,
                  L1_3_L2_1_G2_MINI_ALU_BoothOperand_14,
                  L1_3_L2_1_G2_MINI_ALU_BoothOperand_13,
                  L1_3_L2_1_G2_MINI_ALU_BoothOperand_12,
                  L1_3_L2_1_G2_MINI_ALU_BoothOperand_11,
                  L1_3_L2_1_G2_MINI_ALU_BoothOperand_10,
                  L1_3_L2_1_G2_MINI_ALU_BoothOperand_9,\$dummy [587],
                  \$dummy [588],\$dummy [589],\$dummy [590],\$dummy [591],
                  \$dummy [592],\$dummy [593],\$dummy [594],\$dummy [595]}), .BoothP (
                  {L1_3_L2_1_G2_MINI_ALU_BoothP_16,
                  L1_3_L2_1_G2_MINI_ALU_BoothP_15,
                  L1_3_L2_1_G2_MINI_ALU_BoothP_14,
                  L1_3_L2_1_G2_MINI_ALU_BoothP_13,
                  L1_3_L2_1_G2_MINI_ALU_BoothP_12,
                  L1_3_L2_1_G2_MINI_ALU_BoothP_11,
                  L1_3_L2_1_G2_MINI_ALU_BoothP_10,L1_3_L2_1_G2_MINI_ALU_BoothP_9
                  ,L1_3_L2_1_G2_MINI_ALU_BoothP_8,L1_3_L2_1_G2_MINI_ALU_BoothP_7
                  ,L1_3_L2_1_G2_MINI_ALU_BoothP_6,L1_3_L2_1_G2_MINI_ALU_BoothP_5
                  ,L1_3_L2_1_G2_MINI_ALU_BoothP_4,L1_3_L2_1_G2_MINI_ALU_BoothP_3
                  ,L1_3_L2_1_G2_MINI_ALU_BoothP_2,L1_3_L2_1_G2_MINI_ALU_BoothP_1
                  ,L1_3_L2_1_G2_MINI_ALU_BoothP_0}), .LargeWindowShifted ({
                  \$dummy [596],\$dummy [597],\$dummy [598],\$dummy [599],
                  \$dummy [600],\$dummy [601],\$dummy [602],\$dummy [603],
                  \$dummy [604],\$dummy [605],\$dummy [606],\$dummy [607],
                  \$dummy [608],\$dummy [609],\$dummy [610],\$dummy [611],
                  \$dummy [612]})) ;
    booth_adder_17_unfolded13 L1_3_L2_2_G2_MINI_ALU_BOOTH_ADDER (.AdderFirstOperand (
                              {L1ResultsLarge_8__16,L1ResultsLarge_8__15,
                              L1ResultsLarge_8__14,L1ResultsLarge_8__13,
                              L1ResultsLarge_8__12,L1ResultsLarge_8__11,
                              L1ResultsLarge_8__10,L1ResultsLarge_8__9,
                              L1ResultsLarge_8__8,L1ResultsLarge_8__7,
                              L1ResultsLarge_8__6,L1ResultsLarge_8__5,
                              L1ResultsLarge_8__4,L1ResultsLarge_8__3,
                              L1ResultsLarge_8__2,L1ResultsLarge_8__1,
                              L1ResultsLarge_8__0}), .AdderSecondOperand ({
                              L1ResultsLarge_9__16,L1ResultsLarge_9__15,
                              L1ResultsLarge_9__14,L1ResultsLarge_9__13,
                              L1ResultsLarge_9__12,L1ResultsLarge_9__11,
                              L1ResultsLarge_9__10,L1ResultsLarge_9__9,
                              L1ResultsLarge_9__8,L1ResultsLarge_9__7,
                              L1ResultsLarge_9__6,L1ResultsLarge_9__5,
                              L1ResultsLarge_9__4,L1ResultsLarge_9__3,
                              L1ResultsLarge_9__2,L1ResultsLarge_9__1,
                              L1ResultsLarge_9__0}), .BoothOperand ({
                              L1_3_L2_2_G2_MINI_ALU_BoothOperand_16,
                              L1_3_L2_2_G2_MINI_ALU_BoothOperand_15,
                              L1_3_L2_2_G2_MINI_ALU_BoothOperand_14,
                              L1_3_L2_2_G2_MINI_ALU_BoothOperand_13,
                              L1_3_L2_2_G2_MINI_ALU_BoothOperand_12,
                              L1_3_L2_2_G2_MINI_ALU_BoothOperand_11,
                              L1_3_L2_2_G2_MINI_ALU_BoothOperand_10,
                              L1_3_L2_2_G2_MINI_ALU_BoothOperand_9,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16}), .BoothP ({
                              L1_3_L2_2_G2_MINI_ALU_BoothP_16,
                              L1_3_L2_2_G2_MINI_ALU_BoothP_15,
                              L1_3_L2_2_G2_MINI_ALU_BoothP_14,
                              L1_3_L2_2_G2_MINI_ALU_BoothP_13,
                              L1_3_L2_2_G2_MINI_ALU_BoothP_12,
                              L1_3_L2_2_G2_MINI_ALU_BoothP_11,
                              L1_3_L2_2_G2_MINI_ALU_BoothP_10,
                              L1_3_L2_2_G2_MINI_ALU_BoothP_9,
                              L1_3_L2_2_G2_MINI_ALU_BoothP_8,
                              L1_3_L2_2_G2_MINI_ALU_BoothP_7,
                              L1_3_L2_2_G2_MINI_ALU_BoothP_6,
                              L1_3_L2_2_G2_MINI_ALU_BoothP_5,
                              L1_3_L2_2_G2_MINI_ALU_BoothP_4,
                              L1_3_L2_2_G2_MINI_ALU_BoothP_3,
                              L1_3_L2_2_G2_MINI_ALU_BoothP_2,
                              L1_3_L2_2_G2_MINI_ALU_BoothP_1,
                              L1_3_L2_2_G2_MINI_ALU_BoothP_0}), .SelOperand (
                              nx3284), .Operation (
                              L1_3_L2_2_G2_MINI_ALU_BoothXORCheck), .AdderResult (
                              {L2ResultsLarge_4__16,L2ResultsLarge_4__15,
                              L2ResultsLarge_4__14,L2ResultsLarge_4__13,
                              L2ResultsLarge_4__12,L2ResultsLarge_4__11,
                              L2ResultsLarge_4__10,L2ResultsLarge_4__9,
                              L2ResultsLarge_4__8,L2ResultsLarge_4__7,
                              L2ResultsLarge_4__6,L2ResultsLarge_4__5,
                              L2ResultsLarge_4__4,L2ResultsLarge_4__3,
                              L2ResultsLarge_4__2,L2ResultsLarge_4__1,
                              L2ResultsLarge_4__0}), .AdderBoothResult ({
                              \$dummy [613],
                              L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_15,
                              L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_14,
                              L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_13,
                              L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_12,
                              L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_11,
                              L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_10,
                              L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_9,
                              L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_8,
                              L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_7,
                              L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_6,
                              L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_5,
                              L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_4,
                              L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_3,
                              L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_2,
                              L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_1,
                              L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_0})) ;
    booth_unit_17 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT (.CLK (CLK), .RST (RST), .Start (
                  Start), .Instr (Instr), .LoopingAndResultNotReady (nx3276), .Filter (
                  {FilterDin_3__2__7,FilterDin_3__2__6,FilterDin_3__2__5,
                  FilterDin_3__2__4,FilterDin_3__2__3,FilterDin_3__2__2,
                  FilterDin_3__2__1,FilterDin_3__2__0}), .Window ({
                  WindowDin_3__2__7,WindowDin_3__2__6,WindowDin_3__2__5,
                  WindowDin_3__2__4,WindowDin_3__2__3,WindowDin_3__2__2,
                  WindowDin_3__2__1,WindowDin_3__2__0}), .AdderBoothResult ({
                  L1FirstOperands_12__16,
                  L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_15,
                  L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_14,
                  L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_13,
                  L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_12,
                  L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_11,
                  L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_10,
                  L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_9,
                  L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_8,
                  L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_7,
                  L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_6,
                  L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_5,
                  L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_4,
                  L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_3,
                  L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_2,
                  L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_1,
                  L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_0}), .BoothXORCheck (
                  L1_3_L2_2_G2_MINI_ALU_BoothXORCheck), .BoothResult ({
                  \$dummy [614],\$dummy [615],\$dummy [616],\$dummy [617],
                  \$dummy [618],\$dummy [619],\$dummy [620],\$dummy [621]}), .BoothAddingOperand (
                  {L1_3_L2_2_G2_MINI_ALU_BoothOperand_16,
                  L1_3_L2_2_G2_MINI_ALU_BoothOperand_15,
                  L1_3_L2_2_G2_MINI_ALU_BoothOperand_14,
                  L1_3_L2_2_G2_MINI_ALU_BoothOperand_13,
                  L1_3_L2_2_G2_MINI_ALU_BoothOperand_12,
                  L1_3_L2_2_G2_MINI_ALU_BoothOperand_11,
                  L1_3_L2_2_G2_MINI_ALU_BoothOperand_10,
                  L1_3_L2_2_G2_MINI_ALU_BoothOperand_9,\$dummy [622],
                  \$dummy [623],\$dummy [624],\$dummy [625],\$dummy [626],
                  \$dummy [627],\$dummy [628],\$dummy [629],\$dummy [630]}), .BoothP (
                  {L1_3_L2_2_G2_MINI_ALU_BoothP_16,
                  L1_3_L2_2_G2_MINI_ALU_BoothP_15,
                  L1_3_L2_2_G2_MINI_ALU_BoothP_14,
                  L1_3_L2_2_G2_MINI_ALU_BoothP_13,
                  L1_3_L2_2_G2_MINI_ALU_BoothP_12,
                  L1_3_L2_2_G2_MINI_ALU_BoothP_11,
                  L1_3_L2_2_G2_MINI_ALU_BoothP_10,L1_3_L2_2_G2_MINI_ALU_BoothP_9
                  ,L1_3_L2_2_G2_MINI_ALU_BoothP_8,L1_3_L2_2_G2_MINI_ALU_BoothP_7
                  ,L1_3_L2_2_G2_MINI_ALU_BoothP_6,L1_3_L2_2_G2_MINI_ALU_BoothP_5
                  ,L1_3_L2_2_G2_MINI_ALU_BoothP_4,L1_3_L2_2_G2_MINI_ALU_BoothP_3
                  ,L1_3_L2_2_G2_MINI_ALU_BoothP_2,L1_3_L2_2_G2_MINI_ALU_BoothP_1
                  ,L1_3_L2_2_G2_MINI_ALU_BoothP_0}), .LargeWindowShifted ({
                  \$dummy [631],\$dummy [632],\$dummy [633],\$dummy [634],
                  \$dummy [635],\$dummy [636],\$dummy [637],\$dummy [638],
                  \$dummy [639],\$dummy [640],\$dummy [641],\$dummy [642],
                  \$dummy [643],\$dummy [644],\$dummy [645],\$dummy [646],
                  \$dummy [647]})) ;
    booth_adder_17_unfolded13 L1_3_L2_3_G2_MINI_ALU_BOOTH_ADDER (.AdderFirstOperand (
                              {L1ResultsLarge_10__16,L1ResultsLarge_10__15,
                              L1ResultsLarge_10__14,L1ResultsLarge_10__13,
                              L1ResultsLarge_10__12,L1ResultsLarge_10__11,
                              L1ResultsLarge_10__10,L1ResultsLarge_10__9,
                              L1ResultsLarge_10__8,L1ResultsLarge_10__7,
                              L1ResultsLarge_10__6,L1ResultsLarge_10__5,
                              L1ResultsLarge_10__4,L1ResultsLarge_10__3,
                              L1ResultsLarge_10__2,L1ResultsLarge_10__1,
                              L1ResultsLarge_10__0}), .AdderSecondOperand ({
                              L1ResultsLarge_11__16,L1ResultsLarge_11__15,
                              L1ResultsLarge_11__14,L1ResultsLarge_11__13,
                              L1ResultsLarge_11__12,L1ResultsLarge_11__11,
                              L1ResultsLarge_11__10,L1ResultsLarge_11__9,
                              L1ResultsLarge_11__8,L1ResultsLarge_11__7,
                              L1ResultsLarge_11__6,L1ResultsLarge_11__5,
                              L1ResultsLarge_11__4,L1ResultsLarge_11__3,
                              L1ResultsLarge_11__2,L1ResultsLarge_11__1,
                              L1ResultsLarge_11__0}), .BoothOperand ({
                              L1_3_L2_3_G2_MINI_ALU_BoothOperand_16,
                              L1_3_L2_3_G2_MINI_ALU_BoothOperand_15,
                              L1_3_L2_3_G2_MINI_ALU_BoothOperand_14,
                              L1_3_L2_3_G2_MINI_ALU_BoothOperand_13,
                              L1_3_L2_3_G2_MINI_ALU_BoothOperand_12,
                              L1_3_L2_3_G2_MINI_ALU_BoothOperand_11,
                              L1_3_L2_3_G2_MINI_ALU_BoothOperand_10,
                              L1_3_L2_3_G2_MINI_ALU_BoothOperand_9,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16}), .BoothP ({
                              L1_3_L2_3_G2_MINI_ALU_BoothP_16,
                              L1_3_L2_3_G2_MINI_ALU_BoothP_15,
                              L1_3_L2_3_G2_MINI_ALU_BoothP_14,
                              L1_3_L2_3_G2_MINI_ALU_BoothP_13,
                              L1_3_L2_3_G2_MINI_ALU_BoothP_12,
                              L1_3_L2_3_G2_MINI_ALU_BoothP_11,
                              L1_3_L2_3_G2_MINI_ALU_BoothP_10,
                              L1_3_L2_3_G2_MINI_ALU_BoothP_9,
                              L1_3_L2_3_G2_MINI_ALU_BoothP_8,
                              L1_3_L2_3_G2_MINI_ALU_BoothP_7,
                              L1_3_L2_3_G2_MINI_ALU_BoothP_6,
                              L1_3_L2_3_G2_MINI_ALU_BoothP_5,
                              L1_3_L2_3_G2_MINI_ALU_BoothP_4,
                              L1_3_L2_3_G2_MINI_ALU_BoothP_3,
                              L1_3_L2_3_G2_MINI_ALU_BoothP_2,
                              L1_3_L2_3_G2_MINI_ALU_BoothP_1,
                              L1_3_L2_3_G2_MINI_ALU_BoothP_0}), .SelOperand (
                              nx3284), .Operation (
                              L1_3_L2_3_G2_MINI_ALU_BoothXORCheck), .AdderResult (
                              {L2ResultsLarge_5__16,L2ResultsLarge_5__15,
                              L2ResultsLarge_5__14,L2ResultsLarge_5__13,
                              L2ResultsLarge_5__12,L2ResultsLarge_5__11,
                              L2ResultsLarge_5__10,L2ResultsLarge_5__9,
                              L2ResultsLarge_5__8,L2ResultsLarge_5__7,
                              L2ResultsLarge_5__6,L2ResultsLarge_5__5,
                              L2ResultsLarge_5__4,L2ResultsLarge_5__3,
                              L2ResultsLarge_5__2,L2ResultsLarge_5__1,
                              L2ResultsLarge_5__0}), .AdderBoothResult ({
                              \$dummy [648],
                              L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_15,
                              L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_14,
                              L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_13,
                              L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_12,
                              L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_11,
                              L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_10,
                              L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_9,
                              L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_8,
                              L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_7,
                              L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_6,
                              L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_5,
                              L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_4,
                              L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_3,
                              L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_2,
                              L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_1,
                              L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_0})) ;
    booth_unit_17 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT (.CLK (CLK), .RST (RST), .Start (
                  Start), .Instr (Instr), .LoopingAndResultNotReady (nx3276), .Filter (
                  {FilterDin_3__3__7,FilterDin_3__3__6,FilterDin_3__3__5,
                  FilterDin_3__3__4,FilterDin_3__3__3,FilterDin_3__3__2,
                  FilterDin_3__3__1,FilterDin_3__3__0}), .Window ({
                  WindowDin_3__3__7,WindowDin_3__3__6,WindowDin_3__3__5,
                  WindowDin_3__3__4,WindowDin_3__3__3,WindowDin_3__3__2,
                  WindowDin_3__3__1,WindowDin_3__3__0}), .AdderBoothResult ({
                  L1FirstOperands_12__16,
                  L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_15,
                  L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_14,
                  L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_13,
                  L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_12,
                  L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_11,
                  L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_10,
                  L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_9,
                  L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_8,
                  L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_7,
                  L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_6,
                  L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_5,
                  L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_4,
                  L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_3,
                  L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_2,
                  L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_1,
                  L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_0}), .BoothXORCheck (
                  L1_3_L2_3_G2_MINI_ALU_BoothXORCheck), .BoothResult ({
                  \$dummy [649],\$dummy [650],\$dummy [651],\$dummy [652],
                  \$dummy [653],\$dummy [654],\$dummy [655],\$dummy [656]}), .BoothAddingOperand (
                  {L1_3_L2_3_G2_MINI_ALU_BoothOperand_16,
                  L1_3_L2_3_G2_MINI_ALU_BoothOperand_15,
                  L1_3_L2_3_G2_MINI_ALU_BoothOperand_14,
                  L1_3_L2_3_G2_MINI_ALU_BoothOperand_13,
                  L1_3_L2_3_G2_MINI_ALU_BoothOperand_12,
                  L1_3_L2_3_G2_MINI_ALU_BoothOperand_11,
                  L1_3_L2_3_G2_MINI_ALU_BoothOperand_10,
                  L1_3_L2_3_G2_MINI_ALU_BoothOperand_9,\$dummy [657],
                  \$dummy [658],\$dummy [659],\$dummy [660],\$dummy [661],
                  \$dummy [662],\$dummy [663],\$dummy [664],\$dummy [665]}), .BoothP (
                  {L1_3_L2_3_G2_MINI_ALU_BoothP_16,
                  L1_3_L2_3_G2_MINI_ALU_BoothP_15,
                  L1_3_L2_3_G2_MINI_ALU_BoothP_14,
                  L1_3_L2_3_G2_MINI_ALU_BoothP_13,
                  L1_3_L2_3_G2_MINI_ALU_BoothP_12,
                  L1_3_L2_3_G2_MINI_ALU_BoothP_11,
                  L1_3_L2_3_G2_MINI_ALU_BoothP_10,L1_3_L2_3_G2_MINI_ALU_BoothP_9
                  ,L1_3_L2_3_G2_MINI_ALU_BoothP_8,L1_3_L2_3_G2_MINI_ALU_BoothP_7
                  ,L1_3_L2_3_G2_MINI_ALU_BoothP_6,L1_3_L2_3_G2_MINI_ALU_BoothP_5
                  ,L1_3_L2_3_G2_MINI_ALU_BoothP_4,L1_3_L2_3_G2_MINI_ALU_BoothP_3
                  ,L1_3_L2_3_G2_MINI_ALU_BoothP_2,L1_3_L2_3_G2_MINI_ALU_BoothP_1
                  ,L1_3_L2_3_G2_MINI_ALU_BoothP_0}), .LargeWindowShifted ({
                  \$dummy [666],\$dummy [667],\$dummy [668],\$dummy [669],
                  \$dummy [670],\$dummy [671],\$dummy [672],\$dummy [673],
                  \$dummy [674],\$dummy [675],\$dummy [676],\$dummy [677],
                  \$dummy [678],\$dummy [679],\$dummy [680],\$dummy [681],
                  \$dummy [682]})) ;
    booth_adder_17_unfolded13 L1_3_L2_4_G3_MINI_ALU_BOOTH_ADDER (.AdderFirstOperand (
                              {L2ResultsLarge_0__16,L2ResultsLarge_0__15,
                              L2ResultsLarge_0__14,L2ResultsLarge_0__13,
                              L2ResultsLarge_0__12,L2ResultsLarge_0__11,
                              L2ResultsLarge_0__10,L2ResultsLarge_0__9,
                              L2ResultsLarge_0__8,L2ResultsLarge_0__7,
                              L2ResultsLarge_0__6,L2ResultsLarge_0__5,
                              L2ResultsLarge_0__4,L2ResultsLarge_0__3,
                              L2ResultsLarge_0__2,L2ResultsLarge_0__1,
                              L2ResultsLarge_0__0}), .AdderSecondOperand ({
                              L2ResultsLarge_1__16,L2ResultsLarge_1__15,
                              L2ResultsLarge_1__14,L2ResultsLarge_1__13,
                              L2ResultsLarge_1__12,L2ResultsLarge_1__11,
                              L2ResultsLarge_1__10,L2ResultsLarge_1__9,
                              L2ResultsLarge_1__8,L2ResultsLarge_1__7,
                              L2ResultsLarge_1__6,L2ResultsLarge_1__5,
                              L2ResultsLarge_1__4,L2ResultsLarge_1__3,
                              L2ResultsLarge_1__2,L2ResultsLarge_1__1,
                              L2ResultsLarge_1__0}), .BoothOperand ({
                              L1_3_L2_4_G3_MINI_ALU_BoothOperand_16,
                              L1_3_L2_4_G3_MINI_ALU_BoothOperand_15,
                              L1_3_L2_4_G3_MINI_ALU_BoothOperand_14,
                              L1_3_L2_4_G3_MINI_ALU_BoothOperand_13,
                              L1_3_L2_4_G3_MINI_ALU_BoothOperand_12,
                              L1_3_L2_4_G3_MINI_ALU_BoothOperand_11,
                              L1_3_L2_4_G3_MINI_ALU_BoothOperand_10,
                              L1_3_L2_4_G3_MINI_ALU_BoothOperand_9,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16}), .BoothP ({
                              L1_3_L2_4_G3_MINI_ALU_BoothP_16,
                              L1_3_L2_4_G3_MINI_ALU_BoothP_15,
                              L1_3_L2_4_G3_MINI_ALU_BoothP_14,
                              L1_3_L2_4_G3_MINI_ALU_BoothP_13,
                              L1_3_L2_4_G3_MINI_ALU_BoothP_12,
                              L1_3_L2_4_G3_MINI_ALU_BoothP_11,
                              L1_3_L2_4_G3_MINI_ALU_BoothP_10,
                              L1_3_L2_4_G3_MINI_ALU_BoothP_9,
                              L1_3_L2_4_G3_MINI_ALU_BoothP_8,
                              L1_3_L2_4_G3_MINI_ALU_BoothP_7,
                              L1_3_L2_4_G3_MINI_ALU_BoothP_6,
                              L1_3_L2_4_G3_MINI_ALU_BoothP_5,
                              L1_3_L2_4_G3_MINI_ALU_BoothP_4,
                              L1_3_L2_4_G3_MINI_ALU_BoothP_3,
                              L1_3_L2_4_G3_MINI_ALU_BoothP_2,
                              L1_3_L2_4_G3_MINI_ALU_BoothP_1,
                              L1_3_L2_4_G3_MINI_ALU_BoothP_0}), .SelOperand (
                              nx3284), .Operation (
                              L1_3_L2_4_G3_MINI_ALU_BoothXORCheck), .AdderResult (
                              {L3ResultsLarge_0__16,L3ResultsLarge_0__15,
                              L3ResultsLarge_0__14,L3ResultsLarge_0__13,
                              L3ResultsLarge_0__12,L3ResultsLarge_0__11,
                              L3ResultsLarge_0__10,L3ResultsLarge_0__9,
                              L3ResultsLarge_0__8,L3ResultsLarge_0__7,
                              L3ResultsLarge_0__6,L3ResultsLarge_0__5,
                              L3ResultsLarge_0__4,L3ResultsLarge_0__3,
                              L3ResultsLarge_0__2,L3ResultsLarge_0__1,
                              L3ResultsLarge_0__0}), .AdderBoothResult ({
                              \$dummy [683],
                              L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_15,
                              L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_14,
                              L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_13,
                              L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_12,
                              L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_11,
                              L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_10,
                              L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_9,
                              L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_8,
                              L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_7,
                              L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_6,
                              L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_5,
                              L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_4,
                              L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_3,
                              L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_2,
                              L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_1,
                              L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_0})) ;
    booth_unit_17 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT (.CLK (CLK), .RST (RST), .Start (
                  Start), .Instr (Instr), .LoopingAndResultNotReady (nx3276), .Filter (
                  {FilterDin_3__4__7,FilterDin_3__4__6,FilterDin_3__4__5,
                  FilterDin_3__4__4,FilterDin_3__4__3,FilterDin_3__4__2,
                  FilterDin_3__4__1,FilterDin_3__4__0}), .Window ({
                  WindowDin_3__4__7,WindowDin_3__4__6,WindowDin_3__4__5,
                  WindowDin_3__4__4,WindowDin_3__4__3,WindowDin_3__4__2,
                  WindowDin_3__4__1,WindowDin_3__4__0}), .AdderBoothResult ({
                  L1FirstOperands_12__16,
                  L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_15,
                  L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_14,
                  L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_13,
                  L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_12,
                  L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_11,
                  L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_10,
                  L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_9,
                  L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_8,
                  L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_7,
                  L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_6,
                  L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_5,
                  L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_4,
                  L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_3,
                  L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_2,
                  L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_1,
                  L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_0}), .BoothXORCheck (
                  L1_3_L2_4_G3_MINI_ALU_BoothXORCheck), .BoothResult ({
                  \$dummy [684],\$dummy [685],\$dummy [686],\$dummy [687],
                  \$dummy [688],\$dummy [689],\$dummy [690],\$dummy [691]}), .BoothAddingOperand (
                  {L1_3_L2_4_G3_MINI_ALU_BoothOperand_16,
                  L1_3_L2_4_G3_MINI_ALU_BoothOperand_15,
                  L1_3_L2_4_G3_MINI_ALU_BoothOperand_14,
                  L1_3_L2_4_G3_MINI_ALU_BoothOperand_13,
                  L1_3_L2_4_G3_MINI_ALU_BoothOperand_12,
                  L1_3_L2_4_G3_MINI_ALU_BoothOperand_11,
                  L1_3_L2_4_G3_MINI_ALU_BoothOperand_10,
                  L1_3_L2_4_G3_MINI_ALU_BoothOperand_9,\$dummy [692],
                  \$dummy [693],\$dummy [694],\$dummy [695],\$dummy [696],
                  \$dummy [697],\$dummy [698],\$dummy [699],\$dummy [700]}), .BoothP (
                  {L1_3_L2_4_G3_MINI_ALU_BoothP_16,
                  L1_3_L2_4_G3_MINI_ALU_BoothP_15,
                  L1_3_L2_4_G3_MINI_ALU_BoothP_14,
                  L1_3_L2_4_G3_MINI_ALU_BoothP_13,
                  L1_3_L2_4_G3_MINI_ALU_BoothP_12,
                  L1_3_L2_4_G3_MINI_ALU_BoothP_11,
                  L1_3_L2_4_G3_MINI_ALU_BoothP_10,L1_3_L2_4_G3_MINI_ALU_BoothP_9
                  ,L1_3_L2_4_G3_MINI_ALU_BoothP_8,L1_3_L2_4_G3_MINI_ALU_BoothP_7
                  ,L1_3_L2_4_G3_MINI_ALU_BoothP_6,L1_3_L2_4_G3_MINI_ALU_BoothP_5
                  ,L1_3_L2_4_G3_MINI_ALU_BoothP_4,L1_3_L2_4_G3_MINI_ALU_BoothP_3
                  ,L1_3_L2_4_G3_MINI_ALU_BoothP_2,L1_3_L2_4_G3_MINI_ALU_BoothP_1
                  ,L1_3_L2_4_G3_MINI_ALU_BoothP_0}), .LargeWindowShifted ({
                  \$dummy [701],\$dummy [702],\$dummy [703],\$dummy [704],
                  \$dummy [705],\$dummy [706],\$dummy [707],\$dummy [708],
                  \$dummy [709],\$dummy [710],\$dummy [711],\$dummy [712],
                  \$dummy [713],\$dummy [714],\$dummy [715],\$dummy [716],
                  \$dummy [717]})) ;
    booth_adder_17_unfolded13 L1_4_L2_0_G3_MINI_ALU_BOOTH_ADDER (.AdderFirstOperand (
                              {L2ResultsLarge_2__16,L2ResultsLarge_2__15,
                              L2ResultsLarge_2__14,L2ResultsLarge_2__13,
                              L2ResultsLarge_2__12,L2ResultsLarge_2__11,
                              L2ResultsLarge_2__10,L2ResultsLarge_2__9,
                              L2ResultsLarge_2__8,L2ResultsLarge_2__7,
                              L2ResultsLarge_2__6,L2ResultsLarge_2__5,
                              L2ResultsLarge_2__4,L2ResultsLarge_2__3,
                              L2ResultsLarge_2__2,L2ResultsLarge_2__1,
                              L2ResultsLarge_2__0}), .AdderSecondOperand ({
                              L2ResultsLarge_3__16,L2ResultsLarge_3__15,
                              L2ResultsLarge_3__14,L2ResultsLarge_3__13,
                              L2ResultsLarge_3__12,L2ResultsLarge_3__11,
                              L2ResultsLarge_3__10,L2ResultsLarge_3__9,
                              L2ResultsLarge_3__8,L2ResultsLarge_3__7,
                              L2ResultsLarge_3__6,L2ResultsLarge_3__5,
                              L2ResultsLarge_3__4,L2ResultsLarge_3__3,
                              L2ResultsLarge_3__2,L2ResultsLarge_3__1,
                              L2ResultsLarge_3__0}), .BoothOperand ({
                              L1_4_L2_0_G3_MINI_ALU_BoothOperand_16,
                              L1_4_L2_0_G3_MINI_ALU_BoothOperand_15,
                              L1_4_L2_0_G3_MINI_ALU_BoothOperand_14,
                              L1_4_L2_0_G3_MINI_ALU_BoothOperand_13,
                              L1_4_L2_0_G3_MINI_ALU_BoothOperand_12,
                              L1_4_L2_0_G3_MINI_ALU_BoothOperand_11,
                              L1_4_L2_0_G3_MINI_ALU_BoothOperand_10,
                              L1_4_L2_0_G3_MINI_ALU_BoothOperand_9,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16}), .BoothP ({
                              L1_4_L2_0_G3_MINI_ALU_BoothP_16,
                              L1_4_L2_0_G3_MINI_ALU_BoothP_15,
                              L1_4_L2_0_G3_MINI_ALU_BoothP_14,
                              L1_4_L2_0_G3_MINI_ALU_BoothP_13,
                              L1_4_L2_0_G3_MINI_ALU_BoothP_12,
                              L1_4_L2_0_G3_MINI_ALU_BoothP_11,
                              L1_4_L2_0_G3_MINI_ALU_BoothP_10,
                              L1_4_L2_0_G3_MINI_ALU_BoothP_9,
                              L1_4_L2_0_G3_MINI_ALU_BoothP_8,
                              L1_4_L2_0_G3_MINI_ALU_BoothP_7,
                              L1_4_L2_0_G3_MINI_ALU_BoothP_6,
                              L1_4_L2_0_G3_MINI_ALU_BoothP_5,
                              L1_4_L2_0_G3_MINI_ALU_BoothP_4,
                              L1_4_L2_0_G3_MINI_ALU_BoothP_3,
                              L1_4_L2_0_G3_MINI_ALU_BoothP_2,
                              L1_4_L2_0_G3_MINI_ALU_BoothP_1,
                              L1_4_L2_0_G3_MINI_ALU_BoothP_0}), .SelOperand (
                              nx3284), .Operation (
                              L1_4_L2_0_G3_MINI_ALU_BoothXORCheck), .AdderResult (
                              {L3ResultsLarge_1__16,L3ResultsLarge_1__15,
                              L3ResultsLarge_1__14,L3ResultsLarge_1__13,
                              L3ResultsLarge_1__12,L3ResultsLarge_1__11,
                              L3ResultsLarge_1__10,L3ResultsLarge_1__9,
                              L3ResultsLarge_1__8,L3ResultsLarge_1__7,
                              L3ResultsLarge_1__6,L3ResultsLarge_1__5,
                              L3ResultsLarge_1__4,L3ResultsLarge_1__3,
                              L3ResultsLarge_1__2,L3ResultsLarge_1__1,
                              L3ResultsLarge_1__0}), .AdderBoothResult ({
                              \$dummy [718],
                              L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_15,
                              L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_14,
                              L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_13,
                              L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_12,
                              L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_11,
                              L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_10,
                              L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_9,
                              L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_8,
                              L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_7,
                              L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_6,
                              L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_5,
                              L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_4,
                              L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_3,
                              L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_2,
                              L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_1,
                              L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_0})) ;
    booth_unit_17 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT (.CLK (CLK), .RST (RST), .Start (
                  Start), .Instr (Instr), .LoopingAndResultNotReady (nx3276), .Filter (
                  {FilterDin_4__0__7,FilterDin_4__0__6,FilterDin_4__0__5,
                  FilterDin_4__0__4,FilterDin_4__0__3,FilterDin_4__0__2,
                  FilterDin_4__0__1,FilterDin_4__0__0}), .Window ({
                  WindowDin_4__0__7,WindowDin_4__0__6,WindowDin_4__0__5,
                  WindowDin_4__0__4,WindowDin_4__0__3,WindowDin_4__0__2,
                  WindowDin_4__0__1,WindowDin_4__0__0}), .AdderBoothResult ({
                  L1FirstOperands_12__16,
                  L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_15,
                  L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_14,
                  L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_13,
                  L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_12,
                  L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_11,
                  L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_10,
                  L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_9,
                  L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_8,
                  L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_7,
                  L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_6,
                  L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_5,
                  L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_4,
                  L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_3,
                  L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_2,
                  L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_1,
                  L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_0}), .BoothXORCheck (
                  L1_4_L2_0_G3_MINI_ALU_BoothXORCheck), .BoothResult ({
                  \$dummy [719],\$dummy [720],\$dummy [721],\$dummy [722],
                  \$dummy [723],\$dummy [724],\$dummy [725],\$dummy [726]}), .BoothAddingOperand (
                  {L1_4_L2_0_G3_MINI_ALU_BoothOperand_16,
                  L1_4_L2_0_G3_MINI_ALU_BoothOperand_15,
                  L1_4_L2_0_G3_MINI_ALU_BoothOperand_14,
                  L1_4_L2_0_G3_MINI_ALU_BoothOperand_13,
                  L1_4_L2_0_G3_MINI_ALU_BoothOperand_12,
                  L1_4_L2_0_G3_MINI_ALU_BoothOperand_11,
                  L1_4_L2_0_G3_MINI_ALU_BoothOperand_10,
                  L1_4_L2_0_G3_MINI_ALU_BoothOperand_9,\$dummy [727],
                  \$dummy [728],\$dummy [729],\$dummy [730],\$dummy [731],
                  \$dummy [732],\$dummy [733],\$dummy [734],\$dummy [735]}), .BoothP (
                  {L1_4_L2_0_G3_MINI_ALU_BoothP_16,
                  L1_4_L2_0_G3_MINI_ALU_BoothP_15,
                  L1_4_L2_0_G3_MINI_ALU_BoothP_14,
                  L1_4_L2_0_G3_MINI_ALU_BoothP_13,
                  L1_4_L2_0_G3_MINI_ALU_BoothP_12,
                  L1_4_L2_0_G3_MINI_ALU_BoothP_11,
                  L1_4_L2_0_G3_MINI_ALU_BoothP_10,L1_4_L2_0_G3_MINI_ALU_BoothP_9
                  ,L1_4_L2_0_G3_MINI_ALU_BoothP_8,L1_4_L2_0_G3_MINI_ALU_BoothP_7
                  ,L1_4_L2_0_G3_MINI_ALU_BoothP_6,L1_4_L2_0_G3_MINI_ALU_BoothP_5
                  ,L1_4_L2_0_G3_MINI_ALU_BoothP_4,L1_4_L2_0_G3_MINI_ALU_BoothP_3
                  ,L1_4_L2_0_G3_MINI_ALU_BoothP_2,L1_4_L2_0_G3_MINI_ALU_BoothP_1
                  ,L1_4_L2_0_G3_MINI_ALU_BoothP_0}), .LargeWindowShifted ({
                  \$dummy [736],\$dummy [737],\$dummy [738],\$dummy [739],
                  \$dummy [740],\$dummy [741],\$dummy [742],\$dummy [743],
                  \$dummy [744],\$dummy [745],\$dummy [746],\$dummy [747],
                  \$dummy [748],\$dummy [749],\$dummy [750],\$dummy [751],
                  \$dummy [752]})) ;
    booth_adder_17_unfolded13 L1_4_L2_1_G3_MINI_ALU_BOOTH_ADDER (.AdderFirstOperand (
                              {L2ResultsLarge_4__16,L2ResultsLarge_4__15,
                              L2ResultsLarge_4__14,L2ResultsLarge_4__13,
                              L2ResultsLarge_4__12,L2ResultsLarge_4__11,
                              L2ResultsLarge_4__10,L2ResultsLarge_4__9,
                              L2ResultsLarge_4__8,L2ResultsLarge_4__7,
                              L2ResultsLarge_4__6,L2ResultsLarge_4__5,
                              L2ResultsLarge_4__4,L2ResultsLarge_4__3,
                              L2ResultsLarge_4__2,L2ResultsLarge_4__1,
                              L2ResultsLarge_4__0}), .AdderSecondOperand ({
                              L2ResultsLarge_5__16,L2ResultsLarge_5__15,
                              L2ResultsLarge_5__14,L2ResultsLarge_5__13,
                              L2ResultsLarge_5__12,L2ResultsLarge_5__11,
                              L2ResultsLarge_5__10,L2ResultsLarge_5__9,
                              L2ResultsLarge_5__8,L2ResultsLarge_5__7,
                              L2ResultsLarge_5__6,L2ResultsLarge_5__5,
                              L2ResultsLarge_5__4,L2ResultsLarge_5__3,
                              L2ResultsLarge_5__2,L2ResultsLarge_5__1,
                              L2ResultsLarge_5__0}), .BoothOperand ({
                              L1_4_L2_1_G3_MINI_ALU_BoothOperand_16,
                              L1_4_L2_1_G3_MINI_ALU_BoothOperand_15,
                              L1_4_L2_1_G3_MINI_ALU_BoothOperand_14,
                              L1_4_L2_1_G3_MINI_ALU_BoothOperand_13,
                              L1_4_L2_1_G3_MINI_ALU_BoothOperand_12,
                              L1_4_L2_1_G3_MINI_ALU_BoothOperand_11,
                              L1_4_L2_1_G3_MINI_ALU_BoothOperand_10,
                              L1_4_L2_1_G3_MINI_ALU_BoothOperand_9,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16}), .BoothP ({
                              L1_4_L2_1_G3_MINI_ALU_BoothP_16,
                              L1_4_L2_1_G3_MINI_ALU_BoothP_15,
                              L1_4_L2_1_G3_MINI_ALU_BoothP_14,
                              L1_4_L2_1_G3_MINI_ALU_BoothP_13,
                              L1_4_L2_1_G3_MINI_ALU_BoothP_12,
                              L1_4_L2_1_G3_MINI_ALU_BoothP_11,
                              L1_4_L2_1_G3_MINI_ALU_BoothP_10,
                              L1_4_L2_1_G3_MINI_ALU_BoothP_9,
                              L1_4_L2_1_G3_MINI_ALU_BoothP_8,
                              L1_4_L2_1_G3_MINI_ALU_BoothP_7,
                              L1_4_L2_1_G3_MINI_ALU_BoothP_6,
                              L1_4_L2_1_G3_MINI_ALU_BoothP_5,
                              L1_4_L2_1_G3_MINI_ALU_BoothP_4,
                              L1_4_L2_1_G3_MINI_ALU_BoothP_3,
                              L1_4_L2_1_G3_MINI_ALU_BoothP_2,
                              L1_4_L2_1_G3_MINI_ALU_BoothP_1,
                              L1_4_L2_1_G3_MINI_ALU_BoothP_0}), .SelOperand (
                              nx3286), .Operation (
                              L1_4_L2_1_G3_MINI_ALU_BoothXORCheck), .AdderResult (
                              {L3ResultsLarge_2__16,L3ResultsLarge_2__15,
                              L3ResultsLarge_2__14,L3ResultsLarge_2__13,
                              L3ResultsLarge_2__12,L3ResultsLarge_2__11,
                              L3ResultsLarge_2__10,L3ResultsLarge_2__9,
                              L3ResultsLarge_2__8,L3ResultsLarge_2__7,
                              L3ResultsLarge_2__6,L3ResultsLarge_2__5,
                              L3ResultsLarge_2__4,L3ResultsLarge_2__3,
                              L3ResultsLarge_2__2,L3ResultsLarge_2__1,
                              L3ResultsLarge_2__0}), .AdderBoothResult ({
                              \$dummy [753],
                              L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_15,
                              L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_14,
                              L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_13,
                              L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_12,
                              L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_11,
                              L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_10,
                              L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_9,
                              L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_8,
                              L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_7,
                              L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_6,
                              L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_5,
                              L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_4,
                              L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_3,
                              L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_2,
                              L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_1,
                              L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_0})) ;
    booth_unit_17 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT (.CLK (CLK), .RST (RST), .Start (
                  Start), .Instr (Instr), .LoopingAndResultNotReady (nx3278), .Filter (
                  {FilterDin_4__1__7,FilterDin_4__1__6,FilterDin_4__1__5,
                  FilterDin_4__1__4,FilterDin_4__1__3,FilterDin_4__1__2,
                  FilterDin_4__1__1,FilterDin_4__1__0}), .Window ({
                  WindowDin_4__1__7,WindowDin_4__1__6,WindowDin_4__1__5,
                  WindowDin_4__1__4,WindowDin_4__1__3,WindowDin_4__1__2,
                  WindowDin_4__1__1,WindowDin_4__1__0}), .AdderBoothResult ({
                  L1FirstOperands_12__16,
                  L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_15,
                  L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_14,
                  L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_13,
                  L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_12,
                  L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_11,
                  L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_10,
                  L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_9,
                  L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_8,
                  L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_7,
                  L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_6,
                  L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_5,
                  L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_4,
                  L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_3,
                  L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_2,
                  L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_1,
                  L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_0}), .BoothXORCheck (
                  L1_4_L2_1_G3_MINI_ALU_BoothXORCheck), .BoothResult ({
                  \$dummy [754],\$dummy [755],\$dummy [756],\$dummy [757],
                  \$dummy [758],\$dummy [759],\$dummy [760],\$dummy [761]}), .BoothAddingOperand (
                  {L1_4_L2_1_G3_MINI_ALU_BoothOperand_16,
                  L1_4_L2_1_G3_MINI_ALU_BoothOperand_15,
                  L1_4_L2_1_G3_MINI_ALU_BoothOperand_14,
                  L1_4_L2_1_G3_MINI_ALU_BoothOperand_13,
                  L1_4_L2_1_G3_MINI_ALU_BoothOperand_12,
                  L1_4_L2_1_G3_MINI_ALU_BoothOperand_11,
                  L1_4_L2_1_G3_MINI_ALU_BoothOperand_10,
                  L1_4_L2_1_G3_MINI_ALU_BoothOperand_9,\$dummy [762],
                  \$dummy [763],\$dummy [764],\$dummy [765],\$dummy [766],
                  \$dummy [767],\$dummy [768],\$dummy [769],\$dummy [770]}), .BoothP (
                  {L1_4_L2_1_G3_MINI_ALU_BoothP_16,
                  L1_4_L2_1_G3_MINI_ALU_BoothP_15,
                  L1_4_L2_1_G3_MINI_ALU_BoothP_14,
                  L1_4_L2_1_G3_MINI_ALU_BoothP_13,
                  L1_4_L2_1_G3_MINI_ALU_BoothP_12,
                  L1_4_L2_1_G3_MINI_ALU_BoothP_11,
                  L1_4_L2_1_G3_MINI_ALU_BoothP_10,L1_4_L2_1_G3_MINI_ALU_BoothP_9
                  ,L1_4_L2_1_G3_MINI_ALU_BoothP_8,L1_4_L2_1_G3_MINI_ALU_BoothP_7
                  ,L1_4_L2_1_G3_MINI_ALU_BoothP_6,L1_4_L2_1_G3_MINI_ALU_BoothP_5
                  ,L1_4_L2_1_G3_MINI_ALU_BoothP_4,L1_4_L2_1_G3_MINI_ALU_BoothP_3
                  ,L1_4_L2_1_G3_MINI_ALU_BoothP_2,L1_4_L2_1_G3_MINI_ALU_BoothP_1
                  ,L1_4_L2_1_G3_MINI_ALU_BoothP_0}), .LargeWindowShifted ({
                  \$dummy [771],\$dummy [772],\$dummy [773],\$dummy [774],
                  \$dummy [775],\$dummy [776],\$dummy [777],\$dummy [778],
                  \$dummy [779],\$dummy [780],\$dummy [781],\$dummy [782],
                  \$dummy [783],\$dummy [784],\$dummy [785],\$dummy [786],
                  \$dummy [787]})) ;
    booth_adder_17_unfolded13 L1_4_L2_2_G4_MINI_ALU_BOOTH_ADDER (.AdderFirstOperand (
                              {L3ResultsLarge_0__16,L3ResultsLarge_0__15,
                              L3ResultsLarge_0__14,L3ResultsLarge_0__13,
                              L3ResultsLarge_0__12,L3ResultsLarge_0__11,
                              L3ResultsLarge_0__10,L3ResultsLarge_0__9,
                              L3ResultsLarge_0__8,L3ResultsLarge_0__7,
                              L3ResultsLarge_0__6,L3ResultsLarge_0__5,
                              L3ResultsLarge_0__4,L3ResultsLarge_0__3,
                              L3ResultsLarge_0__2,L3ResultsLarge_0__1,
                              L3ResultsLarge_0__0}), .AdderSecondOperand ({
                              L3ResultsLarge_1__16,L3ResultsLarge_1__15,
                              L3ResultsLarge_1__14,L3ResultsLarge_1__13,
                              L3ResultsLarge_1__12,L3ResultsLarge_1__11,
                              L3ResultsLarge_1__10,L3ResultsLarge_1__9,
                              L3ResultsLarge_1__8,L3ResultsLarge_1__7,
                              L3ResultsLarge_1__6,L3ResultsLarge_1__5,
                              L3ResultsLarge_1__4,L3ResultsLarge_1__3,
                              L3ResultsLarge_1__2,L3ResultsLarge_1__1,
                              L3ResultsLarge_1__0}), .BoothOperand ({
                              L1_4_L2_2_G4_MINI_ALU_BoothOperand_16,
                              L1_4_L2_2_G4_MINI_ALU_BoothOperand_15,
                              L1_4_L2_2_G4_MINI_ALU_BoothOperand_14,
                              L1_4_L2_2_G4_MINI_ALU_BoothOperand_13,
                              L1_4_L2_2_G4_MINI_ALU_BoothOperand_12,
                              L1_4_L2_2_G4_MINI_ALU_BoothOperand_11,
                              L1_4_L2_2_G4_MINI_ALU_BoothOperand_10,
                              L1_4_L2_2_G4_MINI_ALU_BoothOperand_9,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16}), .BoothP ({
                              L1_4_L2_2_G4_MINI_ALU_BoothP_16,
                              L1_4_L2_2_G4_MINI_ALU_BoothP_15,
                              L1_4_L2_2_G4_MINI_ALU_BoothP_14,
                              L1_4_L2_2_G4_MINI_ALU_BoothP_13,
                              L1_4_L2_2_G4_MINI_ALU_BoothP_12,
                              L1_4_L2_2_G4_MINI_ALU_BoothP_11,
                              L1_4_L2_2_G4_MINI_ALU_BoothP_10,
                              L1_4_L2_2_G4_MINI_ALU_BoothP_9,
                              L1_4_L2_2_G4_MINI_ALU_BoothP_8,
                              L1_4_L2_2_G4_MINI_ALU_BoothP_7,
                              L1_4_L2_2_G4_MINI_ALU_BoothP_6,
                              L1_4_L2_2_G4_MINI_ALU_BoothP_5,
                              L1_4_L2_2_G4_MINI_ALU_BoothP_4,
                              L1_4_L2_2_G4_MINI_ALU_BoothP_3,
                              L1_4_L2_2_G4_MINI_ALU_BoothP_2,
                              L1_4_L2_2_G4_MINI_ALU_BoothP_1,
                              L1_4_L2_2_G4_MINI_ALU_BoothP_0}), .SelOperand (
                              nx3286), .Operation (
                              L1_4_L2_2_G4_MINI_ALU_BoothXORCheck), .AdderResult (
                              {L4ResultsLarge_0__16,L4ResultsLarge_0__15,
                              L4ResultsLarge_0__14,L4ResultsLarge_0__13,
                              L4ResultsLarge_0__12,L4ResultsLarge_0__11,
                              L4ResultsLarge_0__10,L4ResultsLarge_0__9,
                              L4ResultsLarge_0__8,L4ResultsLarge_0__7,
                              L4ResultsLarge_0__6,L4ResultsLarge_0__5,
                              L4ResultsLarge_0__4,L4ResultsLarge_0__3,
                              L4ResultsLarge_0__2,L4ResultsLarge_0__1,
                              L4ResultsLarge_0__0}), .AdderBoothResult ({
                              \$dummy [788],
                              L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_15,
                              L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_14,
                              L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_13,
                              L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_12,
                              L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_11,
                              L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_10,
                              L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_9,
                              L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_8,
                              L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_7,
                              L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_6,
                              L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_5,
                              L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_4,
                              L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_3,
                              L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_2,
                              L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_1,
                              L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_0})) ;
    booth_unit_17 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT (.CLK (CLK), .RST (RST), .Start (
                  Start), .Instr (Instr), .LoopingAndResultNotReady (nx3278), .Filter (
                  {FilterDin_4__2__7,FilterDin_4__2__6,FilterDin_4__2__5,
                  FilterDin_4__2__4,FilterDin_4__2__3,FilterDin_4__2__2,
                  FilterDin_4__2__1,FilterDin_4__2__0}), .Window ({
                  WindowDin_4__2__7,WindowDin_4__2__6,WindowDin_4__2__5,
                  WindowDin_4__2__4,WindowDin_4__2__3,WindowDin_4__2__2,
                  WindowDin_4__2__1,WindowDin_4__2__0}), .AdderBoothResult ({
                  L1FirstOperands_12__16,
                  L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_15,
                  L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_14,
                  L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_13,
                  L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_12,
                  L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_11,
                  L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_10,
                  L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_9,
                  L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_8,
                  L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_7,
                  L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_6,
                  L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_5,
                  L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_4,
                  L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_3,
                  L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_2,
                  L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_1,
                  L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_0}), .BoothXORCheck (
                  L1_4_L2_2_G4_MINI_ALU_BoothXORCheck), .BoothResult ({
                  \$dummy [789],\$dummy [790],\$dummy [791],\$dummy [792],
                  \$dummy [793],\$dummy [794],\$dummy [795],\$dummy [796]}), .BoothAddingOperand (
                  {L1_4_L2_2_G4_MINI_ALU_BoothOperand_16,
                  L1_4_L2_2_G4_MINI_ALU_BoothOperand_15,
                  L1_4_L2_2_G4_MINI_ALU_BoothOperand_14,
                  L1_4_L2_2_G4_MINI_ALU_BoothOperand_13,
                  L1_4_L2_2_G4_MINI_ALU_BoothOperand_12,
                  L1_4_L2_2_G4_MINI_ALU_BoothOperand_11,
                  L1_4_L2_2_G4_MINI_ALU_BoothOperand_10,
                  L1_4_L2_2_G4_MINI_ALU_BoothOperand_9,\$dummy [797],
                  \$dummy [798],\$dummy [799],\$dummy [800],\$dummy [801],
                  \$dummy [802],\$dummy [803],\$dummy [804],\$dummy [805]}), .BoothP (
                  {L1_4_L2_2_G4_MINI_ALU_BoothP_16,
                  L1_4_L2_2_G4_MINI_ALU_BoothP_15,
                  L1_4_L2_2_G4_MINI_ALU_BoothP_14,
                  L1_4_L2_2_G4_MINI_ALU_BoothP_13,
                  L1_4_L2_2_G4_MINI_ALU_BoothP_12,
                  L1_4_L2_2_G4_MINI_ALU_BoothP_11,
                  L1_4_L2_2_G4_MINI_ALU_BoothP_10,L1_4_L2_2_G4_MINI_ALU_BoothP_9
                  ,L1_4_L2_2_G4_MINI_ALU_BoothP_8,L1_4_L2_2_G4_MINI_ALU_BoothP_7
                  ,L1_4_L2_2_G4_MINI_ALU_BoothP_6,L1_4_L2_2_G4_MINI_ALU_BoothP_5
                  ,L1_4_L2_2_G4_MINI_ALU_BoothP_4,L1_4_L2_2_G4_MINI_ALU_BoothP_3
                  ,L1_4_L2_2_G4_MINI_ALU_BoothP_2,L1_4_L2_2_G4_MINI_ALU_BoothP_1
                  ,L1_4_L2_2_G4_MINI_ALU_BoothP_0}), .LargeWindowShifted ({
                  \$dummy [806],\$dummy [807],\$dummy [808],\$dummy [809],
                  \$dummy [810],\$dummy [811],\$dummy [812],\$dummy [813],
                  \$dummy [814],\$dummy [815],\$dummy [816],\$dummy [817],
                  \$dummy [818],\$dummy [819],\$dummy [820],\$dummy [821],
                  \$dummy [822]})) ;
    booth_adder_17_unfolded13 L1_4_L2_3_G5_MINI_ALU_BOOTH_ADDER (.AdderFirstOperand (
                              {L4ResultsLarge_0__16,L4ResultsLarge_0__15,
                              L4ResultsLarge_0__14,L4ResultsLarge_0__13,
                              L4ResultsLarge_0__12,L4ResultsLarge_0__11,
                              L4ResultsLarge_0__10,L4ResultsLarge_0__9,
                              L4ResultsLarge_0__8,L4ResultsLarge_0__7,
                              L4ResultsLarge_0__6,L4ResultsLarge_0__5,
                              L4ResultsLarge_0__4,L4ResultsLarge_0__3,
                              L4ResultsLarge_0__2,L4ResultsLarge_0__1,
                              L4ResultsLarge_0__0}), .AdderSecondOperand ({
                              L3ResultsLarge_2__16,L3ResultsLarge_2__15,
                              L3ResultsLarge_2__14,L3ResultsLarge_2__13,
                              L3ResultsLarge_2__12,L3ResultsLarge_2__11,
                              L3ResultsLarge_2__10,L3ResultsLarge_2__9,
                              L3ResultsLarge_2__8,L3ResultsLarge_2__7,
                              L3ResultsLarge_2__6,L3ResultsLarge_2__5,
                              L3ResultsLarge_2__4,L3ResultsLarge_2__3,
                              L3ResultsLarge_2__2,L3ResultsLarge_2__1,
                              L3ResultsLarge_2__0}), .BoothOperand ({
                              L1_4_L2_3_G5_MINI_ALU_BoothOperand_16,
                              L1_4_L2_3_G5_MINI_ALU_BoothOperand_15,
                              L1_4_L2_3_G5_MINI_ALU_BoothOperand_14,
                              L1_4_L2_3_G5_MINI_ALU_BoothOperand_13,
                              L1_4_L2_3_G5_MINI_ALU_BoothOperand_12,
                              L1_4_L2_3_G5_MINI_ALU_BoothOperand_11,
                              L1_4_L2_3_G5_MINI_ALU_BoothOperand_10,
                              L1_4_L2_3_G5_MINI_ALU_BoothOperand_9,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16}), .BoothP ({
                              L1_4_L2_3_G5_MINI_ALU_BoothP_16,
                              L1_4_L2_3_G5_MINI_ALU_BoothP_15,
                              L1_4_L2_3_G5_MINI_ALU_BoothP_14,
                              L1_4_L2_3_G5_MINI_ALU_BoothP_13,
                              L1_4_L2_3_G5_MINI_ALU_BoothP_12,
                              L1_4_L2_3_G5_MINI_ALU_BoothP_11,
                              L1_4_L2_3_G5_MINI_ALU_BoothP_10,
                              L1_4_L2_3_G5_MINI_ALU_BoothP_9,
                              L1_4_L2_3_G5_MINI_ALU_BoothP_8,
                              L1_4_L2_3_G5_MINI_ALU_BoothP_7,
                              L1_4_L2_3_G5_MINI_ALU_BoothP_6,
                              L1_4_L2_3_G5_MINI_ALU_BoothP_5,
                              L1_4_L2_3_G5_MINI_ALU_BoothP_4,
                              L1_4_L2_3_G5_MINI_ALU_BoothP_3,
                              L1_4_L2_3_G5_MINI_ALU_BoothP_2,
                              L1_4_L2_3_G5_MINI_ALU_BoothP_1,
                              L1_4_L2_3_G5_MINI_ALU_BoothP_0}), .SelOperand (
                              nx3286), .Operation (
                              L1_4_L2_3_G5_MINI_ALU_BoothXORCheck), .AdderResult (
                              {L5FirstOperands_1__16,L5FirstOperands_1__15,
                              L5FirstOperands_1__14,L5FirstOperands_1__13,
                              L5FirstOperands_1__12,L5FirstOperands_1__11,
                              L5FirstOperands_1__10,L5FirstOperands_1__9,
                              L5FirstOperands_1__8,L5FirstOperands_1__7,
                              L5FirstOperands_1__6,L5FirstOperands_1__5,
                              L5FirstOperands_1__4,L5FirstOperands_1__3,
                              L5FirstOperands_1__2,L5FirstOperands_1__1,
                              L5FirstOperands_1__0}), .AdderBoothResult ({
                              \$dummy [823],
                              L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_15,
                              L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_14,
                              L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_13,
                              L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_12,
                              L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_11,
                              L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_10,
                              L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_9,
                              L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_8,
                              L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_7,
                              L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_6,
                              L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_5,
                              L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_4,
                              L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_3,
                              L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_2,
                              L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_1,
                              L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_0})) ;
    booth_unit_17 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT (.CLK (CLK), .RST (RST), .Start (
                  Start), .Instr (Instr), .LoopingAndResultNotReady (nx3278), .Filter (
                  {FilterDin_4__3__7,FilterDin_4__3__6,FilterDin_4__3__5,
                  FilterDin_4__3__4,FilterDin_4__3__3,FilterDin_4__3__2,
                  FilterDin_4__3__1,FilterDin_4__3__0}), .Window ({
                  WindowDin_4__3__7,WindowDin_4__3__6,WindowDin_4__3__5,
                  WindowDin_4__3__4,WindowDin_4__3__3,WindowDin_4__3__2,
                  WindowDin_4__3__1,WindowDin_4__3__0}), .AdderBoothResult ({
                  L1FirstOperands_12__16,
                  L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_15,
                  L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_14,
                  L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_13,
                  L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_12,
                  L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_11,
                  L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_10,
                  L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_9,
                  L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_8,
                  L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_7,
                  L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_6,
                  L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_5,
                  L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_4,
                  L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_3,
                  L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_2,
                  L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_1,
                  L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_0}), .BoothXORCheck (
                  L1_4_L2_3_G5_MINI_ALU_BoothXORCheck), .BoothResult ({
                  \$dummy [824],\$dummy [825],\$dummy [826],\$dummy [827],
                  \$dummy [828],\$dummy [829],\$dummy [830],\$dummy [831]}), .BoothAddingOperand (
                  {L1_4_L2_3_G5_MINI_ALU_BoothOperand_16,
                  L1_4_L2_3_G5_MINI_ALU_BoothOperand_15,
                  L1_4_L2_3_G5_MINI_ALU_BoothOperand_14,
                  L1_4_L2_3_G5_MINI_ALU_BoothOperand_13,
                  L1_4_L2_3_G5_MINI_ALU_BoothOperand_12,
                  L1_4_L2_3_G5_MINI_ALU_BoothOperand_11,
                  L1_4_L2_3_G5_MINI_ALU_BoothOperand_10,
                  L1_4_L2_3_G5_MINI_ALU_BoothOperand_9,\$dummy [832],
                  \$dummy [833],\$dummy [834],\$dummy [835],\$dummy [836],
                  \$dummy [837],\$dummy [838],\$dummy [839],\$dummy [840]}), .BoothP (
                  {L1_4_L2_3_G5_MINI_ALU_BoothP_16,
                  L1_4_L2_3_G5_MINI_ALU_BoothP_15,
                  L1_4_L2_3_G5_MINI_ALU_BoothP_14,
                  L1_4_L2_3_G5_MINI_ALU_BoothP_13,
                  L1_4_L2_3_G5_MINI_ALU_BoothP_12,
                  L1_4_L2_3_G5_MINI_ALU_BoothP_11,
                  L1_4_L2_3_G5_MINI_ALU_BoothP_10,L1_4_L2_3_G5_MINI_ALU_BoothP_9
                  ,L1_4_L2_3_G5_MINI_ALU_BoothP_8,L1_4_L2_3_G5_MINI_ALU_BoothP_7
                  ,L1_4_L2_3_G5_MINI_ALU_BoothP_6,L1_4_L2_3_G5_MINI_ALU_BoothP_5
                  ,L1_4_L2_3_G5_MINI_ALU_BoothP_4,L1_4_L2_3_G5_MINI_ALU_BoothP_3
                  ,L1_4_L2_3_G5_MINI_ALU_BoothP_2,L1_4_L2_3_G5_MINI_ALU_BoothP_1
                  ,L1_4_L2_3_G5_MINI_ALU_BoothP_0}), .LargeWindowShifted ({
                  \$dummy [841],\$dummy [842],\$dummy [843],\$dummy [844],
                  \$dummy [845],\$dummy [846],\$dummy [847],\$dummy [848],
                  \$dummy [849],\$dummy [850],\$dummy [851],\$dummy [852],
                  \$dummy [853],\$dummy [854],\$dummy [855],\$dummy [856],
                  \$dummy [857]})) ;
    booth_adder_17_unfolded14 L1_4_L2_4_G5_MINI_ALU_BOOTH_ADDER (.AdderFirstOperand (
                              {L5FirstOperands_1__16,L5FirstOperands_1__15,
                              L5FirstOperands_1__14,L5FirstOperands_1__13,
                              L5FirstOperands_1__12,L5FirstOperands_1__11,
                              L5FirstOperands_1__10,L5FirstOperands_1__9,
                              L5FirstOperands_1__8,L5FirstOperands_1__7,
                              L5FirstOperands_1__6,L5FirstOperands_1__5,
                              L5FirstOperands_1__4,L5FirstOperands_1__3,
                              L5FirstOperands_1__2,L5FirstOperands_1__1,
                              L5FirstOperands_1__0}), .AdderSecondOperand ({
                              L1FirstOperands_12__16,
                              L1_4_L2_4_G5_MINI_ALU_OperationResult_15,
                              L1_4_L2_4_G5_MINI_ALU_OperationResult_14,
                              L1_4_L2_4_G5_MINI_ALU_OperationResult_13,
                              L1_4_L2_4_G5_MINI_ALU_OperationResult_12,
                              L1_4_L2_4_G5_MINI_ALU_OperationResult_11,
                              L1_4_L2_4_G5_MINI_ALU_OperationResult_10,
                              L1_4_L2_4_G5_MINI_ALU_OperationResult_9,
                              L1_4_L2_4_G5_MINI_ALU_OperationResult_8,
                              L1_4_L2_4_G5_MINI_ALU_OperationResult_7,
                              L1_4_L2_4_G5_MINI_ALU_OperationResult_6,
                              L1_4_L2_4_G5_MINI_ALU_OperationResult_5,
                              L1_4_L2_4_G5_MINI_ALU_OperationResult_4,
                              L1_4_L2_4_G5_MINI_ALU_OperationResult_3,
                              L1_4_L2_4_G5_MINI_ALU_OperationResult_2,
                              L1_4_L2_4_G5_MINI_ALU_OperationResult_1,
                              L1_4_L2_4_G5_MINI_ALU_OperationResult_0}), .BoothOperand (
                              {L1_4_L2_4_G5_MINI_ALU_BoothOperand_16,
                              L1_4_L2_4_G5_MINI_ALU_BoothOperand_15,
                              L1_4_L2_4_G5_MINI_ALU_BoothOperand_14,
                              L1_4_L2_4_G5_MINI_ALU_BoothOperand_13,
                              L1_4_L2_4_G5_MINI_ALU_BoothOperand_12,
                              L1_4_L2_4_G5_MINI_ALU_BoothOperand_11,
                              L1_4_L2_4_G5_MINI_ALU_BoothOperand_10,
                              L1_4_L2_4_G5_MINI_ALU_BoothOperand_9,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16}), .BoothP ({
                              L1_4_L2_4_G5_MINI_ALU_BoothP_16,
                              L1_4_L2_4_G5_MINI_ALU_BoothP_15,
                              L1_4_L2_4_G5_MINI_ALU_BoothP_14,
                              L1_4_L2_4_G5_MINI_ALU_BoothP_13,
                              L1_4_L2_4_G5_MINI_ALU_BoothP_12,
                              L1_4_L2_4_G5_MINI_ALU_BoothP_11,
                              L1_4_L2_4_G5_MINI_ALU_BoothP_10,
                              L1_4_L2_4_G5_MINI_ALU_BoothP_9,
                              L1_4_L2_4_G5_MINI_ALU_BoothP_8,
                              L1_4_L2_4_G5_MINI_ALU_BoothP_7,
                              L1_4_L2_4_G5_MINI_ALU_BoothP_6,
                              L1_4_L2_4_G5_MINI_ALU_BoothP_5,
                              L1_4_L2_4_G5_MINI_ALU_BoothP_4,
                              L1_4_L2_4_G5_MINI_ALU_BoothP_3,
                              L1_4_L2_4_G5_MINI_ALU_BoothP_2,
                              L1_4_L2_4_G5_MINI_ALU_BoothP_1,
                              L1_4_L2_4_G5_MINI_ALU_BoothP_0}), .SelOperand (
                              nx3286), .Operation (
                              L1_4_L2_4_G5_MINI_ALU_BoothXORCheck), .AdderResult (
                              {\$dummy [858],\$dummy [859],\$dummy [860],
                              \$dummy [861],\$dummy [862],\$dummy [863],
                              \$dummy [864],\$dummy [865],\$dummy [866],
                              L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_7,
                              L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_6,
                              L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_5,
                              L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_4,
                              L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_3,
                              L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_2,
                              L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_1,
                              L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_0}), .AdderBoothResult (
                              {\$dummy [867],
                              L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_15,
                              L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_14,
                              L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_13,
                              L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_12,
                              L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_11,
                              L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_10,
                              L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_9,
                              L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_8,
                              L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_7,
                              L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_6,
                              L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_5,
                              L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_4,
                              L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_3,
                              L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_2,
                              L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_1,
                              L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_0})) ;
    booth_unit_17 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT (.CLK (CLK), .RST (RST), .Start (
                  Start), .Instr (Instr), .LoopingAndResultNotReady (nx3278), .Filter (
                  {FilterDin_4__4__7,FilterDin_4__4__6,FilterDin_4__4__5,
                  FilterDin_4__4__4,FilterDin_4__4__3,FilterDin_4__4__2,
                  FilterDin_4__4__1,FilterDin_4__4__0}), .Window ({
                  WindowDin_4__4__7,WindowDin_4__4__6,WindowDin_4__4__5,
                  WindowDin_4__4__4,WindowDin_4__4__3,WindowDin_4__4__2,
                  WindowDin_4__4__1,WindowDin_4__4__0}), .AdderBoothResult ({
                  L1FirstOperands_12__16,
                  L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_15,
                  L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_14,
                  L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_13,
                  L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_12,
                  L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_11,
                  L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_10,
                  L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_9,
                  L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_8,
                  L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_7,
                  L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_6,
                  L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_5,
                  L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_4,
                  L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_3,
                  L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_2,
                  L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_1,
                  L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_0}), .BoothXORCheck (
                  L1_4_L2_4_G5_MINI_ALU_BoothXORCheck), .BoothResult ({
                  \$dummy [868],\$dummy [869],\$dummy [870],\$dummy [871],
                  \$dummy [872],\$dummy [873],\$dummy [874],\$dummy [875]}), .BoothAddingOperand (
                  {L1_4_L2_4_G5_MINI_ALU_BoothOperand_16,
                  L1_4_L2_4_G5_MINI_ALU_BoothOperand_15,
                  L1_4_L2_4_G5_MINI_ALU_BoothOperand_14,
                  L1_4_L2_4_G5_MINI_ALU_BoothOperand_13,
                  L1_4_L2_4_G5_MINI_ALU_BoothOperand_12,
                  L1_4_L2_4_G5_MINI_ALU_BoothOperand_11,
                  L1_4_L2_4_G5_MINI_ALU_BoothOperand_10,
                  L1_4_L2_4_G5_MINI_ALU_BoothOperand_9,\$dummy [876],
                  \$dummy [877],\$dummy [878],\$dummy [879],\$dummy [880],
                  \$dummy [881],\$dummy [882],\$dummy [883],\$dummy [884]}), .BoothP (
                  {L1_4_L2_4_G5_MINI_ALU_BoothP_16,
                  L1_4_L2_4_G5_MINI_ALU_BoothP_15,
                  L1_4_L2_4_G5_MINI_ALU_BoothP_14,
                  L1_4_L2_4_G5_MINI_ALU_BoothP_13,
                  L1_4_L2_4_G5_MINI_ALU_BoothP_12,
                  L1_4_L2_4_G5_MINI_ALU_BoothP_11,
                  L1_4_L2_4_G5_MINI_ALU_BoothP_10,L1_4_L2_4_G5_MINI_ALU_BoothP_9
                  ,L1_4_L2_4_G5_MINI_ALU_BoothP_8,L1_4_L2_4_G5_MINI_ALU_BoothP_7
                  ,L1_4_L2_4_G5_MINI_ALU_BoothP_6,L1_4_L2_4_G5_MINI_ALU_BoothP_5
                  ,L1_4_L2_4_G5_MINI_ALU_BoothP_4,L1_4_L2_4_G5_MINI_ALU_BoothP_3
                  ,L1_4_L2_4_G5_MINI_ALU_BoothP_2,L1_4_L2_4_G5_MINI_ALU_BoothP_1
                  ,L1_4_L2_4_G5_MINI_ALU_BoothP_0}), .LargeWindowShifted ({
                  \$dummy [885],\$dummy [886],\$dummy [887],\$dummy [888],
                  \$dummy [889],\$dummy [890],\$dummy [891],\$dummy [892],
                  \$dummy [893],\$dummy [894],\$dummy [895],\$dummy [896],
                  \$dummy [897],\$dummy [898],\$dummy [899],\$dummy [900],
                  \$dummy [901]})) ;
    nor02ii ix2852 (.Y (NOT__145383), .A0 (Instr), .A1 (nx2853)) ;
    nand03 ix2854 (.Y (nx2853), .A0 (CounterOut_0), .A1 (CounterOut_3), .A2 (
           nx2873)) ;
    dffr reg_CounterOut_0 (.Q (CounterOut_0), .QB (NOT_CounterOut_0), .D (
         NOT_CounterOut_0), .CLK (nx1032), .R (nx1036)) ;
    or02 ix1037 (.Y (nx1036), .A0 (Start), .A1 (RST)) ;
    dffr reg_CounterOut_3 (.Q (CounterOut_3), .QB (\$dummy [902]), .D (nx1066), 
         .CLK (nx1032), .R (nx1036)) ;
    xnor2 ix1067 (.Y (nx1066), .A0 (CounterOut_3), .A1 (nx2865)) ;
    nand03 ix2866 (.Y (nx2865), .A0 (CounterOut_2), .A1 (CounterOut_1), .A2 (
           CounterOut_0)) ;
    dffr reg_CounterOut_2 (.Q (CounterOut_2), .QB (\$dummy [903]), .D (nx1058), 
         .CLK (nx1032), .R (nx1036)) ;
    xnor2 ix1059 (.Y (nx1058), .A0 (CounterOut_2), .A1 (nx2869)) ;
    dffr reg_CounterOut_1 (.Q (CounterOut_1), .QB (nx2873), .D (nx1046), .CLK (
         nx1032), .R (nx1036)) ;
    fake_gnd ix2302 (.Y (L1FirstOperands_12__16)) ;
    mux21_ni ix109 (.Y (L1_4_L2_4_G5_MINI_ALU_OperationResult_0), .A0 (
             L1_4_L2_4_G5_MINI_ALU_BoothP_1), .A1 (WindowDin_4__4__0), .S0 (
             Instr)) ;
    mux21_ni ix117 (.Y (L1_4_L2_4_G5_MINI_ALU_OperationResult_1), .A0 (
             L1_4_L2_4_G5_MINI_ALU_BoothP_2), .A1 (WindowDin_4__4__1), .S0 (
             Instr)) ;
    mux21_ni ix125 (.Y (L1_4_L2_4_G5_MINI_ALU_OperationResult_2), .A0 (
             L1_4_L2_4_G5_MINI_ALU_BoothP_3), .A1 (WindowDin_4__4__2), .S0 (
             Instr)) ;
    mux21_ni ix133 (.Y (L1_4_L2_4_G5_MINI_ALU_OperationResult_3), .A0 (
             L1_4_L2_4_G5_MINI_ALU_BoothP_4), .A1 (WindowDin_4__4__3), .S0 (
             Instr)) ;
    mux21_ni ix141 (.Y (L1_4_L2_4_G5_MINI_ALU_OperationResult_4), .A0 (
             L1_4_L2_4_G5_MINI_ALU_BoothP_5), .A1 (WindowDin_4__4__4), .S0 (
             Instr)) ;
    mux21_ni ix149 (.Y (L1_4_L2_4_G5_MINI_ALU_OperationResult_5), .A0 (
             L1_4_L2_4_G5_MINI_ALU_BoothP_6), .A1 (WindowDin_4__4__5), .S0 (
             Instr)) ;
    mux21_ni ix157 (.Y (L1_4_L2_4_G5_MINI_ALU_OperationResult_6), .A0 (
             L1_4_L2_4_G5_MINI_ALU_BoothP_7), .A1 (WindowDin_4__4__6), .S0 (
             Instr)) ;
    mux21_ni ix165 (.Y (L1_4_L2_4_G5_MINI_ALU_OperationResult_7), .A0 (
             L1_4_L2_4_G5_MINI_ALU_BoothP_8), .A1 (WindowDin_4__4__7), .S0 (
             Instr)) ;
    nor02ii ix73 (.Y (L1_4_L2_4_G5_MINI_ALU_OperationResult_8), .A0 (Instr), .A1 (
            L1_4_L2_4_G5_MINI_ALU_BoothP_9)) ;
    nor02ii ix77 (.Y (L1_4_L2_4_G5_MINI_ALU_OperationResult_9), .A0 (Instr), .A1 (
            L1_4_L2_4_G5_MINI_ALU_BoothP_10)) ;
    nor02ii ix81 (.Y (L1_4_L2_4_G5_MINI_ALU_OperationResult_10), .A0 (Instr), .A1 (
            L1_4_L2_4_G5_MINI_ALU_BoothP_11)) ;
    nor02ii ix85 (.Y (L1_4_L2_4_G5_MINI_ALU_OperationResult_11), .A0 (Instr), .A1 (
            L1_4_L2_4_G5_MINI_ALU_BoothP_12)) ;
    nor02ii ix89 (.Y (L1_4_L2_4_G5_MINI_ALU_OperationResult_12), .A0 (Instr), .A1 (
            L1_4_L2_4_G5_MINI_ALU_BoothP_13)) ;
    nor02ii ix93 (.Y (L1_4_L2_4_G5_MINI_ALU_OperationResult_13), .A0 (Instr), .A1 (
            L1_4_L2_4_G5_MINI_ALU_BoothP_14)) ;
    nor02ii ix97 (.Y (L1_4_L2_4_G5_MINI_ALU_OperationResult_14), .A0 (Instr), .A1 (
            L1_4_L2_4_G5_MINI_ALU_BoothP_15)) ;
    nor02ii ix101 (.Y (L1_4_L2_4_G5_MINI_ALU_OperationResult_15), .A0 (Instr), .A1 (
            L1_4_L2_4_G5_MINI_ALU_BoothP_16)) ;
    mux21_ni ix1121 (.Y (L1_2_L2_1_G1_MINI_ALU_OperationResult_0), .A0 (
             L1_2_L2_1_G1_MINI_ALU_BoothP_1), .A1 (WindowDin_2__1__0), .S0 (
             Instr)) ;
    mux21_ni ix1129 (.Y (L1_2_L2_1_G1_MINI_ALU_OperationResult_1), .A0 (
             L1_2_L2_1_G1_MINI_ALU_BoothP_2), .A1 (WindowDin_2__1__1), .S0 (
             Instr)) ;
    mux21_ni ix1137 (.Y (L1_2_L2_1_G1_MINI_ALU_OperationResult_2), .A0 (
             L1_2_L2_1_G1_MINI_ALU_BoothP_3), .A1 (WindowDin_2__1__2), .S0 (
             Instr)) ;
    mux21_ni ix1145 (.Y (L1_2_L2_1_G1_MINI_ALU_OperationResult_3), .A0 (
             L1_2_L2_1_G1_MINI_ALU_BoothP_4), .A1 (WindowDin_2__1__3), .S0 (
             Instr)) ;
    mux21_ni ix1153 (.Y (L1_2_L2_1_G1_MINI_ALU_OperationResult_4), .A0 (
             L1_2_L2_1_G1_MINI_ALU_BoothP_5), .A1 (WindowDin_2__1__4), .S0 (
             Instr)) ;
    mux21_ni ix1161 (.Y (L1_2_L2_1_G1_MINI_ALU_OperationResult_5), .A0 (
             L1_2_L2_1_G1_MINI_ALU_BoothP_6), .A1 (WindowDin_2__1__5), .S0 (
             Instr)) ;
    mux21_ni ix1169 (.Y (L1_2_L2_1_G1_MINI_ALU_OperationResult_6), .A0 (
             L1_2_L2_1_G1_MINI_ALU_BoothP_7), .A1 (WindowDin_2__1__6), .S0 (
             Instr)) ;
    mux21_ni ix1177 (.Y (L1_2_L2_1_G1_MINI_ALU_OperationResult_7), .A0 (
             L1_2_L2_1_G1_MINI_ALU_BoothP_8), .A1 (WindowDin_2__1__7), .S0 (
             Instr)) ;
    nor02ii ix1085 (.Y (L1_2_L2_1_G1_MINI_ALU_OperationResult_8), .A0 (Instr), .A1 (
            L1_2_L2_1_G1_MINI_ALU_BoothP_9)) ;
    nor02ii ix1089 (.Y (L1_2_L2_1_G1_MINI_ALU_OperationResult_9), .A0 (Instr), .A1 (
            L1_2_L2_1_G1_MINI_ALU_BoothP_10)) ;
    nor02ii ix1093 (.Y (L1_2_L2_1_G1_MINI_ALU_OperationResult_10), .A0 (Instr), 
            .A1 (L1_2_L2_1_G1_MINI_ALU_BoothP_11)) ;
    nor02ii ix1097 (.Y (L1_2_L2_1_G1_MINI_ALU_OperationResult_11), .A0 (Instr), 
            .A1 (L1_2_L2_1_G1_MINI_ALU_BoothP_12)) ;
    nor02ii ix1101 (.Y (L1_2_L2_1_G1_MINI_ALU_OperationResult_12), .A0 (Instr), 
            .A1 (L1_2_L2_1_G1_MINI_ALU_BoothP_13)) ;
    nor02ii ix1105 (.Y (L1_2_L2_1_G1_MINI_ALU_OperationResult_13), .A0 (Instr), 
            .A1 (L1_2_L2_1_G1_MINI_ALU_BoothP_14)) ;
    nor02ii ix1109 (.Y (L1_2_L2_1_G1_MINI_ALU_OperationResult_14), .A0 (Instr), 
            .A1 (L1_2_L2_1_G1_MINI_ALU_BoothP_15)) ;
    nor02ii ix1113 (.Y (L1_2_L2_1_G1_MINI_ALU_OperationResult_15), .A0 (Instr), 
            .A1 (L1_2_L2_1_G1_MINI_ALU_BoothP_16)) ;
    mux21_ni ix1217 (.Y (L1_2_L2_0_G1_MINI_ALU_OperationResult_0), .A0 (
             L1_2_L2_0_G1_MINI_ALU_BoothP_1), .A1 (WindowDin_2__0__0), .S0 (
             Instr)) ;
    mux21_ni ix1225 (.Y (L1_2_L2_0_G1_MINI_ALU_OperationResult_1), .A0 (
             L1_2_L2_0_G1_MINI_ALU_BoothP_2), .A1 (WindowDin_2__0__1), .S0 (
             Instr)) ;
    mux21_ni ix1233 (.Y (L1_2_L2_0_G1_MINI_ALU_OperationResult_2), .A0 (
             L1_2_L2_0_G1_MINI_ALU_BoothP_3), .A1 (WindowDin_2__0__2), .S0 (
             Instr)) ;
    mux21_ni ix1241 (.Y (L1_2_L2_0_G1_MINI_ALU_OperationResult_3), .A0 (
             L1_2_L2_0_G1_MINI_ALU_BoothP_4), .A1 (WindowDin_2__0__3), .S0 (
             Instr)) ;
    mux21_ni ix1249 (.Y (L1_2_L2_0_G1_MINI_ALU_OperationResult_4), .A0 (
             L1_2_L2_0_G1_MINI_ALU_BoothP_5), .A1 (WindowDin_2__0__4), .S0 (
             Instr)) ;
    mux21_ni ix1257 (.Y (L1_2_L2_0_G1_MINI_ALU_OperationResult_5), .A0 (
             L1_2_L2_0_G1_MINI_ALU_BoothP_6), .A1 (WindowDin_2__0__5), .S0 (
             Instr)) ;
    mux21_ni ix1265 (.Y (L1_2_L2_0_G1_MINI_ALU_OperationResult_6), .A0 (
             L1_2_L2_0_G1_MINI_ALU_BoothP_7), .A1 (WindowDin_2__0__6), .S0 (
             Instr)) ;
    mux21_ni ix1273 (.Y (L1_2_L2_0_G1_MINI_ALU_OperationResult_7), .A0 (
             L1_2_L2_0_G1_MINI_ALU_BoothP_8), .A1 (WindowDin_2__0__7), .S0 (
             Instr)) ;
    nor02ii ix1181 (.Y (L1_2_L2_0_G1_MINI_ALU_OperationResult_8), .A0 (Instr), .A1 (
            L1_2_L2_0_G1_MINI_ALU_BoothP_9)) ;
    nor02ii ix1185 (.Y (L1_2_L2_0_G1_MINI_ALU_OperationResult_9), .A0 (Instr), .A1 (
            L1_2_L2_0_G1_MINI_ALU_BoothP_10)) ;
    nor02ii ix1189 (.Y (L1_2_L2_0_G1_MINI_ALU_OperationResult_10), .A0 (Instr), 
            .A1 (L1_2_L2_0_G1_MINI_ALU_BoothP_11)) ;
    nor02ii ix1193 (.Y (L1_2_L2_0_G1_MINI_ALU_OperationResult_11), .A0 (Instr), 
            .A1 (L1_2_L2_0_G1_MINI_ALU_BoothP_12)) ;
    nor02ii ix1197 (.Y (L1_2_L2_0_G1_MINI_ALU_OperationResult_12), .A0 (Instr), 
            .A1 (L1_2_L2_0_G1_MINI_ALU_BoothP_13)) ;
    nor02ii ix1201 (.Y (L1_2_L2_0_G1_MINI_ALU_OperationResult_13), .A0 (Instr), 
            .A1 (L1_2_L2_0_G1_MINI_ALU_BoothP_14)) ;
    nor02ii ix1205 (.Y (L1_2_L2_0_G1_MINI_ALU_OperationResult_14), .A0 (Instr), 
            .A1 (L1_2_L2_0_G1_MINI_ALU_BoothP_15)) ;
    nor02ii ix1209 (.Y (L1_2_L2_0_G1_MINI_ALU_OperationResult_15), .A0 (Instr), 
            .A1 (L1_2_L2_0_G1_MINI_ALU_BoothP_16)) ;
    mux21_ni ix1313 (.Y (L1_1_L2_4_G1_MINI_ALU_OperationResult_0), .A0 (
             L1_1_L2_4_G1_MINI_ALU_BoothP_1), .A1 (WindowDin_1__4__0), .S0 (
             Instr)) ;
    mux21_ni ix1321 (.Y (L1_1_L2_4_G1_MINI_ALU_OperationResult_1), .A0 (
             L1_1_L2_4_G1_MINI_ALU_BoothP_2), .A1 (WindowDin_1__4__1), .S0 (
             Instr)) ;
    mux21_ni ix1329 (.Y (L1_1_L2_4_G1_MINI_ALU_OperationResult_2), .A0 (
             L1_1_L2_4_G1_MINI_ALU_BoothP_3), .A1 (WindowDin_1__4__2), .S0 (
             Instr)) ;
    mux21_ni ix1337 (.Y (L1_1_L2_4_G1_MINI_ALU_OperationResult_3), .A0 (
             L1_1_L2_4_G1_MINI_ALU_BoothP_4), .A1 (WindowDin_1__4__3), .S0 (
             Instr)) ;
    mux21_ni ix1345 (.Y (L1_1_L2_4_G1_MINI_ALU_OperationResult_4), .A0 (
             L1_1_L2_4_G1_MINI_ALU_BoothP_5), .A1 (WindowDin_1__4__4), .S0 (
             Instr)) ;
    mux21_ni ix1353 (.Y (L1_1_L2_4_G1_MINI_ALU_OperationResult_5), .A0 (
             L1_1_L2_4_G1_MINI_ALU_BoothP_6), .A1 (WindowDin_1__4__5), .S0 (
             Instr)) ;
    mux21_ni ix1361 (.Y (L1_1_L2_4_G1_MINI_ALU_OperationResult_6), .A0 (
             L1_1_L2_4_G1_MINI_ALU_BoothP_7), .A1 (WindowDin_1__4__6), .S0 (
             Instr)) ;
    mux21_ni ix1369 (.Y (L1_1_L2_4_G1_MINI_ALU_OperationResult_7), .A0 (
             L1_1_L2_4_G1_MINI_ALU_BoothP_8), .A1 (WindowDin_1__4__7), .S0 (
             Instr)) ;
    nor02ii ix1277 (.Y (L1_1_L2_4_G1_MINI_ALU_OperationResult_8), .A0 (Instr), .A1 (
            L1_1_L2_4_G1_MINI_ALU_BoothP_9)) ;
    nor02ii ix1281 (.Y (L1_1_L2_4_G1_MINI_ALU_OperationResult_9), .A0 (Instr), .A1 (
            L1_1_L2_4_G1_MINI_ALU_BoothP_10)) ;
    nor02ii ix1285 (.Y (L1_1_L2_4_G1_MINI_ALU_OperationResult_10), .A0 (Instr), 
            .A1 (L1_1_L2_4_G1_MINI_ALU_BoothP_11)) ;
    nor02ii ix1289 (.Y (L1_1_L2_4_G1_MINI_ALU_OperationResult_11), .A0 (Instr), 
            .A1 (L1_1_L2_4_G1_MINI_ALU_BoothP_12)) ;
    nor02ii ix1293 (.Y (L1_1_L2_4_G1_MINI_ALU_OperationResult_12), .A0 (Instr), 
            .A1 (L1_1_L2_4_G1_MINI_ALU_BoothP_13)) ;
    nor02ii ix1297 (.Y (L1_1_L2_4_G1_MINI_ALU_OperationResult_13), .A0 (Instr), 
            .A1 (L1_1_L2_4_G1_MINI_ALU_BoothP_14)) ;
    nor02ii ix1301 (.Y (L1_1_L2_4_G1_MINI_ALU_OperationResult_14), .A0 (Instr), 
            .A1 (L1_1_L2_4_G1_MINI_ALU_BoothP_15)) ;
    nor02ii ix1305 (.Y (L1_1_L2_4_G1_MINI_ALU_OperationResult_15), .A0 (Instr), 
            .A1 (L1_1_L2_4_G1_MINI_ALU_BoothP_16)) ;
    mux21_ni ix1409 (.Y (L1_1_L2_3_G1_MINI_ALU_OperationResult_0), .A0 (
             L1_1_L2_3_G1_MINI_ALU_BoothP_1), .A1 (WindowDin_1__3__0), .S0 (
             Instr)) ;
    mux21_ni ix1417 (.Y (L1_1_L2_3_G1_MINI_ALU_OperationResult_1), .A0 (
             L1_1_L2_3_G1_MINI_ALU_BoothP_2), .A1 (WindowDin_1__3__1), .S0 (
             Instr)) ;
    mux21_ni ix1425 (.Y (L1_1_L2_3_G1_MINI_ALU_OperationResult_2), .A0 (
             L1_1_L2_3_G1_MINI_ALU_BoothP_3), .A1 (WindowDin_1__3__2), .S0 (
             Instr)) ;
    mux21_ni ix1433 (.Y (L1_1_L2_3_G1_MINI_ALU_OperationResult_3), .A0 (
             L1_1_L2_3_G1_MINI_ALU_BoothP_4), .A1 (WindowDin_1__3__3), .S0 (
             Instr)) ;
    mux21_ni ix1441 (.Y (L1_1_L2_3_G1_MINI_ALU_OperationResult_4), .A0 (
             L1_1_L2_3_G1_MINI_ALU_BoothP_5), .A1 (WindowDin_1__3__4), .S0 (
             Instr)) ;
    mux21_ni ix1449 (.Y (L1_1_L2_3_G1_MINI_ALU_OperationResult_5), .A0 (
             L1_1_L2_3_G1_MINI_ALU_BoothP_6), .A1 (WindowDin_1__3__5), .S0 (
             Instr)) ;
    mux21_ni ix1457 (.Y (L1_1_L2_3_G1_MINI_ALU_OperationResult_6), .A0 (
             L1_1_L2_3_G1_MINI_ALU_BoothP_7), .A1 (WindowDin_1__3__6), .S0 (
             Instr)) ;
    mux21_ni ix1465 (.Y (L1_1_L2_3_G1_MINI_ALU_OperationResult_7), .A0 (
             L1_1_L2_3_G1_MINI_ALU_BoothP_8), .A1 (WindowDin_1__3__7), .S0 (
             Instr)) ;
    nor02ii ix1373 (.Y (L1_1_L2_3_G1_MINI_ALU_OperationResult_8), .A0 (Instr), .A1 (
            L1_1_L2_3_G1_MINI_ALU_BoothP_9)) ;
    nor02ii ix1377 (.Y (L1_1_L2_3_G1_MINI_ALU_OperationResult_9), .A0 (Instr), .A1 (
            L1_1_L2_3_G1_MINI_ALU_BoothP_10)) ;
    nor02ii ix1381 (.Y (L1_1_L2_3_G1_MINI_ALU_OperationResult_10), .A0 (Instr), 
            .A1 (L1_1_L2_3_G1_MINI_ALU_BoothP_11)) ;
    nor02ii ix1385 (.Y (L1_1_L2_3_G1_MINI_ALU_OperationResult_11), .A0 (Instr), 
            .A1 (L1_1_L2_3_G1_MINI_ALU_BoothP_12)) ;
    nor02ii ix1389 (.Y (L1_1_L2_3_G1_MINI_ALU_OperationResult_12), .A0 (Instr), 
            .A1 (L1_1_L2_3_G1_MINI_ALU_BoothP_13)) ;
    nor02ii ix1393 (.Y (L1_1_L2_3_G1_MINI_ALU_OperationResult_13), .A0 (Instr), 
            .A1 (L1_1_L2_3_G1_MINI_ALU_BoothP_14)) ;
    nor02ii ix1397 (.Y (L1_1_L2_3_G1_MINI_ALU_OperationResult_14), .A0 (Instr), 
            .A1 (L1_1_L2_3_G1_MINI_ALU_BoothP_15)) ;
    nor02ii ix1401 (.Y (L1_1_L2_3_G1_MINI_ALU_OperationResult_15), .A0 (Instr), 
            .A1 (L1_1_L2_3_G1_MINI_ALU_BoothP_16)) ;
    mux21_ni ix1505 (.Y (L1_1_L2_2_G1_MINI_ALU_OperationResult_0), .A0 (
             L1_1_L2_2_G1_MINI_ALU_BoothP_1), .A1 (WindowDin_1__2__0), .S0 (
             Instr)) ;
    mux21_ni ix1513 (.Y (L1_1_L2_2_G1_MINI_ALU_OperationResult_1), .A0 (
             L1_1_L2_2_G1_MINI_ALU_BoothP_2), .A1 (WindowDin_1__2__1), .S0 (
             Instr)) ;
    mux21_ni ix1521 (.Y (L1_1_L2_2_G1_MINI_ALU_OperationResult_2), .A0 (
             L1_1_L2_2_G1_MINI_ALU_BoothP_3), .A1 (WindowDin_1__2__2), .S0 (
             Instr)) ;
    mux21_ni ix1529 (.Y (L1_1_L2_2_G1_MINI_ALU_OperationResult_3), .A0 (
             L1_1_L2_2_G1_MINI_ALU_BoothP_4), .A1 (WindowDin_1__2__3), .S0 (
             Instr)) ;
    mux21_ni ix1537 (.Y (L1_1_L2_2_G1_MINI_ALU_OperationResult_4), .A0 (
             L1_1_L2_2_G1_MINI_ALU_BoothP_5), .A1 (WindowDin_1__2__4), .S0 (
             Instr)) ;
    mux21_ni ix1545 (.Y (L1_1_L2_2_G1_MINI_ALU_OperationResult_5), .A0 (
             L1_1_L2_2_G1_MINI_ALU_BoothP_6), .A1 (WindowDin_1__2__5), .S0 (
             Instr)) ;
    mux21_ni ix1553 (.Y (L1_1_L2_2_G1_MINI_ALU_OperationResult_6), .A0 (
             L1_1_L2_2_G1_MINI_ALU_BoothP_7), .A1 (WindowDin_1__2__6), .S0 (
             Instr)) ;
    mux21_ni ix1561 (.Y (L1_1_L2_2_G1_MINI_ALU_OperationResult_7), .A0 (
             L1_1_L2_2_G1_MINI_ALU_BoothP_8), .A1 (WindowDin_1__2__7), .S0 (
             Instr)) ;
    nor02ii ix1469 (.Y (L1_1_L2_2_G1_MINI_ALU_OperationResult_8), .A0 (Instr), .A1 (
            L1_1_L2_2_G1_MINI_ALU_BoothP_9)) ;
    nor02ii ix1473 (.Y (L1_1_L2_2_G1_MINI_ALU_OperationResult_9), .A0 (Instr), .A1 (
            L1_1_L2_2_G1_MINI_ALU_BoothP_10)) ;
    nor02ii ix1477 (.Y (L1_1_L2_2_G1_MINI_ALU_OperationResult_10), .A0 (Instr), 
            .A1 (L1_1_L2_2_G1_MINI_ALU_BoothP_11)) ;
    nor02ii ix1481 (.Y (L1_1_L2_2_G1_MINI_ALU_OperationResult_11), .A0 (Instr), 
            .A1 (L1_1_L2_2_G1_MINI_ALU_BoothP_12)) ;
    nor02ii ix1485 (.Y (L1_1_L2_2_G1_MINI_ALU_OperationResult_12), .A0 (Instr), 
            .A1 (L1_1_L2_2_G1_MINI_ALU_BoothP_13)) ;
    nor02ii ix1489 (.Y (L1_1_L2_2_G1_MINI_ALU_OperationResult_13), .A0 (Instr), 
            .A1 (L1_1_L2_2_G1_MINI_ALU_BoothP_14)) ;
    nor02ii ix1493 (.Y (L1_1_L2_2_G1_MINI_ALU_OperationResult_14), .A0 (Instr), 
            .A1 (L1_1_L2_2_G1_MINI_ALU_BoothP_15)) ;
    nor02ii ix1497 (.Y (L1_1_L2_2_G1_MINI_ALU_OperationResult_15), .A0 (Instr), 
            .A1 (L1_1_L2_2_G1_MINI_ALU_BoothP_16)) ;
    mux21_ni ix1601 (.Y (L1_1_L2_1_G1_MINI_ALU_OperationResult_0), .A0 (
             L1_1_L2_1_G1_MINI_ALU_BoothP_1), .A1 (WindowDin_1__1__0), .S0 (
             Instr)) ;
    mux21_ni ix1609 (.Y (L1_1_L2_1_G1_MINI_ALU_OperationResult_1), .A0 (
             L1_1_L2_1_G1_MINI_ALU_BoothP_2), .A1 (WindowDin_1__1__1), .S0 (
             Instr)) ;
    mux21_ni ix1617 (.Y (L1_1_L2_1_G1_MINI_ALU_OperationResult_2), .A0 (
             L1_1_L2_1_G1_MINI_ALU_BoothP_3), .A1 (WindowDin_1__1__2), .S0 (
             Instr)) ;
    mux21_ni ix1625 (.Y (L1_1_L2_1_G1_MINI_ALU_OperationResult_3), .A0 (
             L1_1_L2_1_G1_MINI_ALU_BoothP_4), .A1 (WindowDin_1__1__3), .S0 (
             Instr)) ;
    mux21_ni ix1633 (.Y (L1_1_L2_1_G1_MINI_ALU_OperationResult_4), .A0 (
             L1_1_L2_1_G1_MINI_ALU_BoothP_5), .A1 (WindowDin_1__1__4), .S0 (
             Instr)) ;
    mux21_ni ix1641 (.Y (L1_1_L2_1_G1_MINI_ALU_OperationResult_5), .A0 (
             L1_1_L2_1_G1_MINI_ALU_BoothP_6), .A1 (WindowDin_1__1__5), .S0 (
             Instr)) ;
    mux21_ni ix1649 (.Y (L1_1_L2_1_G1_MINI_ALU_OperationResult_6), .A0 (
             L1_1_L2_1_G1_MINI_ALU_BoothP_7), .A1 (WindowDin_1__1__6), .S0 (
             Instr)) ;
    mux21_ni ix1657 (.Y (L1_1_L2_1_G1_MINI_ALU_OperationResult_7), .A0 (
             L1_1_L2_1_G1_MINI_ALU_BoothP_8), .A1 (WindowDin_1__1__7), .S0 (
             Instr)) ;
    nor02ii ix1565 (.Y (L1_1_L2_1_G1_MINI_ALU_OperationResult_8), .A0 (Instr), .A1 (
            L1_1_L2_1_G1_MINI_ALU_BoothP_9)) ;
    nor02ii ix1569 (.Y (L1_1_L2_1_G1_MINI_ALU_OperationResult_9), .A0 (Instr), .A1 (
            L1_1_L2_1_G1_MINI_ALU_BoothP_10)) ;
    nor02ii ix1573 (.Y (L1_1_L2_1_G1_MINI_ALU_OperationResult_10), .A0 (Instr), 
            .A1 (L1_1_L2_1_G1_MINI_ALU_BoothP_11)) ;
    nor02ii ix1577 (.Y (L1_1_L2_1_G1_MINI_ALU_OperationResult_11), .A0 (Instr), 
            .A1 (L1_1_L2_1_G1_MINI_ALU_BoothP_12)) ;
    nor02ii ix1581 (.Y (L1_1_L2_1_G1_MINI_ALU_OperationResult_12), .A0 (Instr), 
            .A1 (L1_1_L2_1_G1_MINI_ALU_BoothP_13)) ;
    nor02ii ix1585 (.Y (L1_1_L2_1_G1_MINI_ALU_OperationResult_13), .A0 (Instr), 
            .A1 (L1_1_L2_1_G1_MINI_ALU_BoothP_14)) ;
    nor02ii ix1589 (.Y (L1_1_L2_1_G1_MINI_ALU_OperationResult_14), .A0 (Instr), 
            .A1 (L1_1_L2_1_G1_MINI_ALU_BoothP_15)) ;
    nor02ii ix1593 (.Y (L1_1_L2_1_G1_MINI_ALU_OperationResult_15), .A0 (Instr), 
            .A1 (L1_1_L2_1_G1_MINI_ALU_BoothP_16)) ;
    mux21_ni ix1697 (.Y (L1_1_L2_0_G1_MINI_ALU_OperationResult_0), .A0 (
             L1_1_L2_0_G1_MINI_ALU_BoothP_1), .A1 (WindowDin_1__0__0), .S0 (
             Instr)) ;
    mux21_ni ix1705 (.Y (L1_1_L2_0_G1_MINI_ALU_OperationResult_1), .A0 (
             L1_1_L2_0_G1_MINI_ALU_BoothP_2), .A1 (WindowDin_1__0__1), .S0 (
             Instr)) ;
    mux21_ni ix1713 (.Y (L1_1_L2_0_G1_MINI_ALU_OperationResult_2), .A0 (
             L1_1_L2_0_G1_MINI_ALU_BoothP_3), .A1 (WindowDin_1__0__2), .S0 (
             Instr)) ;
    mux21_ni ix1721 (.Y (L1_1_L2_0_G1_MINI_ALU_OperationResult_3), .A0 (
             L1_1_L2_0_G1_MINI_ALU_BoothP_4), .A1 (WindowDin_1__0__3), .S0 (
             Instr)) ;
    mux21_ni ix1729 (.Y (L1_1_L2_0_G1_MINI_ALU_OperationResult_4), .A0 (
             L1_1_L2_0_G1_MINI_ALU_BoothP_5), .A1 (WindowDin_1__0__4), .S0 (
             Instr)) ;
    mux21_ni ix1737 (.Y (L1_1_L2_0_G1_MINI_ALU_OperationResult_5), .A0 (
             L1_1_L2_0_G1_MINI_ALU_BoothP_6), .A1 (WindowDin_1__0__5), .S0 (
             Instr)) ;
    mux21_ni ix1745 (.Y (L1_1_L2_0_G1_MINI_ALU_OperationResult_6), .A0 (
             L1_1_L2_0_G1_MINI_ALU_BoothP_7), .A1 (WindowDin_1__0__6), .S0 (
             Instr)) ;
    mux21_ni ix1753 (.Y (L1_1_L2_0_G1_MINI_ALU_OperationResult_7), .A0 (
             L1_1_L2_0_G1_MINI_ALU_BoothP_8), .A1 (WindowDin_1__0__7), .S0 (
             Instr)) ;
    nor02ii ix1661 (.Y (L1_1_L2_0_G1_MINI_ALU_OperationResult_8), .A0 (Instr), .A1 (
            L1_1_L2_0_G1_MINI_ALU_BoothP_9)) ;
    nor02ii ix1665 (.Y (L1_1_L2_0_G1_MINI_ALU_OperationResult_9), .A0 (Instr), .A1 (
            L1_1_L2_0_G1_MINI_ALU_BoothP_10)) ;
    nor02ii ix1669 (.Y (L1_1_L2_0_G1_MINI_ALU_OperationResult_10), .A0 (Instr), 
            .A1 (L1_1_L2_0_G1_MINI_ALU_BoothP_11)) ;
    nor02ii ix1673 (.Y (L1_1_L2_0_G1_MINI_ALU_OperationResult_11), .A0 (Instr), 
            .A1 (L1_1_L2_0_G1_MINI_ALU_BoothP_12)) ;
    nor02ii ix1677 (.Y (L1_1_L2_0_G1_MINI_ALU_OperationResult_12), .A0 (Instr), 
            .A1 (L1_1_L2_0_G1_MINI_ALU_BoothP_13)) ;
    nor02ii ix1681 (.Y (L1_1_L2_0_G1_MINI_ALU_OperationResult_13), .A0 (Instr), 
            .A1 (L1_1_L2_0_G1_MINI_ALU_BoothP_14)) ;
    nor02ii ix1685 (.Y (L1_1_L2_0_G1_MINI_ALU_OperationResult_14), .A0 (Instr), 
            .A1 (L1_1_L2_0_G1_MINI_ALU_BoothP_15)) ;
    nor02ii ix1689 (.Y (L1_1_L2_0_G1_MINI_ALU_OperationResult_15), .A0 (Instr), 
            .A1 (L1_1_L2_0_G1_MINI_ALU_BoothP_16)) ;
    mux21_ni ix1793 (.Y (L1_0_L2_4_G1_MINI_ALU_OperationResult_0), .A0 (
             L1_0_L2_4_G1_MINI_ALU_BoothP_1), .A1 (WindowDin_0__4__0), .S0 (
             Instr)) ;
    mux21_ni ix1801 (.Y (L1_0_L2_4_G1_MINI_ALU_OperationResult_1), .A0 (
             L1_0_L2_4_G1_MINI_ALU_BoothP_2), .A1 (WindowDin_0__4__1), .S0 (
             Instr)) ;
    mux21_ni ix1809 (.Y (L1_0_L2_4_G1_MINI_ALU_OperationResult_2), .A0 (
             L1_0_L2_4_G1_MINI_ALU_BoothP_3), .A1 (WindowDin_0__4__2), .S0 (
             Instr)) ;
    mux21_ni ix1817 (.Y (L1_0_L2_4_G1_MINI_ALU_OperationResult_3), .A0 (
             L1_0_L2_4_G1_MINI_ALU_BoothP_4), .A1 (WindowDin_0__4__3), .S0 (
             Instr)) ;
    mux21_ni ix1825 (.Y (L1_0_L2_4_G1_MINI_ALU_OperationResult_4), .A0 (
             L1_0_L2_4_G1_MINI_ALU_BoothP_5), .A1 (WindowDin_0__4__4), .S0 (
             Instr)) ;
    mux21_ni ix1833 (.Y (L1_0_L2_4_G1_MINI_ALU_OperationResult_5), .A0 (
             L1_0_L2_4_G1_MINI_ALU_BoothP_6), .A1 (WindowDin_0__4__5), .S0 (
             Instr)) ;
    mux21_ni ix1841 (.Y (L1_0_L2_4_G1_MINI_ALU_OperationResult_6), .A0 (
             L1_0_L2_4_G1_MINI_ALU_BoothP_7), .A1 (WindowDin_0__4__6), .S0 (
             Instr)) ;
    mux21_ni ix1849 (.Y (L1_0_L2_4_G1_MINI_ALU_OperationResult_7), .A0 (
             L1_0_L2_4_G1_MINI_ALU_BoothP_8), .A1 (WindowDin_0__4__7), .S0 (
             Instr)) ;
    nor02ii ix1757 (.Y (L1_0_L2_4_G1_MINI_ALU_OperationResult_8), .A0 (Instr), .A1 (
            L1_0_L2_4_G1_MINI_ALU_BoothP_9)) ;
    nor02ii ix1761 (.Y (L1_0_L2_4_G1_MINI_ALU_OperationResult_9), .A0 (Instr), .A1 (
            L1_0_L2_4_G1_MINI_ALU_BoothP_10)) ;
    nor02ii ix1765 (.Y (L1_0_L2_4_G1_MINI_ALU_OperationResult_10), .A0 (Instr), 
            .A1 (L1_0_L2_4_G1_MINI_ALU_BoothP_11)) ;
    nor02ii ix1769 (.Y (L1_0_L2_4_G1_MINI_ALU_OperationResult_11), .A0 (Instr), 
            .A1 (L1_0_L2_4_G1_MINI_ALU_BoothP_12)) ;
    nor02ii ix1773 (.Y (L1_0_L2_4_G1_MINI_ALU_OperationResult_12), .A0 (Instr), 
            .A1 (L1_0_L2_4_G1_MINI_ALU_BoothP_13)) ;
    nor02ii ix1777 (.Y (L1_0_L2_4_G1_MINI_ALU_OperationResult_13), .A0 (Instr), 
            .A1 (L1_0_L2_4_G1_MINI_ALU_BoothP_14)) ;
    nor02ii ix1781 (.Y (L1_0_L2_4_G1_MINI_ALU_OperationResult_14), .A0 (Instr), 
            .A1 (L1_0_L2_4_G1_MINI_ALU_BoothP_15)) ;
    nor02ii ix1785 (.Y (L1_0_L2_4_G1_MINI_ALU_OperationResult_15), .A0 (Instr), 
            .A1 (L1_0_L2_4_G1_MINI_ALU_BoothP_16)) ;
    mux21_ni ix1889 (.Y (L1_0_L2_3_G1_MINI_ALU_OperationResult_0), .A0 (
             L1_0_L2_3_G1_MINI_ALU_BoothP_1), .A1 (WindowDin_0__3__0), .S0 (
             Instr)) ;
    mux21_ni ix1897 (.Y (L1_0_L2_3_G1_MINI_ALU_OperationResult_1), .A0 (
             L1_0_L2_3_G1_MINI_ALU_BoothP_2), .A1 (WindowDin_0__3__1), .S0 (
             Instr)) ;
    mux21_ni ix1905 (.Y (L1_0_L2_3_G1_MINI_ALU_OperationResult_2), .A0 (
             L1_0_L2_3_G1_MINI_ALU_BoothP_3), .A1 (WindowDin_0__3__2), .S0 (
             Instr)) ;
    mux21_ni ix1913 (.Y (L1_0_L2_3_G1_MINI_ALU_OperationResult_3), .A0 (
             L1_0_L2_3_G1_MINI_ALU_BoothP_4), .A1 (WindowDin_0__3__3), .S0 (
             Instr)) ;
    mux21_ni ix1921 (.Y (L1_0_L2_3_G1_MINI_ALU_OperationResult_4), .A0 (
             L1_0_L2_3_G1_MINI_ALU_BoothP_5), .A1 (WindowDin_0__3__4), .S0 (
             Instr)) ;
    mux21_ni ix1929 (.Y (L1_0_L2_3_G1_MINI_ALU_OperationResult_5), .A0 (
             L1_0_L2_3_G1_MINI_ALU_BoothP_6), .A1 (WindowDin_0__3__5), .S0 (
             Instr)) ;
    mux21_ni ix1937 (.Y (L1_0_L2_3_G1_MINI_ALU_OperationResult_6), .A0 (
             L1_0_L2_3_G1_MINI_ALU_BoothP_7), .A1 (WindowDin_0__3__6), .S0 (
             Instr)) ;
    mux21_ni ix1945 (.Y (L1_0_L2_3_G1_MINI_ALU_OperationResult_7), .A0 (
             L1_0_L2_3_G1_MINI_ALU_BoothP_8), .A1 (WindowDin_0__3__7), .S0 (
             Instr)) ;
    nor02ii ix1853 (.Y (L1_0_L2_3_G1_MINI_ALU_OperationResult_8), .A0 (Instr), .A1 (
            L1_0_L2_3_G1_MINI_ALU_BoothP_9)) ;
    nor02ii ix1857 (.Y (L1_0_L2_3_G1_MINI_ALU_OperationResult_9), .A0 (Instr), .A1 (
            L1_0_L2_3_G1_MINI_ALU_BoothP_10)) ;
    nor02ii ix1861 (.Y (L1_0_L2_3_G1_MINI_ALU_OperationResult_10), .A0 (Instr), 
            .A1 (L1_0_L2_3_G1_MINI_ALU_BoothP_11)) ;
    nor02ii ix1865 (.Y (L1_0_L2_3_G1_MINI_ALU_OperationResult_11), .A0 (Instr), 
            .A1 (L1_0_L2_3_G1_MINI_ALU_BoothP_12)) ;
    nor02ii ix1869 (.Y (L1_0_L2_3_G1_MINI_ALU_OperationResult_12), .A0 (Instr), 
            .A1 (L1_0_L2_3_G1_MINI_ALU_BoothP_13)) ;
    nor02ii ix1873 (.Y (L1_0_L2_3_G1_MINI_ALU_OperationResult_13), .A0 (Instr), 
            .A1 (L1_0_L2_3_G1_MINI_ALU_BoothP_14)) ;
    nor02ii ix1877 (.Y (L1_0_L2_3_G1_MINI_ALU_OperationResult_14), .A0 (Instr), 
            .A1 (L1_0_L2_3_G1_MINI_ALU_BoothP_15)) ;
    nor02ii ix1881 (.Y (L1_0_L2_3_G1_MINI_ALU_OperationResult_15), .A0 (Instr), 
            .A1 (L1_0_L2_3_G1_MINI_ALU_BoothP_16)) ;
    mux21_ni ix1985 (.Y (L1_0_L2_2_G1_MINI_ALU_OperationResult_0), .A0 (
             L1_0_L2_2_G1_MINI_ALU_BoothP_1), .A1 (WindowDin_0__2__0), .S0 (
             Instr)) ;
    mux21_ni ix1993 (.Y (L1_0_L2_2_G1_MINI_ALU_OperationResult_1), .A0 (
             L1_0_L2_2_G1_MINI_ALU_BoothP_2), .A1 (WindowDin_0__2__1), .S0 (
             Instr)) ;
    mux21_ni ix2001 (.Y (L1_0_L2_2_G1_MINI_ALU_OperationResult_2), .A0 (
             L1_0_L2_2_G1_MINI_ALU_BoothP_3), .A1 (WindowDin_0__2__2), .S0 (
             Instr)) ;
    mux21_ni ix2009 (.Y (L1_0_L2_2_G1_MINI_ALU_OperationResult_3), .A0 (
             L1_0_L2_2_G1_MINI_ALU_BoothP_4), .A1 (WindowDin_0__2__3), .S0 (
             Instr)) ;
    mux21_ni ix2017 (.Y (L1_0_L2_2_G1_MINI_ALU_OperationResult_4), .A0 (
             L1_0_L2_2_G1_MINI_ALU_BoothP_5), .A1 (WindowDin_0__2__4), .S0 (
             Instr)) ;
    mux21_ni ix2025 (.Y (L1_0_L2_2_G1_MINI_ALU_OperationResult_5), .A0 (
             L1_0_L2_2_G1_MINI_ALU_BoothP_6), .A1 (WindowDin_0__2__5), .S0 (
             Instr)) ;
    mux21_ni ix2033 (.Y (L1_0_L2_2_G1_MINI_ALU_OperationResult_6), .A0 (
             L1_0_L2_2_G1_MINI_ALU_BoothP_7), .A1 (WindowDin_0__2__6), .S0 (
             Instr)) ;
    mux21_ni ix2041 (.Y (L1_0_L2_2_G1_MINI_ALU_OperationResult_7), .A0 (
             L1_0_L2_2_G1_MINI_ALU_BoothP_8), .A1 (WindowDin_0__2__7), .S0 (
             Instr)) ;
    nor02ii ix1949 (.Y (L1_0_L2_2_G1_MINI_ALU_OperationResult_8), .A0 (Instr), .A1 (
            L1_0_L2_2_G1_MINI_ALU_BoothP_9)) ;
    nor02ii ix1953 (.Y (L1_0_L2_2_G1_MINI_ALU_OperationResult_9), .A0 (Instr), .A1 (
            L1_0_L2_2_G1_MINI_ALU_BoothP_10)) ;
    nor02ii ix1957 (.Y (L1_0_L2_2_G1_MINI_ALU_OperationResult_10), .A0 (Instr), 
            .A1 (L1_0_L2_2_G1_MINI_ALU_BoothP_11)) ;
    nor02ii ix1961 (.Y (L1_0_L2_2_G1_MINI_ALU_OperationResult_11), .A0 (Instr), 
            .A1 (L1_0_L2_2_G1_MINI_ALU_BoothP_12)) ;
    nor02ii ix1965 (.Y (L1_0_L2_2_G1_MINI_ALU_OperationResult_12), .A0 (Instr), 
            .A1 (L1_0_L2_2_G1_MINI_ALU_BoothP_13)) ;
    nor02ii ix1969 (.Y (L1_0_L2_2_G1_MINI_ALU_OperationResult_13), .A0 (Instr), 
            .A1 (L1_0_L2_2_G1_MINI_ALU_BoothP_14)) ;
    nor02ii ix1973 (.Y (L1_0_L2_2_G1_MINI_ALU_OperationResult_14), .A0 (Instr), 
            .A1 (L1_0_L2_2_G1_MINI_ALU_BoothP_15)) ;
    nor02ii ix1977 (.Y (L1_0_L2_2_G1_MINI_ALU_OperationResult_15), .A0 (Instr), 
            .A1 (L1_0_L2_2_G1_MINI_ALU_BoothP_16)) ;
    mux21_ni ix2081 (.Y (L1_0_L2_1_G1_MINI_ALU_OperationResult_0), .A0 (
             L1_0_L2_1_G1_MINI_ALU_BoothP_1), .A1 (WindowDin_0__1__0), .S0 (
             Instr)) ;
    mux21_ni ix2089 (.Y (L1_0_L2_1_G1_MINI_ALU_OperationResult_1), .A0 (
             L1_0_L2_1_G1_MINI_ALU_BoothP_2), .A1 (WindowDin_0__1__1), .S0 (
             Instr)) ;
    mux21_ni ix2097 (.Y (L1_0_L2_1_G1_MINI_ALU_OperationResult_2), .A0 (
             L1_0_L2_1_G1_MINI_ALU_BoothP_3), .A1 (WindowDin_0__1__2), .S0 (
             Instr)) ;
    mux21_ni ix2105 (.Y (L1_0_L2_1_G1_MINI_ALU_OperationResult_3), .A0 (
             L1_0_L2_1_G1_MINI_ALU_BoothP_4), .A1 (WindowDin_0__1__3), .S0 (
             Instr)) ;
    mux21_ni ix2113 (.Y (L1_0_L2_1_G1_MINI_ALU_OperationResult_4), .A0 (
             L1_0_L2_1_G1_MINI_ALU_BoothP_5), .A1 (WindowDin_0__1__4), .S0 (
             Instr)) ;
    mux21_ni ix2121 (.Y (L1_0_L2_1_G1_MINI_ALU_OperationResult_5), .A0 (
             L1_0_L2_1_G1_MINI_ALU_BoothP_6), .A1 (WindowDin_0__1__5), .S0 (
             Instr)) ;
    mux21_ni ix2129 (.Y (L1_0_L2_1_G1_MINI_ALU_OperationResult_6), .A0 (
             L1_0_L2_1_G1_MINI_ALU_BoothP_7), .A1 (WindowDin_0__1__6), .S0 (
             Instr)) ;
    mux21_ni ix2137 (.Y (L1_0_L2_1_G1_MINI_ALU_OperationResult_7), .A0 (
             L1_0_L2_1_G1_MINI_ALU_BoothP_8), .A1 (WindowDin_0__1__7), .S0 (
             Instr)) ;
    nor02ii ix2045 (.Y (L1_0_L2_1_G1_MINI_ALU_OperationResult_8), .A0 (Instr), .A1 (
            L1_0_L2_1_G1_MINI_ALU_BoothP_9)) ;
    nor02ii ix2049 (.Y (L1_0_L2_1_G1_MINI_ALU_OperationResult_9), .A0 (Instr), .A1 (
            L1_0_L2_1_G1_MINI_ALU_BoothP_10)) ;
    nor02ii ix2053 (.Y (L1_0_L2_1_G1_MINI_ALU_OperationResult_10), .A0 (Instr), 
            .A1 (L1_0_L2_1_G1_MINI_ALU_BoothP_11)) ;
    nor02ii ix2057 (.Y (L1_0_L2_1_G1_MINI_ALU_OperationResult_11), .A0 (Instr), 
            .A1 (L1_0_L2_1_G1_MINI_ALU_BoothP_12)) ;
    nor02ii ix2061 (.Y (L1_0_L2_1_G1_MINI_ALU_OperationResult_12), .A0 (Instr), 
            .A1 (L1_0_L2_1_G1_MINI_ALU_BoothP_13)) ;
    nor02ii ix2065 (.Y (L1_0_L2_1_G1_MINI_ALU_OperationResult_13), .A0 (Instr), 
            .A1 (L1_0_L2_1_G1_MINI_ALU_BoothP_14)) ;
    nor02ii ix2069 (.Y (L1_0_L2_1_G1_MINI_ALU_OperationResult_14), .A0 (Instr), 
            .A1 (L1_0_L2_1_G1_MINI_ALU_BoothP_15)) ;
    nor02ii ix2073 (.Y (L1_0_L2_1_G1_MINI_ALU_OperationResult_15), .A0 (Instr), 
            .A1 (L1_0_L2_1_G1_MINI_ALU_BoothP_16)) ;
    mux21_ni ix2177 (.Y (L1_0_L2_0_G1_MINI_ALU_OperationResult_0), .A0 (
             L1_0_L2_0_G1_MINI_ALU_BoothP_1), .A1 (WindowDin_0__0__0), .S0 (
             Instr)) ;
    mux21_ni ix2185 (.Y (L1_0_L2_0_G1_MINI_ALU_OperationResult_1), .A0 (
             L1_0_L2_0_G1_MINI_ALU_BoothP_2), .A1 (WindowDin_0__0__1), .S0 (
             Instr)) ;
    mux21_ni ix2193 (.Y (L1_0_L2_0_G1_MINI_ALU_OperationResult_2), .A0 (
             L1_0_L2_0_G1_MINI_ALU_BoothP_3), .A1 (WindowDin_0__0__2), .S0 (
             Instr)) ;
    mux21_ni ix2201 (.Y (L1_0_L2_0_G1_MINI_ALU_OperationResult_3), .A0 (
             L1_0_L2_0_G1_MINI_ALU_BoothP_4), .A1 (WindowDin_0__0__3), .S0 (
             Instr)) ;
    mux21_ni ix2209 (.Y (L1_0_L2_0_G1_MINI_ALU_OperationResult_4), .A0 (
             L1_0_L2_0_G1_MINI_ALU_BoothP_5), .A1 (WindowDin_0__0__4), .S0 (
             Instr)) ;
    mux21_ni ix2217 (.Y (L1_0_L2_0_G1_MINI_ALU_OperationResult_5), .A0 (
             L1_0_L2_0_G1_MINI_ALU_BoothP_6), .A1 (WindowDin_0__0__5), .S0 (
             Instr)) ;
    mux21_ni ix2225 (.Y (L1_0_L2_0_G1_MINI_ALU_OperationResult_6), .A0 (
             L1_0_L2_0_G1_MINI_ALU_BoothP_7), .A1 (WindowDin_0__0__6), .S0 (
             Instr)) ;
    mux21_ni ix2233 (.Y (L1_0_L2_0_G1_MINI_ALU_OperationResult_7), .A0 (
             L1_0_L2_0_G1_MINI_ALU_BoothP_8), .A1 (WindowDin_0__0__7), .S0 (
             Instr)) ;
    nor02ii ix2141 (.Y (L1_0_L2_0_G1_MINI_ALU_OperationResult_8), .A0 (Instr), .A1 (
            L1_0_L2_0_G1_MINI_ALU_BoothP_9)) ;
    nor02ii ix2145 (.Y (L1_0_L2_0_G1_MINI_ALU_OperationResult_9), .A0 (Instr), .A1 (
            L1_0_L2_0_G1_MINI_ALU_BoothP_10)) ;
    nor02ii ix2149 (.Y (L1_0_L2_0_G1_MINI_ALU_OperationResult_10), .A0 (Instr), 
            .A1 (L1_0_L2_0_G1_MINI_ALU_BoothP_11)) ;
    nor02ii ix2153 (.Y (L1_0_L2_0_G1_MINI_ALU_OperationResult_11), .A0 (Instr), 
            .A1 (L1_0_L2_0_G1_MINI_ALU_BoothP_12)) ;
    nor02ii ix2157 (.Y (L1_0_L2_0_G1_MINI_ALU_OperationResult_12), .A0 (Instr), 
            .A1 (L1_0_L2_0_G1_MINI_ALU_BoothP_13)) ;
    nor02ii ix2161 (.Y (L1_0_L2_0_G1_MINI_ALU_OperationResult_13), .A0 (Instr), 
            .A1 (L1_0_L2_0_G1_MINI_ALU_BoothP_14)) ;
    nor02ii ix2165 (.Y (L1_0_L2_0_G1_MINI_ALU_OperationResult_14), .A0 (Instr), 
            .A1 (L1_0_L2_0_G1_MINI_ALU_BoothP_15)) ;
    nor02ii ix2169 (.Y (L1_0_L2_0_G1_MINI_ALU_OperationResult_15), .A0 (Instr), 
            .A1 (L1_0_L2_0_G1_MINI_ALU_BoothP_16)) ;
    mux21_ni ix973 (.Y (L1FirstOperands_11__0), .A0 (
             L1_2_L2_2_G1_MINI_ALU_BoothP_1), .A1 (WindowDin_2__2__0), .S0 (
             Instr)) ;
    mux21_ni ix981 (.Y (L1FirstOperands_11__1), .A0 (
             L1_2_L2_2_G1_MINI_ALU_BoothP_2), .A1 (WindowDin_2__2__1), .S0 (
             Instr)) ;
    mux21_ni ix989 (.Y (L1FirstOperands_11__2), .A0 (
             L1_2_L2_2_G1_MINI_ALU_BoothP_3), .A1 (WindowDin_2__2__2), .S0 (
             Instr)) ;
    mux21_ni ix997 (.Y (L1FirstOperands_11__3), .A0 (
             L1_2_L2_2_G1_MINI_ALU_BoothP_4), .A1 (WindowDin_2__2__3), .S0 (
             Instr)) ;
    mux21_ni ix1005 (.Y (L1FirstOperands_11__4), .A0 (
             L1_2_L2_2_G1_MINI_ALU_BoothP_5), .A1 (WindowDin_2__2__4), .S0 (
             Instr)) ;
    mux21_ni ix1013 (.Y (L1FirstOperands_11__5), .A0 (
             L1_2_L2_2_G1_MINI_ALU_BoothP_6), .A1 (WindowDin_2__2__5), .S0 (
             Instr)) ;
    mux21_ni ix1021 (.Y (L1FirstOperands_11__6), .A0 (
             L1_2_L2_2_G1_MINI_ALU_BoothP_7), .A1 (WindowDin_2__2__6), .S0 (
             Instr)) ;
    mux21_ni ix1029 (.Y (L1FirstOperands_11__7), .A0 (
             L1_2_L2_2_G1_MINI_ALU_BoothP_8), .A1 (WindowDin_2__2__7), .S0 (
             Instr)) ;
    nor02ii ix937 (.Y (L1FirstOperands_11__8), .A0 (Instr), .A1 (
            L1_2_L2_2_G1_MINI_ALU_BoothP_9)) ;
    nor02ii ix941 (.Y (L1FirstOperands_11__9), .A0 (Instr), .A1 (
            L1_2_L2_2_G1_MINI_ALU_BoothP_10)) ;
    nor02ii ix945 (.Y (L1FirstOperands_11__10), .A0 (Instr), .A1 (
            L1_2_L2_2_G1_MINI_ALU_BoothP_11)) ;
    nor02ii ix949 (.Y (L1FirstOperands_11__11), .A0 (Instr), .A1 (
            L1_2_L2_2_G1_MINI_ALU_BoothP_12)) ;
    nor02ii ix953 (.Y (L1FirstOperands_11__12), .A0 (Instr), .A1 (
            L1_2_L2_2_G1_MINI_ALU_BoothP_13)) ;
    nor02ii ix957 (.Y (L1FirstOperands_11__13), .A0 (Instr), .A1 (
            L1_2_L2_2_G1_MINI_ALU_BoothP_14)) ;
    nor02ii ix961 (.Y (L1FirstOperands_11__14), .A0 (Instr), .A1 (
            L1_2_L2_2_G1_MINI_ALU_BoothP_15)) ;
    nor02ii ix965 (.Y (L1FirstOperands_11__15), .A0 (Instr), .A1 (
            L1_2_L2_2_G1_MINI_ALU_BoothP_16)) ;
    mux21_ni ix397 (.Y (L1FirstOperands_10__0), .A0 (
             L1_3_L2_3_G2_MINI_ALU_BoothP_1), .A1 (WindowDin_3__3__0), .S0 (
             Instr)) ;
    mux21_ni ix405 (.Y (L1FirstOperands_10__1), .A0 (
             L1_3_L2_3_G2_MINI_ALU_BoothP_2), .A1 (WindowDin_3__3__1), .S0 (
             Instr)) ;
    mux21_ni ix413 (.Y (L1FirstOperands_10__2), .A0 (
             L1_3_L2_3_G2_MINI_ALU_BoothP_3), .A1 (WindowDin_3__3__2), .S0 (
             Instr)) ;
    mux21_ni ix421 (.Y (L1FirstOperands_10__3), .A0 (
             L1_3_L2_3_G2_MINI_ALU_BoothP_4), .A1 (WindowDin_3__3__3), .S0 (
             Instr)) ;
    mux21_ni ix429 (.Y (L1FirstOperands_10__4), .A0 (
             L1_3_L2_3_G2_MINI_ALU_BoothP_5), .A1 (WindowDin_3__3__4), .S0 (
             Instr)) ;
    mux21_ni ix437 (.Y (L1FirstOperands_10__5), .A0 (
             L1_3_L2_3_G2_MINI_ALU_BoothP_6), .A1 (WindowDin_3__3__5), .S0 (
             Instr)) ;
    mux21_ni ix445 (.Y (L1FirstOperands_10__6), .A0 (
             L1_3_L2_3_G2_MINI_ALU_BoothP_7), .A1 (WindowDin_3__3__6), .S0 (
             Instr)) ;
    mux21_ni ix453 (.Y (L1FirstOperands_10__7), .A0 (
             L1_3_L2_3_G2_MINI_ALU_BoothP_8), .A1 (WindowDin_3__3__7), .S0 (
             Instr)) ;
    nor02ii ix361 (.Y (L1FirstOperands_10__8), .A0 (Instr), .A1 (
            L1_3_L2_3_G2_MINI_ALU_BoothP_9)) ;
    nor02ii ix365 (.Y (L1FirstOperands_10__9), .A0 (Instr), .A1 (
            L1_3_L2_3_G2_MINI_ALU_BoothP_10)) ;
    nor02ii ix369 (.Y (L1FirstOperands_10__10), .A0 (Instr), .A1 (
            L1_3_L2_3_G2_MINI_ALU_BoothP_11)) ;
    nor02ii ix373 (.Y (L1FirstOperands_10__11), .A0 (Instr), .A1 (
            L1_3_L2_3_G2_MINI_ALU_BoothP_12)) ;
    nor02ii ix377 (.Y (L1FirstOperands_10__12), .A0 (Instr), .A1 (
            L1_3_L2_3_G2_MINI_ALU_BoothP_13)) ;
    nor02ii ix381 (.Y (L1FirstOperands_10__13), .A0 (Instr), .A1 (
            L1_3_L2_3_G2_MINI_ALU_BoothP_14)) ;
    nor02ii ix385 (.Y (L1FirstOperands_10__14), .A0 (Instr), .A1 (
            L1_3_L2_3_G2_MINI_ALU_BoothP_15)) ;
    nor02ii ix389 (.Y (L1FirstOperands_10__15), .A0 (Instr), .A1 (
            L1_3_L2_3_G2_MINI_ALU_BoothP_16)) ;
    mux21_ni ix493 (.Y (L1FirstOperands_8__0), .A0 (
             L1_3_L2_2_G2_MINI_ALU_BoothP_1), .A1 (WindowDin_3__2__0), .S0 (
             Instr)) ;
    mux21_ni ix501 (.Y (L1FirstOperands_8__1), .A0 (
             L1_3_L2_2_G2_MINI_ALU_BoothP_2), .A1 (WindowDin_3__2__1), .S0 (
             Instr)) ;
    mux21_ni ix509 (.Y (L1FirstOperands_8__2), .A0 (
             L1_3_L2_2_G2_MINI_ALU_BoothP_3), .A1 (WindowDin_3__2__2), .S0 (
             Instr)) ;
    mux21_ni ix517 (.Y (L1FirstOperands_8__3), .A0 (
             L1_3_L2_2_G2_MINI_ALU_BoothP_4), .A1 (WindowDin_3__2__3), .S0 (
             Instr)) ;
    mux21_ni ix525 (.Y (L1FirstOperands_8__4), .A0 (
             L1_3_L2_2_G2_MINI_ALU_BoothP_5), .A1 (WindowDin_3__2__4), .S0 (
             Instr)) ;
    mux21_ni ix533 (.Y (L1FirstOperands_8__5), .A0 (
             L1_3_L2_2_G2_MINI_ALU_BoothP_6), .A1 (WindowDin_3__2__5), .S0 (
             Instr)) ;
    mux21_ni ix541 (.Y (L1FirstOperands_8__6), .A0 (
             L1_3_L2_2_G2_MINI_ALU_BoothP_7), .A1 (WindowDin_3__2__6), .S0 (
             Instr)) ;
    mux21_ni ix549 (.Y (L1FirstOperands_8__7), .A0 (
             L1_3_L2_2_G2_MINI_ALU_BoothP_8), .A1 (WindowDin_3__2__7), .S0 (
             Instr)) ;
    nor02ii ix457 (.Y (L1FirstOperands_8__8), .A0 (Instr), .A1 (
            L1_3_L2_2_G2_MINI_ALU_BoothP_9)) ;
    nor02ii ix461 (.Y (L1FirstOperands_8__9), .A0 (Instr), .A1 (
            L1_3_L2_2_G2_MINI_ALU_BoothP_10)) ;
    nor02ii ix465 (.Y (L1FirstOperands_8__10), .A0 (Instr), .A1 (
            L1_3_L2_2_G2_MINI_ALU_BoothP_11)) ;
    nor02ii ix469 (.Y (L1FirstOperands_8__11), .A0 (Instr), .A1 (
            L1_3_L2_2_G2_MINI_ALU_BoothP_12)) ;
    nor02ii ix473 (.Y (L1FirstOperands_8__12), .A0 (Instr), .A1 (
            L1_3_L2_2_G2_MINI_ALU_BoothP_13)) ;
    nor02ii ix477 (.Y (L1FirstOperands_8__13), .A0 (Instr), .A1 (
            L1_3_L2_2_G2_MINI_ALU_BoothP_14)) ;
    nor02ii ix481 (.Y (L1FirstOperands_8__14), .A0 (Instr), .A1 (
            L1_3_L2_2_G2_MINI_ALU_BoothP_15)) ;
    nor02ii ix485 (.Y (L1FirstOperands_8__15), .A0 (Instr), .A1 (
            L1_3_L2_2_G2_MINI_ALU_BoothP_16)) ;
    mux21_ni ix205 (.Y (L1FirstOperands_7__0), .A0 (
             L1_4_L2_3_G5_MINI_ALU_BoothP_1), .A1 (WindowDin_4__3__0), .S0 (
             Instr)) ;
    mux21_ni ix213 (.Y (L1FirstOperands_7__1), .A0 (
             L1_4_L2_3_G5_MINI_ALU_BoothP_2), .A1 (WindowDin_4__3__1), .S0 (
             Instr)) ;
    mux21_ni ix221 (.Y (L1FirstOperands_7__2), .A0 (
             L1_4_L2_3_G5_MINI_ALU_BoothP_3), .A1 (WindowDin_4__3__2), .S0 (
             Instr)) ;
    mux21_ni ix229 (.Y (L1FirstOperands_7__3), .A0 (
             L1_4_L2_3_G5_MINI_ALU_BoothP_4), .A1 (WindowDin_4__3__3), .S0 (
             Instr)) ;
    mux21_ni ix237 (.Y (L1FirstOperands_7__4), .A0 (
             L1_4_L2_3_G5_MINI_ALU_BoothP_5), .A1 (WindowDin_4__3__4), .S0 (
             Instr)) ;
    mux21_ni ix245 (.Y (L1FirstOperands_7__5), .A0 (
             L1_4_L2_3_G5_MINI_ALU_BoothP_6), .A1 (WindowDin_4__3__5), .S0 (
             Instr)) ;
    mux21_ni ix253 (.Y (L1FirstOperands_7__6), .A0 (
             L1_4_L2_3_G5_MINI_ALU_BoothP_7), .A1 (WindowDin_4__3__6), .S0 (
             Instr)) ;
    mux21_ni ix261 (.Y (L1FirstOperands_7__7), .A0 (
             L1_4_L2_3_G5_MINI_ALU_BoothP_8), .A1 (WindowDin_4__3__7), .S0 (
             Instr)) ;
    nor02ii ix169 (.Y (L1FirstOperands_7__8), .A0 (Instr), .A1 (
            L1_4_L2_3_G5_MINI_ALU_BoothP_9)) ;
    nor02ii ix173 (.Y (L1FirstOperands_7__9), .A0 (Instr), .A1 (
            L1_4_L2_3_G5_MINI_ALU_BoothP_10)) ;
    nor02ii ix177 (.Y (L1FirstOperands_7__10), .A0 (Instr), .A1 (
            L1_4_L2_3_G5_MINI_ALU_BoothP_11)) ;
    nor02ii ix181 (.Y (L1FirstOperands_7__11), .A0 (Instr), .A1 (
            L1_4_L2_3_G5_MINI_ALU_BoothP_12)) ;
    nor02ii ix185 (.Y (L1FirstOperands_7__12), .A0 (Instr), .A1 (
            L1_4_L2_3_G5_MINI_ALU_BoothP_13)) ;
    nor02ii ix189 (.Y (L1FirstOperands_7__13), .A0 (Instr), .A1 (
            L1_4_L2_3_G5_MINI_ALU_BoothP_14)) ;
    nor02ii ix193 (.Y (L1FirstOperands_7__14), .A0 (Instr), .A1 (
            L1_4_L2_3_G5_MINI_ALU_BoothP_15)) ;
    nor02ii ix197 (.Y (L1FirstOperands_7__15), .A0 (Instr), .A1 (
            L1_4_L2_3_G5_MINI_ALU_BoothP_16)) ;
    mux21_ni ix589 (.Y (L1FirstOperands_6__0), .A0 (
             L1_3_L2_1_G2_MINI_ALU_BoothP_1), .A1 (WindowDin_3__1__0), .S0 (
             Instr)) ;
    mux21_ni ix597 (.Y (L1FirstOperands_6__1), .A0 (
             L1_3_L2_1_G2_MINI_ALU_BoothP_2), .A1 (WindowDin_3__1__1), .S0 (
             Instr)) ;
    mux21_ni ix605 (.Y (L1FirstOperands_6__2), .A0 (
             L1_3_L2_1_G2_MINI_ALU_BoothP_3), .A1 (WindowDin_3__1__2), .S0 (
             Instr)) ;
    mux21_ni ix613 (.Y (L1FirstOperands_6__3), .A0 (
             L1_3_L2_1_G2_MINI_ALU_BoothP_4), .A1 (WindowDin_3__1__3), .S0 (
             Instr)) ;
    mux21_ni ix621 (.Y (L1FirstOperands_6__4), .A0 (
             L1_3_L2_1_G2_MINI_ALU_BoothP_5), .A1 (WindowDin_3__1__4), .S0 (
             Instr)) ;
    mux21_ni ix629 (.Y (L1FirstOperands_6__5), .A0 (
             L1_3_L2_1_G2_MINI_ALU_BoothP_6), .A1 (WindowDin_3__1__5), .S0 (
             Instr)) ;
    mux21_ni ix637 (.Y (L1FirstOperands_6__6), .A0 (
             L1_3_L2_1_G2_MINI_ALU_BoothP_7), .A1 (WindowDin_3__1__6), .S0 (
             Instr)) ;
    mux21_ni ix645 (.Y (L1FirstOperands_6__7), .A0 (
             L1_3_L2_1_G2_MINI_ALU_BoothP_8), .A1 (WindowDin_3__1__7), .S0 (
             Instr)) ;
    nor02ii ix553 (.Y (L1FirstOperands_6__8), .A0 (Instr), .A1 (
            L1_3_L2_1_G2_MINI_ALU_BoothP_9)) ;
    nor02ii ix557 (.Y (L1FirstOperands_6__9), .A0 (Instr), .A1 (
            L1_3_L2_1_G2_MINI_ALU_BoothP_10)) ;
    nor02ii ix561 (.Y (L1FirstOperands_6__10), .A0 (Instr), .A1 (
            L1_3_L2_1_G2_MINI_ALU_BoothP_11)) ;
    nor02ii ix565 (.Y (L1FirstOperands_6__11), .A0 (Instr), .A1 (
            L1_3_L2_1_G2_MINI_ALU_BoothP_12)) ;
    nor02ii ix569 (.Y (L1FirstOperands_6__12), .A0 (Instr), .A1 (
            L1_3_L2_1_G2_MINI_ALU_BoothP_13)) ;
    nor02ii ix573 (.Y (L1FirstOperands_6__13), .A0 (Instr), .A1 (
            L1_3_L2_1_G2_MINI_ALU_BoothP_14)) ;
    nor02ii ix577 (.Y (L1FirstOperands_6__14), .A0 (Instr), .A1 (
            L1_3_L2_1_G2_MINI_ALU_BoothP_15)) ;
    nor02ii ix581 (.Y (L1FirstOperands_6__15), .A0 (Instr), .A1 (
            L1_3_L2_1_G2_MINI_ALU_BoothP_16)) ;
    mux21_ni ix685 (.Y (L1FirstOperands_4__0), .A0 (
             L1_3_L2_0_G2_MINI_ALU_BoothP_1), .A1 (WindowDin_3__0__0), .S0 (
             Instr)) ;
    mux21_ni ix693 (.Y (L1FirstOperands_4__1), .A0 (
             L1_3_L2_0_G2_MINI_ALU_BoothP_2), .A1 (WindowDin_3__0__1), .S0 (
             Instr)) ;
    mux21_ni ix701 (.Y (L1FirstOperands_4__2), .A0 (
             L1_3_L2_0_G2_MINI_ALU_BoothP_3), .A1 (WindowDin_3__0__2), .S0 (
             Instr)) ;
    mux21_ni ix709 (.Y (L1FirstOperands_4__3), .A0 (
             L1_3_L2_0_G2_MINI_ALU_BoothP_4), .A1 (WindowDin_3__0__3), .S0 (
             Instr)) ;
    mux21_ni ix717 (.Y (L1FirstOperands_4__4), .A0 (
             L1_3_L2_0_G2_MINI_ALU_BoothP_5), .A1 (WindowDin_3__0__4), .S0 (
             Instr)) ;
    mux21_ni ix725 (.Y (L1FirstOperands_4__5), .A0 (
             L1_3_L2_0_G2_MINI_ALU_BoothP_6), .A1 (WindowDin_3__0__5), .S0 (
             Instr)) ;
    mux21_ni ix733 (.Y (L1FirstOperands_4__6), .A0 (
             L1_3_L2_0_G2_MINI_ALU_BoothP_7), .A1 (WindowDin_3__0__6), .S0 (
             Instr)) ;
    mux21_ni ix741 (.Y (L1FirstOperands_4__7), .A0 (
             L1_3_L2_0_G2_MINI_ALU_BoothP_8), .A1 (WindowDin_3__0__7), .S0 (
             Instr)) ;
    nor02ii ix649 (.Y (L1FirstOperands_4__8), .A0 (Instr), .A1 (
            L1_3_L2_0_G2_MINI_ALU_BoothP_9)) ;
    nor02ii ix653 (.Y (L1FirstOperands_4__9), .A0 (Instr), .A1 (
            L1_3_L2_0_G2_MINI_ALU_BoothP_10)) ;
    nor02ii ix657 (.Y (L1FirstOperands_4__10), .A0 (Instr), .A1 (
            L1_3_L2_0_G2_MINI_ALU_BoothP_11)) ;
    nor02ii ix661 (.Y (L1FirstOperands_4__11), .A0 (Instr), .A1 (
            L1_3_L2_0_G2_MINI_ALU_BoothP_12)) ;
    nor02ii ix665 (.Y (L1FirstOperands_4__12), .A0 (Instr), .A1 (
            L1_3_L2_0_G2_MINI_ALU_BoothP_13)) ;
    nor02ii ix669 (.Y (L1FirstOperands_4__13), .A0 (Instr), .A1 (
            L1_3_L2_0_G2_MINI_ALU_BoothP_14)) ;
    nor02ii ix673 (.Y (L1FirstOperands_4__14), .A0 (Instr), .A1 (
            L1_3_L2_0_G2_MINI_ALU_BoothP_15)) ;
    nor02ii ix677 (.Y (L1FirstOperands_4__15), .A0 (Instr), .A1 (
            L1_3_L2_0_G2_MINI_ALU_BoothP_16)) ;
    mux21_ni ix301 (.Y (L1FirstOperands_3__0), .A0 (
             L1_4_L2_2_G4_MINI_ALU_BoothP_1), .A1 (WindowDin_4__2__0), .S0 (
             Instr)) ;
    mux21_ni ix309 (.Y (L1FirstOperands_3__1), .A0 (
             L1_4_L2_2_G4_MINI_ALU_BoothP_2), .A1 (WindowDin_4__2__1), .S0 (
             Instr)) ;
    mux21_ni ix317 (.Y (L1FirstOperands_3__2), .A0 (
             L1_4_L2_2_G4_MINI_ALU_BoothP_3), .A1 (WindowDin_4__2__2), .S0 (
             Instr)) ;
    mux21_ni ix325 (.Y (L1FirstOperands_3__3), .A0 (
             L1_4_L2_2_G4_MINI_ALU_BoothP_4), .A1 (WindowDin_4__2__3), .S0 (
             Instr)) ;
    mux21_ni ix333 (.Y (L1FirstOperands_3__4), .A0 (
             L1_4_L2_2_G4_MINI_ALU_BoothP_5), .A1 (WindowDin_4__2__4), .S0 (
             Instr)) ;
    mux21_ni ix341 (.Y (L1FirstOperands_3__5), .A0 (
             L1_4_L2_2_G4_MINI_ALU_BoothP_6), .A1 (WindowDin_4__2__5), .S0 (
             Instr)) ;
    mux21_ni ix349 (.Y (L1FirstOperands_3__6), .A0 (
             L1_4_L2_2_G4_MINI_ALU_BoothP_7), .A1 (WindowDin_4__2__6), .S0 (
             Instr)) ;
    mux21_ni ix357 (.Y (L1FirstOperands_3__7), .A0 (
             L1_4_L2_2_G4_MINI_ALU_BoothP_8), .A1 (WindowDin_4__2__7), .S0 (
             Instr)) ;
    nor02ii ix265 (.Y (L1FirstOperands_3__8), .A0 (Instr), .A1 (
            L1_4_L2_2_G4_MINI_ALU_BoothP_9)) ;
    nor02ii ix269 (.Y (L1FirstOperands_3__9), .A0 (Instr), .A1 (
            L1_4_L2_2_G4_MINI_ALU_BoothP_10)) ;
    nor02ii ix273 (.Y (L1FirstOperands_3__10), .A0 (Instr), .A1 (
            L1_4_L2_2_G4_MINI_ALU_BoothP_11)) ;
    nor02ii ix277 (.Y (L1FirstOperands_3__11), .A0 (Instr), .A1 (
            L1_4_L2_2_G4_MINI_ALU_BoothP_12)) ;
    nor02ii ix281 (.Y (L1FirstOperands_3__12), .A0 (Instr), .A1 (
            L1_4_L2_2_G4_MINI_ALU_BoothP_13)) ;
    nor02ii ix285 (.Y (L1FirstOperands_3__13), .A0 (Instr), .A1 (
            L1_4_L2_2_G4_MINI_ALU_BoothP_14)) ;
    nor02ii ix289 (.Y (L1FirstOperands_3__14), .A0 (Instr), .A1 (
            L1_4_L2_2_G4_MINI_ALU_BoothP_15)) ;
    nor02ii ix293 (.Y (L1FirstOperands_3__15), .A0 (Instr), .A1 (
            L1_4_L2_2_G4_MINI_ALU_BoothP_16)) ;
    mux21_ni ix781 (.Y (L1FirstOperands_2__0), .A0 (
             L1_2_L2_4_G2_MINI_ALU_BoothP_1), .A1 (WindowDin_2__4__0), .S0 (
             Instr)) ;
    mux21_ni ix789 (.Y (L1FirstOperands_2__1), .A0 (
             L1_2_L2_4_G2_MINI_ALU_BoothP_2), .A1 (WindowDin_2__4__1), .S0 (
             Instr)) ;
    mux21_ni ix797 (.Y (L1FirstOperands_2__2), .A0 (
             L1_2_L2_4_G2_MINI_ALU_BoothP_3), .A1 (WindowDin_2__4__2), .S0 (
             Instr)) ;
    mux21_ni ix805 (.Y (L1FirstOperands_2__3), .A0 (
             L1_2_L2_4_G2_MINI_ALU_BoothP_4), .A1 (WindowDin_2__4__3), .S0 (
             Instr)) ;
    mux21_ni ix813 (.Y (L1FirstOperands_2__4), .A0 (
             L1_2_L2_4_G2_MINI_ALU_BoothP_5), .A1 (WindowDin_2__4__4), .S0 (
             Instr)) ;
    mux21_ni ix821 (.Y (L1FirstOperands_2__5), .A0 (
             L1_2_L2_4_G2_MINI_ALU_BoothP_6), .A1 (WindowDin_2__4__5), .S0 (
             Instr)) ;
    mux21_ni ix829 (.Y (L1FirstOperands_2__6), .A0 (
             L1_2_L2_4_G2_MINI_ALU_BoothP_7), .A1 (WindowDin_2__4__6), .S0 (
             Instr)) ;
    mux21_ni ix837 (.Y (L1FirstOperands_2__7), .A0 (
             L1_2_L2_4_G2_MINI_ALU_BoothP_8), .A1 (WindowDin_2__4__7), .S0 (
             Instr)) ;
    nor02ii ix745 (.Y (L1FirstOperands_2__8), .A0 (Instr), .A1 (
            L1_2_L2_4_G2_MINI_ALU_BoothP_9)) ;
    nor02ii ix749 (.Y (L1FirstOperands_2__9), .A0 (Instr), .A1 (
            L1_2_L2_4_G2_MINI_ALU_BoothP_10)) ;
    nor02ii ix753 (.Y (L1FirstOperands_2__10), .A0 (Instr), .A1 (
            L1_2_L2_4_G2_MINI_ALU_BoothP_11)) ;
    nor02ii ix757 (.Y (L1FirstOperands_2__11), .A0 (Instr), .A1 (
            L1_2_L2_4_G2_MINI_ALU_BoothP_12)) ;
    nor02ii ix761 (.Y (L1FirstOperands_2__12), .A0 (Instr), .A1 (
            L1_2_L2_4_G2_MINI_ALU_BoothP_13)) ;
    nor02ii ix765 (.Y (L1FirstOperands_2__13), .A0 (Instr), .A1 (
            L1_2_L2_4_G2_MINI_ALU_BoothP_14)) ;
    nor02ii ix769 (.Y (L1FirstOperands_2__14), .A0 (Instr), .A1 (
            L1_2_L2_4_G2_MINI_ALU_BoothP_15)) ;
    nor02ii ix773 (.Y (L1FirstOperands_2__15), .A0 (Instr), .A1 (
            L1_2_L2_4_G2_MINI_ALU_BoothP_16)) ;
    mux21_ni ix877 (.Y (L1FirstOperands_0__0), .A0 (
             L1_2_L2_3_G2_MINI_ALU_BoothP_1), .A1 (WindowDin_2__3__0), .S0 (
             Instr)) ;
    mux21_ni ix885 (.Y (L1FirstOperands_0__1), .A0 (
             L1_2_L2_3_G2_MINI_ALU_BoothP_2), .A1 (WindowDin_2__3__1), .S0 (
             Instr)) ;
    mux21_ni ix893 (.Y (L1FirstOperands_0__2), .A0 (
             L1_2_L2_3_G2_MINI_ALU_BoothP_3), .A1 (WindowDin_2__3__2), .S0 (
             Instr)) ;
    mux21_ni ix901 (.Y (L1FirstOperands_0__3), .A0 (
             L1_2_L2_3_G2_MINI_ALU_BoothP_4), .A1 (WindowDin_2__3__3), .S0 (
             Instr)) ;
    mux21_ni ix909 (.Y (L1FirstOperands_0__4), .A0 (
             L1_2_L2_3_G2_MINI_ALU_BoothP_5), .A1 (WindowDin_2__3__4), .S0 (
             Instr)) ;
    mux21_ni ix917 (.Y (L1FirstOperands_0__5), .A0 (
             L1_2_L2_3_G2_MINI_ALU_BoothP_6), .A1 (WindowDin_2__3__5), .S0 (
             Instr)) ;
    mux21_ni ix925 (.Y (L1FirstOperands_0__6), .A0 (
             L1_2_L2_3_G2_MINI_ALU_BoothP_7), .A1 (WindowDin_2__3__6), .S0 (
             Instr)) ;
    mux21_ni ix933 (.Y (L1FirstOperands_0__7), .A0 (
             L1_2_L2_3_G2_MINI_ALU_BoothP_8), .A1 (WindowDin_2__3__7), .S0 (
             Instr)) ;
    nor02ii ix841 (.Y (L1FirstOperands_0__8), .A0 (Instr), .A1 (
            L1_2_L2_3_G2_MINI_ALU_BoothP_9)) ;
    nor02ii ix845 (.Y (L1FirstOperands_0__9), .A0 (Instr), .A1 (
            L1_2_L2_3_G2_MINI_ALU_BoothP_10)) ;
    nor02ii ix849 (.Y (L1FirstOperands_0__10), .A0 (Instr), .A1 (
            L1_2_L2_3_G2_MINI_ALU_BoothP_11)) ;
    nor02ii ix853 (.Y (L1FirstOperands_0__11), .A0 (Instr), .A1 (
            L1_2_L2_3_G2_MINI_ALU_BoothP_12)) ;
    nor02ii ix857 (.Y (L1FirstOperands_0__12), .A0 (Instr), .A1 (
            L1_2_L2_3_G2_MINI_ALU_BoothP_13)) ;
    nor02ii ix861 (.Y (L1FirstOperands_0__13), .A0 (Instr), .A1 (
            L1_2_L2_3_G2_MINI_ALU_BoothP_14)) ;
    nor02ii ix865 (.Y (L1FirstOperands_0__14), .A0 (Instr), .A1 (
            L1_2_L2_3_G2_MINI_ALU_BoothP_15)) ;
    nor02ii ix869 (.Y (L1FirstOperands_0__15), .A0 (Instr), .A1 (
            L1_2_L2_3_G2_MINI_ALU_BoothP_16)) ;
    nor02ii ix2243 (.Y (LoopingAndResultNotReady), .A0 (nx3230), .A1 (nx2853)) ;
    nor04 ix3231 (.Y (nx3230), .A0 (CounterOut_0), .A1 (CounterOut_1), .A2 (
          CounterOut_2), .A3 (CounterOut_3)) ;
    oai21 ix29 (.Y (Result[0]), .A0 (nx3233), .A1 (Instr), .B0 (nx3235)) ;
    inv01 ix3234 (.Y (nx3233), .A (L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_0)) ;
    aoi32 ix3236 (.Y (nx3235), .A0 (L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_5), .A1 (
          FilterSize), .A2 (Instr), .B0 (
          L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_3), .B1 (nx22)) ;
    nor02ii ix23 (.Y (nx22), .A0 (FilterSize), .A1 (Instr)) ;
    oai21 ix41 (.Y (Result[1]), .A0 (nx3239), .A1 (Instr), .B0 (nx3241)) ;
    inv01 ix3240 (.Y (nx3239), .A (L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_1)) ;
    aoi32 ix3242 (.Y (nx3241), .A0 (L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_6), .A1 (
          FilterSize), .A2 (Instr), .B0 (
          L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_4), .B1 (nx22)) ;
    oai21 ix53 (.Y (Result[2]), .A0 (nx3244), .A1 (Instr), .B0 (nx3246)) ;
    inv01 ix3245 (.Y (nx3244), .A (L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_2)) ;
    aoi32 ix3247 (.Y (nx3246), .A0 (L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_7), .A1 (
          FilterSize), .A2 (Instr), .B0 (
          L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_5), .B1 (nx22)) ;
    nor02ii ix3 (.Y (Result[5]), .A0 (Instr), .A1 (
            L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_5)) ;
    nor02ii ix7 (.Y (Result[6]), .A0 (Instr), .A1 (
            L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_6)) ;
    nor02ii ix11 (.Y (Result[7]), .A0 (Instr), .A1 (
            L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_7)) ;
    inv01 ix1079 (.Y (Done), .A (NOT__145383)) ;
    inv01 ix3269 (.Y (nx3270), .A (LoopingAndResultNotReady)) ;
    inv01 ix3271 (.Y (nx3272), .A (nx3270)) ;
    inv01 ix3273 (.Y (nx3274), .A (nx3270)) ;
    inv01 ix3275 (.Y (nx3276), .A (nx3270)) ;
    inv01 ix3277 (.Y (nx3278), .A (nx3270)) ;
    inv01 ix3279 (.Y (nx3280), .A (Done)) ;
    inv01 ix3281 (.Y (nx3282), .A (Done)) ;
    inv01 ix3283 (.Y (nx3284), .A (Done)) ;
    inv01 ix3285 (.Y (nx3286), .A (Done)) ;
    and02 ix1033 (.Y (nx1032), .A0 (NOT__145383), .A1 (CLK)) ;
    or02 ix2870 (.Y (nx2869), .A0 (nx2873), .A1 (NOT_CounterOut_0)) ;
    xnor2 ix1047 (.Y (nx1046), .A0 (nx2873), .A1 (CounterOut_0)) ;
    ao22 ix61 (.Y (Result[3]), .A0 (L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_6), .A1 (
         nx22), .B0 (L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_3), .B1 (nx3292)) ;
    inv01 ix3291 (.Y (nx3292), .A (Instr)) ;
    ao22 ix69 (.Y (Result[4]), .A0 (L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_7), .A1 (
         nx22), .B0 (L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_4), .B1 (nx3292)) ;
endmodule


module booth_adder_17_unfolded14 ( AdderFirstOperand, AdderSecondOperand, 
                                   BoothOperand, BoothP, SelOperand, Operation, 
                                   AdderResult, AdderBoothResult ) ;

    input [16:0]AdderFirstOperand ;
    input [16:0]AdderSecondOperand ;
    input [16:0]BoothOperand ;
    input [16:0]BoothP ;
    input SelOperand ;
    input Operation ;
    output [16:0]AdderResult ;
    output [16:0]AdderBoothResult ;

    wire AdderResult_16_rename, AdderResult_15_rename, AdderResult_14_rename, 
         AdderResult_13_rename, AdderResult_12_rename, AdderResult_11_rename, 
         AdderResult_10_rename, AdderResult_9_rename, AdderResult_8_rename, 
         FirstOperand_16, FirstOperand_15, FirstOperand_14, FirstOperand_13, 
         FirstOperand_12, FirstOperand_11, FirstOperand_10, FirstOperand_9, 
         FirstOperand_8, FirstOperand_7, FirstOperand_6, FirstOperand_5, 
         FirstOperand_4, FirstOperand_3, FirstOperand_2, FirstOperand_1, 
         FirstOperand_0, SecondOperand_16, SecondOperand_15, SecondOperand_14, 
         SecondOperand_13, SecondOperand_12, SecondOperand_11, SecondOperand_10, 
         SecondOperand_9, SecondOperand_8, SecondOperand_7, SecondOperand_6, 
         SecondOperand_5, SecondOperand_4, SecondOperand_3, SecondOperand_2, 
         SecondOperand_1, SecondOperand_0, nx224, nx227, nx229, nx231, nx233, 
         nx235, nx237, nx239, nx241, nx243;
    wire [0:0] \$dummy ;




    assign AdderResult[16] = AdderBoothResult[16] ;
    assign AdderResult[15] = AdderBoothResult[16] ;
    assign AdderResult[14] = AdderBoothResult[16] ;
    assign AdderResult[13] = AdderBoothResult[16] ;
    assign AdderResult[12] = AdderBoothResult[16] ;
    assign AdderResult[11] = AdderBoothResult[16] ;
    assign AdderResult[10] = AdderBoothResult[16] ;
    assign AdderResult[9] = AdderBoothResult[16] ;
    assign AdderResult[8] = AdderBoothResult[16] ;
    adder_17 ADDER (.A ({FirstOperand_16,FirstOperand_15,FirstOperand_14,
             FirstOperand_13,FirstOperand_12,FirstOperand_11,FirstOperand_10,
             FirstOperand_9,FirstOperand_8,FirstOperand_7,FirstOperand_6,
             FirstOperand_5,FirstOperand_4,FirstOperand_3,FirstOperand_2,
             FirstOperand_1,FirstOperand_0}), .B ({SecondOperand_16,
             SecondOperand_15,SecondOperand_14,SecondOperand_13,SecondOperand_12
             ,SecondOperand_11,SecondOperand_10,SecondOperand_9,SecondOperand_8,
             SecondOperand_7,SecondOperand_6,SecondOperand_5,SecondOperand_4,
             SecondOperand_3,SecondOperand_2,SecondOperand_1,SecondOperand_0}), 
             .Cin (AdderBoothResult[16]), .Sum ({AdderResult_16_rename,
             AdderResult_15_rename,AdderResult_14_rename,AdderResult_13_rename,
             AdderResult_12_rename,AdderResult_11_rename,AdderResult_10_rename,
             AdderResult_9_rename,AdderResult_8_rename,AdderResult[7],
             AdderResult[6],AdderResult[5],AdderResult[4],AdderResult[3],
             AdderResult[2],AdderResult[1],AdderResult[0]}), .Cout (\$dummy [0])
             ) ;
    fake_gnd ix47 (.Y (AdderBoothResult[16])) ;
    mux21_ni ix137 (.Y (SecondOperand_0), .A0 (AdderSecondOperand[0]), .A1 (
             BoothP[0]), .S0 (nx235)) ;
    mux21_ni ix145 (.Y (SecondOperand_1), .A0 (AdderSecondOperand[1]), .A1 (
             BoothP[1]), .S0 (nx235)) ;
    mux21_ni ix153 (.Y (SecondOperand_2), .A0 (AdderSecondOperand[2]), .A1 (
             BoothP[2]), .S0 (nx235)) ;
    mux21_ni ix161 (.Y (SecondOperand_3), .A0 (AdderSecondOperand[3]), .A1 (
             BoothP[3]), .S0 (nx235)) ;
    mux21_ni ix169 (.Y (SecondOperand_4), .A0 (AdderSecondOperand[4]), .A1 (
             BoothP[4]), .S0 (nx235)) ;
    mux21_ni ix177 (.Y (SecondOperand_5), .A0 (AdderSecondOperand[5]), .A1 (
             BoothP[5]), .S0 (nx235)) ;
    mux21_ni ix185 (.Y (SecondOperand_6), .A0 (AdderSecondOperand[6]), .A1 (
             BoothP[6]), .S0 (nx235)) ;
    mux21_ni ix193 (.Y (SecondOperand_7), .A0 (AdderSecondOperand[7]), .A1 (
             BoothP[7]), .S0 (nx237)) ;
    mux21_ni ix201 (.Y (SecondOperand_8), .A0 (AdderSecondOperand[8]), .A1 (
             BoothP[8]), .S0 (nx237)) ;
    mux21_ni ix209 (.Y (SecondOperand_9), .A0 (AdderSecondOperand[9]), .A1 (
             BoothP[9]), .S0 (nx237)) ;
    mux21_ni ix217 (.Y (SecondOperand_10), .A0 (AdderSecondOperand[10]), .A1 (
             BoothP[10]), .S0 (nx237)) ;
    mux21_ni ix225 (.Y (SecondOperand_11), .A0 (AdderSecondOperand[11]), .A1 (
             BoothP[11]), .S0 (nx237)) ;
    mux21_ni ix233 (.Y (SecondOperand_12), .A0 (AdderSecondOperand[12]), .A1 (
             BoothP[12]), .S0 (nx237)) ;
    mux21_ni ix241 (.Y (SecondOperand_13), .A0 (AdderSecondOperand[13]), .A1 (
             BoothP[13]), .S0 (nx237)) ;
    mux21_ni ix249 (.Y (SecondOperand_14), .A0 (AdderSecondOperand[14]), .A1 (
             BoothP[14]), .S0 (nx239)) ;
    mux21_ni ix257 (.Y (SecondOperand_15), .A0 (AdderSecondOperand[15]), .A1 (
             BoothP[15]), .S0 (nx239)) ;
    nor02ii ix261 (.Y (FirstOperand_0), .A0 (nx239), .A1 (AdderFirstOperand[0])
            ) ;
    nor02ii ix265 (.Y (FirstOperand_1), .A0 (nx239), .A1 (AdderFirstOperand[1])
            ) ;
    nor02ii ix269 (.Y (FirstOperand_2), .A0 (nx239), .A1 (AdderFirstOperand[2])
            ) ;
    nor02ii ix273 (.Y (FirstOperand_3), .A0 (nx239), .A1 (AdderFirstOperand[3])
            ) ;
    nor02ii ix277 (.Y (FirstOperand_4), .A0 (nx239), .A1 (AdderFirstOperand[4])
            ) ;
    nor02ii ix281 (.Y (FirstOperand_5), .A0 (nx241), .A1 (AdderFirstOperand[5])
            ) ;
    nor02ii ix285 (.Y (FirstOperand_6), .A0 (nx241), .A1 (AdderFirstOperand[6])
            ) ;
    nor02ii ix289 (.Y (FirstOperand_7), .A0 (nx241), .A1 (AdderFirstOperand[7])
            ) ;
    nor02ii ix293 (.Y (FirstOperand_8), .A0 (nx241), .A1 (AdderFirstOperand[8])
            ) ;
    mux21_ni ix301 (.Y (FirstOperand_9), .A0 (AdderFirstOperand[9]), .A1 (
             BoothOperand[9]), .S0 (nx241)) ;
    mux21_ni ix309 (.Y (FirstOperand_10), .A0 (AdderFirstOperand[10]), .A1 (
             BoothOperand[10]), .S0 (nx241)) ;
    mux21_ni ix317 (.Y (FirstOperand_11), .A0 (AdderFirstOperand[11]), .A1 (
             BoothOperand[11]), .S0 (nx241)) ;
    mux21_ni ix325 (.Y (FirstOperand_12), .A0 (AdderFirstOperand[12]), .A1 (
             BoothOperand[12]), .S0 (nx243)) ;
    mux21_ni ix333 (.Y (FirstOperand_13), .A0 (AdderFirstOperand[13]), .A1 (
             BoothOperand[13]), .S0 (nx243)) ;
    mux21_ni ix341 (.Y (FirstOperand_14), .A0 (AdderFirstOperand[14]), .A1 (
             BoothOperand[14]), .S0 (nx243)) ;
    mux21_ni ix349 (.Y (FirstOperand_15), .A0 (AdderFirstOperand[15]), .A1 (
             BoothOperand[15]), .S0 (nx243)) ;
    mux21_ni ix357 (.Y (FirstOperand_16), .A0 (AdderFirstOperand[16]), .A1 (
             BoothOperand[16]), .S0 (nx243)) ;
    mux21_ni ix7 (.Y (AdderBoothResult[0]), .A0 (BoothP[1]), .A1 (AdderResult[1]
             ), .S0 (nx227)) ;
    mux21_ni ix15 (.Y (AdderBoothResult[1]), .A0 (BoothP[2]), .A1 (
             AdderResult[2]), .S0 (nx227)) ;
    mux21_ni ix23 (.Y (AdderBoothResult[2]), .A0 (BoothP[3]), .A1 (
             AdderResult[3]), .S0 (nx227)) ;
    mux21_ni ix31 (.Y (AdderBoothResult[3]), .A0 (BoothP[4]), .A1 (
             AdderResult[4]), .S0 (nx227)) ;
    mux21_ni ix39 (.Y (AdderBoothResult[4]), .A0 (BoothP[5]), .A1 (
             AdderResult[5]), .S0 (nx227)) ;
    mux21_ni ix49 (.Y (AdderBoothResult[5]), .A0 (BoothP[6]), .A1 (
             AdderResult[6]), .S0 (nx227)) ;
    mux21_ni ix55 (.Y (AdderBoothResult[6]), .A0 (BoothP[7]), .A1 (
             AdderResult[7]), .S0 (nx227)) ;
    mux21_ni ix63 (.Y (AdderBoothResult[7]), .A0 (BoothP[8]), .A1 (
             AdderResult_8_rename), .S0 (nx229)) ;
    mux21_ni ix71 (.Y (AdderBoothResult[8]), .A0 (BoothP[9]), .A1 (
             AdderResult_9_rename), .S0 (nx229)) ;
    mux21_ni ix79 (.Y (AdderBoothResult[9]), .A0 (BoothP[10]), .A1 (
             AdderResult_10_rename), .S0 (nx229)) ;
    mux21_ni ix87 (.Y (AdderBoothResult[10]), .A0 (BoothP[11]), .A1 (
             AdderResult_11_rename), .S0 (nx229)) ;
    mux21_ni ix95 (.Y (AdderBoothResult[11]), .A0 (BoothP[12]), .A1 (
             AdderResult_12_rename), .S0 (nx229)) ;
    mux21_ni ix103 (.Y (AdderBoothResult[12]), .A0 (BoothP[13]), .A1 (
             AdderResult_13_rename), .S0 (nx229)) ;
    mux21_ni ix111 (.Y (AdderBoothResult[13]), .A0 (BoothP[14]), .A1 (
             AdderResult_14_rename), .S0 (nx229)) ;
    mux21_ni ix119 (.Y (AdderBoothResult[14]), .A0 (BoothP[15]), .A1 (
             AdderResult_15_rename), .S0 (nx231)) ;
    mux21_ni ix127 (.Y (AdderBoothResult[15]), .A0 (BoothP[16]), .A1 (
             AdderResult_16_rename), .S0 (nx231)) ;
    and02 ix129 (.Y (SecondOperand_16), .A0 (nx243), .A1 (BoothP[16])) ;
    inv01 ix223 (.Y (nx224), .A (Operation)) ;
    inv02 ix226 (.Y (nx227), .A (nx224)) ;
    inv02 ix228 (.Y (nx229), .A (nx224)) ;
    inv02 ix230 (.Y (nx231), .A (nx224)) ;
    inv01 ix232 (.Y (nx233), .A (SelOperand)) ;
    inv02 ix234 (.Y (nx235), .A (nx233)) ;
    inv02 ix236 (.Y (nx237), .A (nx233)) ;
    inv02 ix238 (.Y (nx239), .A (nx233)) ;
    inv02 ix240 (.Y (nx241), .A (nx233)) ;
    inv02 ix242 (.Y (nx243), .A (nx233)) ;
endmodule


module booth_adder_17_unfolded13 ( AdderFirstOperand, AdderSecondOperand, 
                                   BoothOperand, BoothP, SelOperand, Operation, 
                                   AdderResult, AdderBoothResult ) ;

    input [16:0]AdderFirstOperand ;
    input [16:0]AdderSecondOperand ;
    input [16:0]BoothOperand ;
    input [16:0]BoothP ;
    input SelOperand ;
    input Operation ;
    output [16:0]AdderResult ;
    output [16:0]AdderBoothResult ;

    wire FirstOperand_16, FirstOperand_15, FirstOperand_14, FirstOperand_13, 
         FirstOperand_12, FirstOperand_11, FirstOperand_10, FirstOperand_9, 
         FirstOperand_8, FirstOperand_7, FirstOperand_6, FirstOperand_5, 
         FirstOperand_4, FirstOperand_3, FirstOperand_2, FirstOperand_1, 
         FirstOperand_0, SecondOperand_16, SecondOperand_15, SecondOperand_14, 
         SecondOperand_13, SecondOperand_12, SecondOperand_11, SecondOperand_10, 
         SecondOperand_9, SecondOperand_8, SecondOperand_7, SecondOperand_6, 
         SecondOperand_5, SecondOperand_4, SecondOperand_3, SecondOperand_2, 
         SecondOperand_1, SecondOperand_0, nx220, nx222, nx225, nx227, nx229, 
         nx231, nx233, nx235, nx237, nx239;
    wire [0:0] \$dummy ;




    adder_17 ADDER (.A ({FirstOperand_16,FirstOperand_15,FirstOperand_14,
             FirstOperand_13,FirstOperand_12,FirstOperand_11,FirstOperand_10,
             FirstOperand_9,FirstOperand_8,FirstOperand_7,FirstOperand_6,
             FirstOperand_5,FirstOperand_4,FirstOperand_3,FirstOperand_2,
             FirstOperand_1,FirstOperand_0}), .B ({SecondOperand_16,
             SecondOperand_15,SecondOperand_14,SecondOperand_13,SecondOperand_12
             ,SecondOperand_11,SecondOperand_10,SecondOperand_9,SecondOperand_8,
             SecondOperand_7,SecondOperand_6,SecondOperand_5,SecondOperand_4,
             SecondOperand_3,SecondOperand_2,SecondOperand_1,SecondOperand_0}), 
             .Cin (AdderBoothResult[16]), .Sum ({AdderResult[16],AdderResult[15]
             ,AdderResult[14],AdderResult[13],AdderResult[12],AdderResult[11],
             AdderResult[10],AdderResult[9],AdderResult[8],AdderResult[7],
             AdderResult[6],AdderResult[5],AdderResult[4],AdderResult[3],
             AdderResult[2],AdderResult[1],AdderResult[0]}), .Cout (\$dummy [0])
             ) ;
    fake_gnd ix45 (.Y (AdderBoothResult[16])) ;
    mux21_ni ix135 (.Y (SecondOperand_0), .A0 (AdderSecondOperand[0]), .A1 (
             BoothP[0]), .S0 (nx231)) ;
    mux21_ni ix143 (.Y (SecondOperand_1), .A0 (AdderSecondOperand[1]), .A1 (
             BoothP[1]), .S0 (nx231)) ;
    mux21_ni ix151 (.Y (SecondOperand_2), .A0 (AdderSecondOperand[2]), .A1 (
             BoothP[2]), .S0 (nx231)) ;
    mux21_ni ix159 (.Y (SecondOperand_3), .A0 (AdderSecondOperand[3]), .A1 (
             BoothP[3]), .S0 (nx231)) ;
    mux21_ni ix167 (.Y (SecondOperand_4), .A0 (AdderSecondOperand[4]), .A1 (
             BoothP[4]), .S0 (nx231)) ;
    mux21_ni ix175 (.Y (SecondOperand_5), .A0 (AdderSecondOperand[5]), .A1 (
             BoothP[5]), .S0 (nx231)) ;
    mux21_ni ix183 (.Y (SecondOperand_6), .A0 (AdderSecondOperand[6]), .A1 (
             BoothP[6]), .S0 (nx231)) ;
    mux21_ni ix191 (.Y (SecondOperand_7), .A0 (AdderSecondOperand[7]), .A1 (
             BoothP[7]), .S0 (nx233)) ;
    mux21_ni ix199 (.Y (SecondOperand_8), .A0 (AdderSecondOperand[8]), .A1 (
             BoothP[8]), .S0 (nx233)) ;
    mux21_ni ix207 (.Y (SecondOperand_9), .A0 (AdderSecondOperand[9]), .A1 (
             BoothP[9]), .S0 (nx233)) ;
    mux21_ni ix215 (.Y (SecondOperand_10), .A0 (AdderSecondOperand[10]), .A1 (
             BoothP[10]), .S0 (nx233)) ;
    mux21_ni ix223 (.Y (SecondOperand_11), .A0 (AdderSecondOperand[11]), .A1 (
             BoothP[11]), .S0 (nx233)) ;
    mux21_ni ix231 (.Y (SecondOperand_12), .A0 (AdderSecondOperand[12]), .A1 (
             BoothP[12]), .S0 (nx233)) ;
    mux21_ni ix239 (.Y (SecondOperand_13), .A0 (AdderSecondOperand[13]), .A1 (
             BoothP[13]), .S0 (nx233)) ;
    mux21_ni ix247 (.Y (SecondOperand_14), .A0 (AdderSecondOperand[14]), .A1 (
             BoothP[14]), .S0 (nx235)) ;
    mux21_ni ix255 (.Y (SecondOperand_15), .A0 (AdderSecondOperand[15]), .A1 (
             BoothP[15]), .S0 (nx235)) ;
    mux21_ni ix263 (.Y (SecondOperand_16), .A0 (AdderSecondOperand[16]), .A1 (
             BoothP[16]), .S0 (nx235)) ;
    nor02ii ix267 (.Y (FirstOperand_0), .A0 (nx235), .A1 (AdderFirstOperand[0])
            ) ;
    nor02ii ix271 (.Y (FirstOperand_1), .A0 (nx235), .A1 (AdderFirstOperand[1])
            ) ;
    nor02ii ix275 (.Y (FirstOperand_2), .A0 (nx235), .A1 (AdderFirstOperand[2])
            ) ;
    nor02ii ix279 (.Y (FirstOperand_3), .A0 (nx235), .A1 (AdderFirstOperand[3])
            ) ;
    nor02ii ix283 (.Y (FirstOperand_4), .A0 (nx237), .A1 (AdderFirstOperand[4])
            ) ;
    nor02ii ix287 (.Y (FirstOperand_5), .A0 (nx237), .A1 (AdderFirstOperand[5])
            ) ;
    nor02ii ix291 (.Y (FirstOperand_6), .A0 (nx237), .A1 (AdderFirstOperand[6])
            ) ;
    nor02ii ix295 (.Y (FirstOperand_7), .A0 (nx237), .A1 (AdderFirstOperand[7])
            ) ;
    nor02ii ix299 (.Y (FirstOperand_8), .A0 (nx237), .A1 (AdderFirstOperand[8])
            ) ;
    mux21_ni ix307 (.Y (FirstOperand_9), .A0 (AdderFirstOperand[9]), .A1 (
             BoothOperand[9]), .S0 (nx237)) ;
    mux21_ni ix315 (.Y (FirstOperand_10), .A0 (AdderFirstOperand[10]), .A1 (
             BoothOperand[10]), .S0 (nx237)) ;
    mux21_ni ix323 (.Y (FirstOperand_11), .A0 (AdderFirstOperand[11]), .A1 (
             BoothOperand[11]), .S0 (nx239)) ;
    mux21_ni ix331 (.Y (FirstOperand_12), .A0 (AdderFirstOperand[12]), .A1 (
             BoothOperand[12]), .S0 (nx239)) ;
    mux21_ni ix339 (.Y (FirstOperand_13), .A0 (AdderFirstOperand[13]), .A1 (
             BoothOperand[13]), .S0 (nx239)) ;
    mux21_ni ix347 (.Y (FirstOperand_14), .A0 (AdderFirstOperand[14]), .A1 (
             BoothOperand[14]), .S0 (nx239)) ;
    mux21_ni ix355 (.Y (FirstOperand_15), .A0 (AdderFirstOperand[15]), .A1 (
             BoothOperand[15]), .S0 (nx239)) ;
    mux21_ni ix363 (.Y (FirstOperand_16), .A0 (AdderFirstOperand[16]), .A1 (
             BoothOperand[16]), .S0 (nx239)) ;
    mux21_ni ix7 (.Y (AdderBoothResult[0]), .A0 (BoothP[1]), .A1 (AdderResult[1]
             ), .S0 (nx222)) ;
    mux21_ni ix15 (.Y (AdderBoothResult[1]), .A0 (BoothP[2]), .A1 (
             AdderResult[2]), .S0 (nx222)) ;
    mux21_ni ix23 (.Y (AdderBoothResult[2]), .A0 (BoothP[3]), .A1 (
             AdderResult[3]), .S0 (nx222)) ;
    mux21_ni ix31 (.Y (AdderBoothResult[3]), .A0 (BoothP[4]), .A1 (
             AdderResult[4]), .S0 (nx222)) ;
    mux21_ni ix39 (.Y (AdderBoothResult[4]), .A0 (BoothP[5]), .A1 (
             AdderResult[5]), .S0 (nx222)) ;
    mux21_ni ix48 (.Y (AdderBoothResult[5]), .A0 (BoothP[6]), .A1 (
             AdderResult[6]), .S0 (nx222)) ;
    mux21_ni ix55 (.Y (AdderBoothResult[6]), .A0 (BoothP[7]), .A1 (
             AdderResult[7]), .S0 (nx222)) ;
    mux21_ni ix63 (.Y (AdderBoothResult[7]), .A0 (BoothP[8]), .A1 (
             AdderResult[8]), .S0 (nx225)) ;
    mux21_ni ix71 (.Y (AdderBoothResult[8]), .A0 (BoothP[9]), .A1 (
             AdderResult[9]), .S0 (nx225)) ;
    mux21_ni ix79 (.Y (AdderBoothResult[9]), .A0 (BoothP[10]), .A1 (
             AdderResult[10]), .S0 (nx225)) ;
    mux21_ni ix87 (.Y (AdderBoothResult[10]), .A0 (BoothP[11]), .A1 (
             AdderResult[11]), .S0 (nx225)) ;
    mux21_ni ix95 (.Y (AdderBoothResult[11]), .A0 (BoothP[12]), .A1 (
             AdderResult[12]), .S0 (nx225)) ;
    mux21_ni ix103 (.Y (AdderBoothResult[12]), .A0 (BoothP[13]), .A1 (
             AdderResult[13]), .S0 (nx225)) ;
    mux21_ni ix111 (.Y (AdderBoothResult[13]), .A0 (BoothP[14]), .A1 (
             AdderResult[14]), .S0 (nx225)) ;
    mux21_ni ix119 (.Y (AdderBoothResult[14]), .A0 (BoothP[15]), .A1 (
             AdderResult[15]), .S0 (nx227)) ;
    mux21_ni ix127 (.Y (AdderBoothResult[15]), .A0 (BoothP[16]), .A1 (
             AdderResult[16]), .S0 (nx227)) ;
    inv01 ix219 (.Y (nx220), .A (Operation)) ;
    inv02 ix221 (.Y (nx222), .A (nx220)) ;
    inv02 ix224 (.Y (nx225), .A (nx220)) ;
    inv02 ix226 (.Y (nx227), .A (nx220)) ;
    inv01 ix228 (.Y (nx229), .A (SelOperand)) ;
    inv02 ix230 (.Y (nx231), .A (nx229)) ;
    inv02 ix232 (.Y (nx233), .A (nx229)) ;
    inv02 ix234 (.Y (nx235), .A (nx229)) ;
    inv02 ix236 (.Y (nx237), .A (nx229)) ;
    inv02 ix238 (.Y (nx239), .A (nx229)) ;
endmodule


module booth_unit_17_unfolded4 ( CLK, RST, Start, Instr, 
                                 LoopingAndResultNotReady, Filter, Window, 
                                 AdderBoothResult, BoothXORCheck, BoothResult, 
                                 BoothAddingOperand, BoothP, LargeWindowShifted
                                  ) ;

    input CLK ;
    input RST ;
    input Start ;
    input Instr ;
    input LoopingAndResultNotReady ;
    input [7:0]Filter ;
    input [7:0]Window ;
    input [16:0]AdderBoothResult ;
    output BoothXORCheck ;
    output [7:0]BoothResult ;
    output [16:0]BoothAddingOperand ;
    output [16:0]BoothP ;
    output [16:0]LargeWindowShifted ;

    wire BoothP_0_rename, RegisterPEN, RegisterPDin_16, RegisterPDin_15, 
         RegisterPDin_14, RegisterPDin_13, RegisterPDin_12, RegisterPDin_11, 
         RegisterPDin_10, RegisterPDin_9, RegisterPDin_8, RegisterPDin_7, 
         RegisterPDin_6, RegisterPDin_5, RegisterPDin_4, RegisterPDin_3, 
         RegisterPDin_2, RegisterPDin_1, RegisterPDin_0, RegisterSDout_10, nx12, 
         nx20, RegisterADout_10, RegisterSDout_11, nx52, nx60, RegisterADout_11, 
         RegisterSDout_12, nx92, nx100, RegisterADout_12, RegisterSDout_13, 
         nx132, nx140, RegisterADout_13, RegisterSDout_14, nx172, nx180, 
         RegisterADout_14, RegisterSDout_15, nx212, nx220, RegisterADout_15, 
         RegisterSDout_16, nx246, RegisterADout_16, nx69, nx79, nx89, nx99, 
         nx109, nx119, nx129, nx139, nx149, nx159, nx169, nx179, nx189, nx199, 
         nx209, nx224, nx226, nx235, nx249, nx261, nx273, nx286, nx299, nx315, 
         nx324, nx326, nx328;
    wire [14:0] \$dummy ;




    assign BoothResult[7] = LargeWindowShifted[16] ;
    assign BoothResult[6] = LargeWindowShifted[16] ;
    assign BoothResult[5] = LargeWindowShifted[16] ;
    assign BoothResult[4] = LargeWindowShifted[16] ;
    assign BoothResult[3] = LargeWindowShifted[16] ;
    assign BoothResult[2] = LargeWindowShifted[16] ;
    assign BoothResult[1] = LargeWindowShifted[16] ;
    assign BoothResult[0] = LargeWindowShifted[16] ;
    assign BoothAddingOperand[8] = LargeWindowShifted[16] ;
    assign BoothAddingOperand[7] = LargeWindowShifted[16] ;
    assign BoothAddingOperand[6] = LargeWindowShifted[16] ;
    assign BoothAddingOperand[5] = LargeWindowShifted[16] ;
    assign BoothAddingOperand[4] = LargeWindowShifted[16] ;
    assign BoothAddingOperand[3] = LargeWindowShifted[16] ;
    assign BoothAddingOperand[2] = LargeWindowShifted[16] ;
    assign BoothAddingOperand[1] = LargeWindowShifted[16] ;
    assign BoothAddingOperand[0] = LargeWindowShifted[16] ;
    assign BoothP[0] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[15] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[14] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[13] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[12] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[11] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[10] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[9] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[8] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[7] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[6] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[5] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[4] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[3] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[2] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[1] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[0] = LargeWindowShifted[16] ;
    register_edge_17 REGISTER_P (.CLK (CLK), .RST (RST), .EN (RegisterPEN), .Din (
                     {RegisterPDin_16,RegisterPDin_15,RegisterPDin_14,
                     RegisterPDin_13,RegisterPDin_12,RegisterPDin_11,
                     RegisterPDin_10,RegisterPDin_9,RegisterPDin_8,
                     RegisterPDin_7,RegisterPDin_6,RegisterPDin_5,RegisterPDin_4
                     ,RegisterPDin_3,RegisterPDin_2,RegisterPDin_1,
                     RegisterPDin_0}), .Dout ({BoothP[16],BoothP[15],BoothP[14],
                     BoothP[13],BoothP[12],BoothP[11],BoothP[10],BoothP[9],
                     BoothP[8],BoothP[7],BoothP[6],BoothP[5],BoothP[4],BoothP[3]
                     ,BoothP[2],BoothP[1],BoothP_0_rename})) ;
    mux_4x1_17 P_INPUT_DATA_MUX (.A ({LargeWindowShifted[16],
               AdderBoothResult[15],AdderBoothResult[14],AdderBoothResult[13],
               AdderBoothResult[12],AdderBoothResult[11],AdderBoothResult[10],
               AdderBoothResult[9],AdderBoothResult[8],AdderBoothResult[7],
               AdderBoothResult[6],AdderBoothResult[5],AdderBoothResult[4],
               AdderBoothResult[3],AdderBoothResult[2],AdderBoothResult[1],
               AdderBoothResult[0]}), .B ({LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16]}), .C ({
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],Window[7],Window[6]
               ,Window[5],Window[4],Window[3],Window[2],Window[1],Window[0],
               LargeWindowShifted[16]}), .D ({LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16]}), .S ({Start,Instr
               }), .Dout ({RegisterPDin_16,RegisterPDin_15,RegisterPDin_14,
               RegisterPDin_13,RegisterPDin_12,RegisterPDin_11,RegisterPDin_10,
               RegisterPDin_9,RegisterPDin_8,RegisterPDin_7,RegisterPDin_6,
               RegisterPDin_5,RegisterPDin_4,RegisterPDin_3,RegisterPDin_2,
               RegisterPDin_1,RegisterPDin_0})) ;
    fake_gnd ix43 (.Y (LargeWindowShifted[16])) ;
    dff REGISTER_A_reg_Dout_9 (.Q (BoothAddingOperand[9]), .QB (\$dummy [0]), .D (
        nx209), .CLK (CLK)) ;
    ao32 ix210 (.Y (nx209), .A0 (nx324), .A1 (Filter[0]), .A2 (Start), .B0 (
         BoothAddingOperand[9]), .B1 (nx326)) ;
    inv01 ix225 (.Y (nx224), .A (RST)) ;
    nor02_2x ix227 (.Y (nx226), .A0 (Start), .A1 (RST)) ;
    or02 ix287 (.Y (RegisterPEN), .A0 (Start), .A1 (LoopingAndResultNotReady)) ;
    dff REGISTER_S_reg_Dout_10 (.Q (RegisterSDout_10), .QB (\$dummy [1]), .D (
        nx69), .CLK (CLK)) ;
    mux21_ni ix70 (.Y (nx69), .A0 (nx20), .A1 (RegisterSDout_10), .S0 (nx326)) ;
    aoi21 ix21 (.Y (nx20), .A0 (Filter[1]), .A1 (Filter[0]), .B0 (nx235)) ;
    or02 ix236 (.Y (nx235), .A0 (RST), .A1 (nx12)) ;
    nor02_2x ix13 (.Y (nx12), .A0 (Filter[0]), .A1 (Filter[1])) ;
    dff REGISTER_A_reg_Dout_10 (.Q (RegisterADout_10), .QB (\$dummy [2]), .D (
        nx79), .CLK (CLK)) ;
    ao32 ix80 (.Y (nx79), .A0 (nx324), .A1 (Filter[1]), .A2 (Start), .B0 (
         RegisterADout_10), .B1 (nx326)) ;
    dff REGISTER_S_reg_Dout_11 (.Q (RegisterSDout_11), .QB (\$dummy [3]), .D (
        nx89), .CLK (CLK)) ;
    mux21_ni ix90 (.Y (nx89), .A0 (nx60), .A1 (RegisterSDout_11), .S0 (nx326)) ;
    nor03_2x ix61 (.Y (nx60), .A0 (nx249), .A1 (RST), .A2 (nx52)) ;
    nor02ii ix250 (.Y (nx249), .A0 (nx12), .A1 (Filter[2])) ;
    nor03_2x ix53 (.Y (nx52), .A0 (Filter[2]), .A1 (Filter[0]), .A2 (Filter[1])
             ) ;
    dff REGISTER_A_reg_Dout_11 (.Q (RegisterADout_11), .QB (\$dummy [4]), .D (
        nx99), .CLK (CLK)) ;
    ao32 ix100 (.Y (nx99), .A0 (nx324), .A1 (Filter[2]), .A2 (Start), .B0 (
         RegisterADout_11), .B1 (nx326)) ;
    dff REGISTER_S_reg_Dout_12 (.Q (RegisterSDout_12), .QB (\$dummy [5]), .D (
        nx109), .CLK (CLK)) ;
    mux21_ni ix110 (.Y (nx109), .A0 (nx100), .A1 (RegisterSDout_12), .S0 (nx326)
             ) ;
    nor03_2x ix101 (.Y (nx100), .A0 (nx261), .A1 (RST), .A2 (nx92)) ;
    nor02ii ix262 (.Y (nx261), .A0 (nx52), .A1 (Filter[3])) ;
    nor04 ix93 (.Y (nx92), .A0 (Filter[3]), .A1 (Filter[2]), .A2 (Filter[0]), .A3 (
          Filter[1])) ;
    dff REGISTER_A_reg_Dout_12 (.Q (RegisterADout_12), .QB (\$dummy [6]), .D (
        nx119), .CLK (CLK)) ;
    ao32 ix120 (.Y (nx119), .A0 (nx324), .A1 (Filter[3]), .A2 (Start), .B0 (
         RegisterADout_12), .B1 (nx326)) ;
    dff REGISTER_S_reg_Dout_13 (.Q (RegisterSDout_13), .QB (\$dummy [7]), .D (
        nx129), .CLK (CLK)) ;
    mux21_ni ix130 (.Y (nx129), .A0 (nx140), .A1 (RegisterSDout_13), .S0 (nx328)
             ) ;
    nor03_2x ix141 (.Y (nx140), .A0 (nx273), .A1 (RST), .A2 (nx132)) ;
    nor02ii ix274 (.Y (nx273), .A0 (nx92), .A1 (Filter[4])) ;
    nor02ii ix133 (.Y (nx132), .A0 (Filter[4]), .A1 (nx92)) ;
    dff REGISTER_A_reg_Dout_13 (.Q (RegisterADout_13), .QB (\$dummy [8]), .D (
        nx139), .CLK (CLK)) ;
    ao32 ix140 (.Y (nx139), .A0 (nx324), .A1 (Filter[4]), .A2 (Start), .B0 (
         RegisterADout_13), .B1 (nx328)) ;
    dff REGISTER_S_reg_Dout_14 (.Q (RegisterSDout_14), .QB (\$dummy [9]), .D (
        nx149), .CLK (CLK)) ;
    mux21_ni ix150 (.Y (nx149), .A0 (nx180), .A1 (RegisterSDout_14), .S0 (nx328)
             ) ;
    nor03_2x ix181 (.Y (nx180), .A0 (nx286), .A1 (RST), .A2 (nx172)) ;
    nor02ii ix288 (.Y (nx286), .A0 (nx132), .A1 (Filter[5])) ;
    nor02ii ix173 (.Y (nx172), .A0 (Filter[5]), .A1 (nx132)) ;
    dff REGISTER_A_reg_Dout_14 (.Q (RegisterADout_14), .QB (\$dummy [10]), .D (
        nx159), .CLK (CLK)) ;
    ao32 ix160 (.Y (nx159), .A0 (nx324), .A1 (Filter[5]), .A2 (Start), .B0 (
         RegisterADout_14), .B1 (nx328)) ;
    dff REGISTER_S_reg_Dout_15 (.Q (RegisterSDout_15), .QB (\$dummy [11]), .D (
        nx169), .CLK (CLK)) ;
    mux21_ni ix170 (.Y (nx169), .A0 (nx220), .A1 (RegisterSDout_15), .S0 (nx328)
             ) ;
    nor03_2x ix221 (.Y (nx220), .A0 (nx299), .A1 (RST), .A2 (nx212)) ;
    nor02ii ix300 (.Y (nx299), .A0 (nx172), .A1 (Filter[6])) ;
    nor02ii ix213 (.Y (nx212), .A0 (Filter[6]), .A1 (nx172)) ;
    dff REGISTER_A_reg_Dout_15 (.Q (RegisterADout_15), .QB (\$dummy [12]), .D (
        nx179), .CLK (CLK)) ;
    ao32 ix180 (.Y (nx179), .A0 (nx324), .A1 (Filter[6]), .A2 (Start), .B0 (
         RegisterADout_15), .B1 (nx328)) ;
    dff REGISTER_S_reg_Dout_16 (.Q (RegisterSDout_16), .QB (\$dummy [13]), .D (
        nx189), .CLK (CLK)) ;
    ao32 ix190 (.Y (nx189), .A0 (nx224), .A1 (nx246), .A2 (Start), .B0 (
         RegisterSDout_16), .B1 (nx328)) ;
    xnor2 ix247 (.Y (nx246), .A0 (Filter[7]), .A1 (nx212)) ;
    dff REGISTER_A_reg_Dout_16 (.Q (RegisterADout_16), .QB (\$dummy [14]), .D (
        nx199), .CLK (CLK)) ;
    ao32 ix200 (.Y (nx199), .A0 (nx224), .A1 (Filter[7]), .A2 (Start), .B0 (
         RegisterADout_16), .B1 (nx226)) ;
    inv02 ix316 (.Y (nx315), .A (BoothP_0_rename)) ;
    inv01 ix323 (.Y (nx324), .A (RST)) ;
    nor02_2x ix325 (.Y (nx326), .A0 (Start), .A1 (RST)) ;
    nor02_2x ix327 (.Y (nx328), .A0 (Start), .A1 (RST)) ;
    mux21_ni ix46 (.Y (BoothAddingOperand[10]), .A0 (RegisterADout_10), .A1 (
             RegisterSDout_10), .S0 (nx315)) ;
    mux21_ni ix85 (.Y (BoothAddingOperand[11]), .A0 (RegisterADout_11), .A1 (
             RegisterSDout_11), .S0 (nx315)) ;
    mux21_ni ix125 (.Y (BoothAddingOperand[12]), .A0 (RegisterADout_12), .A1 (
             RegisterSDout_12), .S0 (nx315)) ;
    mux21_ni ix165 (.Y (BoothAddingOperand[13]), .A0 (RegisterADout_13), .A1 (
             RegisterSDout_13), .S0 (nx315)) ;
    mux21_ni ix205 (.Y (BoothAddingOperand[14]), .A0 (RegisterADout_14), .A1 (
             RegisterSDout_14), .S0 (nx315)) ;
    mux21_ni ix245 (.Y (BoothAddingOperand[15]), .A0 (RegisterADout_15), .A1 (
             RegisterSDout_15), .S0 (nx315)) ;
    mux21_ni ix275 (.Y (BoothAddingOperand[16]), .A0 (RegisterADout_16), .A1 (
             RegisterSDout_16), .S0 (nx315)) ;
    xor2 ix289 (.Y (BoothXORCheck), .A0 (BoothP[1]), .A1 (BoothP_0_rename)) ;
endmodule


module booth_adder_17_unfolded12 ( AdderFirstOperand, AdderSecondOperand, 
                                   BoothOperand, BoothP, SelOperand, Operation, 
                                   AdderResult, AdderBoothResult ) ;

    input [16:0]AdderFirstOperand ;
    input [16:0]AdderSecondOperand ;
    input [16:0]BoothOperand ;
    input [16:0]BoothP ;
    input SelOperand ;
    input Operation ;
    output [16:0]AdderResult ;
    output [16:0]AdderBoothResult ;

    wire AdderResult_16_rename, AdderResult_15_rename, AdderResult_14_rename, 
         AdderResult_13_rename, AdderResult_12_rename, AdderResult_11_rename, 
         AdderResult_10_rename, AdderResult_9_rename, FirstOperand_16, 
         FirstOperand_15, FirstOperand_14, FirstOperand_13, FirstOperand_12, 
         FirstOperand_11, FirstOperand_10, FirstOperand_9, SecondOperand_16, 
         SecondOperand_15, SecondOperand_14, SecondOperand_13, SecondOperand_12, 
         SecondOperand_11, SecondOperand_10, SecondOperand_9, SecondOperand_8, 
         SecondOperand_7, SecondOperand_6, SecondOperand_5, SecondOperand_4, 
         nx143, nx153, nx155, nx158, nx161, nx164, nx167, nx182, nx184, nx186, 
         nx188, nx190, nx192, nx194;
    wire [9:0] \$dummy ;




    assign AdderResult[16] = AdderBoothResult[16] ;
    assign AdderResult[15] = AdderBoothResult[16] ;
    assign AdderResult[14] = AdderBoothResult[16] ;
    assign AdderResult[13] = AdderBoothResult[16] ;
    assign AdderResult[12] = AdderBoothResult[16] ;
    assign AdderResult[11] = AdderBoothResult[16] ;
    assign AdderResult[10] = AdderBoothResult[16] ;
    assign AdderResult[9] = AdderBoothResult[16] ;
    assign AdderResult[8] = AdderBoothResult[16] ;
    assign AdderResult[7] = AdderBoothResult[16] ;
    assign AdderResult[6] = AdderBoothResult[16] ;
    assign AdderResult[5] = AdderBoothResult[16] ;
    assign AdderResult[4] = AdderBoothResult[16] ;
    assign AdderResult[3] = AdderBoothResult[16] ;
    assign AdderResult[2] = AdderBoothResult[16] ;
    assign AdderResult[1] = AdderBoothResult[16] ;
    assign AdderResult[0] = AdderBoothResult[16] ;
    adder_17_unfolded4 ADDER (.A ({FirstOperand_16,FirstOperand_15,
                       FirstOperand_14,FirstOperand_13,FirstOperand_12,
                       FirstOperand_11,FirstOperand_10,FirstOperand_9,
                       AdderBoothResult[16],AdderBoothResult[16],
                       AdderBoothResult[16],AdderBoothResult[16],
                       AdderBoothResult[16],AdderBoothResult[16],
                       AdderBoothResult[16],AdderBoothResult[16],
                       AdderBoothResult[16]}), .B ({SecondOperand_16,
                       SecondOperand_15,SecondOperand_14,SecondOperand_13,
                       SecondOperand_12,SecondOperand_11,SecondOperand_10,
                       SecondOperand_9,SecondOperand_8,SecondOperand_7,
                       SecondOperand_6,SecondOperand_5,SecondOperand_4,
                       AdderBoothResult[16],AdderBoothResult[16],
                       AdderBoothResult[16],AdderBoothResult[16]}), .Cin (
                       AdderBoothResult[16]), .Sum ({AdderResult_16_rename,
                       AdderResult_15_rename,AdderResult_14_rename,
                       AdderResult_13_rename,AdderResult_12_rename,
                       AdderResult_11_rename,AdderResult_10_rename,
                       AdderResult_9_rename,\$dummy [0],\$dummy [1],\$dummy [2],
                       \$dummy [3],\$dummy [4],\$dummy [5],\$dummy [6],
                       \$dummy [7],\$dummy [8]}), .Cout (\$dummy [9])) ;
    fake_gnd ix59 (.Y (AdderBoothResult[16])) ;
    and02 ix15 (.Y (SecondOperand_4), .A0 (BoothP[4]), .A1 (nx186)) ;
    and02 ix25 (.Y (SecondOperand_5), .A0 (BoothP[5]), .A1 (nx186)) ;
    and02 ix35 (.Y (SecondOperand_6), .A0 (BoothP[6]), .A1 (nx186)) ;
    and02 ix45 (.Y (SecondOperand_7), .A0 (BoothP[7]), .A1 (nx186)) ;
    and02 ix55 (.Y (SecondOperand_8), .A0 (BoothP[8]), .A1 (nx186)) ;
    and02 ix125 (.Y (SecondOperand_9), .A0 (BoothP[9]), .A1 (nx186)) ;
    and02 ix127 (.Y (SecondOperand_10), .A0 (BoothP[10]), .A1 (nx186)) ;
    and02 ix129 (.Y (SecondOperand_11), .A0 (BoothP[11]), .A1 (nx188)) ;
    and02 ix131 (.Y (SecondOperand_12), .A0 (BoothP[12]), .A1 (nx188)) ;
    and02 ix133 (.Y (SecondOperand_13), .A0 (BoothP[13]), .A1 (nx188)) ;
    and02 ix135 (.Y (SecondOperand_14), .A0 (BoothP[14]), .A1 (nx188)) ;
    and02 ix137 (.Y (SecondOperand_15), .A0 (BoothP[15]), .A1 (nx188)) ;
    and02 ix139 (.Y (SecondOperand_16), .A0 (BoothP[16]), .A1 (nx188)) ;
    and02 ix141 (.Y (FirstOperand_9), .A0 (BoothOperand[9]), .A1 (nx188)) ;
    and02 ix143 (.Y (FirstOperand_10), .A0 (BoothOperand[10]), .A1 (nx190)) ;
    and02 ix145 (.Y (FirstOperand_11), .A0 (BoothOperand[11]), .A1 (nx190)) ;
    and02 ix147 (.Y (FirstOperand_12), .A0 (BoothOperand[12]), .A1 (nx190)) ;
    and02 ix149 (.Y (FirstOperand_13), .A0 (BoothOperand[13]), .A1 (nx190)) ;
    and02 ix151 (.Y (FirstOperand_14), .A0 (BoothOperand[14]), .A1 (nx190)) ;
    and02 ix153 (.Y (FirstOperand_15), .A0 (BoothOperand[15]), .A1 (nx190)) ;
    and02 ix155 (.Y (FirstOperand_16), .A0 (nx190), .A1 (BoothOperand[16])) ;
    nor02ii ix5 (.Y (AdderBoothResult[0]), .A0 (nx143), .A1 (BoothP[1])) ;
    nor02ii ix7 (.Y (AdderBoothResult[1]), .A0 (nx143), .A1 (BoothP[2])) ;
    nor02ii ix9 (.Y (AdderBoothResult[2]), .A0 (nx143), .A1 (BoothP[3])) ;
    aoi21 ix19 (.Y (AdderBoothResult[3]), .A0 (nx182), .A1 (nx194), .B0 (nx155)
          ) ;
    inv01 ix154 (.Y (nx153), .A (SelOperand)) ;
    inv01 ix156 (.Y (nx155), .A (BoothP[4])) ;
    aoi21 ix29 (.Y (AdderBoothResult[4]), .A0 (nx182), .A1 (nx194), .B0 (nx158)
          ) ;
    inv01 ix159 (.Y (nx158), .A (BoothP[5])) ;
    aoi21 ix39 (.Y (AdderBoothResult[5]), .A0 (nx182), .A1 (nx194), .B0 (nx161)
          ) ;
    inv01 ix162 (.Y (nx161), .A (BoothP[6])) ;
    aoi21 ix49 (.Y (AdderBoothResult[6]), .A0 (nx182), .A1 (nx194), .B0 (nx164)
          ) ;
    inv01 ix165 (.Y (nx164), .A (BoothP[7])) ;
    aoi21 ix61 (.Y (AdderBoothResult[7]), .A0 (nx182), .A1 (nx194), .B0 (nx167)
          ) ;
    inv01 ix168 (.Y (nx167), .A (BoothP[8])) ;
    mux21_ni ix67 (.Y (AdderBoothResult[8]), .A0 (BoothP[9]), .A1 (
             AdderResult_9_rename), .S0 (nx182)) ;
    mux21_ni ix75 (.Y (AdderBoothResult[9]), .A0 (BoothP[10]), .A1 (
             AdderResult_10_rename), .S0 (nx182)) ;
    mux21_ni ix83 (.Y (AdderBoothResult[10]), .A0 (BoothP[11]), .A1 (
             AdderResult_11_rename), .S0 (nx184)) ;
    mux21_ni ix91 (.Y (AdderBoothResult[11]), .A0 (BoothP[12]), .A1 (
             AdderResult_12_rename), .S0 (nx184)) ;
    mux21_ni ix99 (.Y (AdderBoothResult[12]), .A0 (BoothP[13]), .A1 (
             AdderResult_13_rename), .S0 (nx184)) ;
    mux21_ni ix107 (.Y (AdderBoothResult[13]), .A0 (BoothP[14]), .A1 (
             AdderResult_14_rename), .S0 (nx184)) ;
    mux21_ni ix115 (.Y (AdderBoothResult[14]), .A0 (BoothP[15]), .A1 (
             AdderResult_15_rename), .S0 (nx184)) ;
    mux21_ni ix123 (.Y (AdderBoothResult[15]), .A0 (BoothP[16]), .A1 (
             AdderResult_16_rename), .S0 (nx184)) ;
    nor02ii ix144 (.Y (nx143), .A0 (nx192), .A1 (nx184)) ;
    buf02 ix181 (.Y (nx182), .A (Operation)) ;
    buf02 ix183 (.Y (nx184), .A (Operation)) ;
    inv02 ix185 (.Y (nx186), .A (nx194)) ;
    inv02 ix187 (.Y (nx188), .A (nx153)) ;
    inv02 ix189 (.Y (nx190), .A (nx153)) ;
    inv02 ix191 (.Y (nx192), .A (nx153)) ;
    inv01 ix193 (.Y (nx194), .A (SelOperand)) ;
endmodule


module adder_17_unfolded4 ( A, B, Cin, Sum, Cout ) ;

    input [16:0]A ;
    input [16:0]B ;
    input Cin ;
    output [16:0]Sum ;
    output Cout ;

    wire nx2, nx16, nx18, nx32, nx34, nx48, nx93, nx95, nx98, nx101, nx105, 
         nx107, nx110, nx113, nx117, nx119, nx122, nx125, nx129, nx131;



    assign Sum[8] = B[8] ;
    assign Sum[7] = B[7] ;
    assign Sum[6] = B[6] ;
    assign Sum[5] = B[5] ;
    assign Sum[4] = B[4] ;
    assign Sum[3] = Cout ;
    assign Sum[2] = Cout ;
    assign Sum[1] = Cout ;
    assign Sum[0] = Cout ;
    fake_gnd ix68 (.Y (Cout)) ;
    xor2 ix71 (.Y (Sum[9]), .A0 (B[9]), .A1 (A[9])) ;
    xor2 ix65 (.Y (Sum[10]), .A0 (nx93), .A1 (nx95)) ;
    nand02 ix94 (.Y (nx93), .A0 (B[9]), .A1 (A[9])) ;
    xnor2 ix96 (.Y (nx95), .A0 (A[10]), .A1 (B[10])) ;
    xor2 ix63 (.Y (Sum[11]), .A0 (nx98), .A1 (nx101)) ;
    aoi32 ix99 (.Y (nx98), .A0 (B[9]), .A1 (A[9]), .A2 (nx2), .B0 (B[10]), .B1 (
          A[10])) ;
    xnor2 ix102 (.Y (nx101), .A0 (A[11]), .A1 (B[11])) ;
    xnor2 ix61 (.Y (Sum[12]), .A0 (nx16), .A1 (nx107)) ;
    oai21 ix17 (.Y (nx16), .A0 (nx98), .A1 (nx101), .B0 (nx105)) ;
    nand02 ix106 (.Y (nx105), .A0 (B[11]), .A1 (A[11])) ;
    xnor2 ix108 (.Y (nx107), .A0 (A[12]), .A1 (B[12])) ;
    xor2 ix59 (.Y (Sum[13]), .A0 (nx110), .A1 (nx113)) ;
    aoi22 ix111 (.Y (nx110), .A0 (B[12]), .A1 (A[12]), .B0 (nx16), .B1 (nx18)) ;
    xnor2 ix114 (.Y (nx113), .A0 (A[13]), .A1 (B[13])) ;
    xnor2 ix57 (.Y (Sum[14]), .A0 (nx32), .A1 (nx119)) ;
    oai21 ix33 (.Y (nx32), .A0 (nx110), .A1 (nx113), .B0 (nx117)) ;
    nand02 ix118 (.Y (nx117), .A0 (B[13]), .A1 (A[13])) ;
    xnor2 ix120 (.Y (nx119), .A0 (A[14]), .A1 (B[14])) ;
    xor2 ix55 (.Y (Sum[15]), .A0 (nx122), .A1 (nx125)) ;
    aoi22 ix123 (.Y (nx122), .A0 (B[14]), .A1 (A[14]), .B0 (nx32), .B1 (nx34)) ;
    xnor2 ix126 (.Y (nx125), .A0 (A[15]), .A1 (B[15])) ;
    xnor2 ix53 (.Y (Sum[16]), .A0 (nx48), .A1 (nx131)) ;
    oai21 ix49 (.Y (nx48), .A0 (nx122), .A1 (nx125), .B0 (nx129)) ;
    nand02 ix130 (.Y (nx129), .A0 (B[15]), .A1 (A[15])) ;
    xnor2 ix132 (.Y (nx131), .A0 (A[16]), .A1 (B[16])) ;
    inv01 ix35 (.Y (nx34), .A (nx119)) ;
    inv01 ix19 (.Y (nx18), .A (nx107)) ;
    inv01 ix3 (.Y (nx2), .A (nx95)) ;
endmodule


module booth_unit_17 ( CLK, RST, Start, Instr, LoopingAndResultNotReady, Filter, 
                       Window, AdderBoothResult, BoothXORCheck, BoothResult, 
                       BoothAddingOperand, BoothP, LargeWindowShifted ) ;

    input CLK ;
    input RST ;
    input Start ;
    input Instr ;
    input LoopingAndResultNotReady ;
    input [7:0]Filter ;
    input [7:0]Window ;
    input [16:0]AdderBoothResult ;
    output BoothXORCheck ;
    output [7:0]BoothResult ;
    output [16:0]BoothAddingOperand ;
    output [16:0]BoothP ;
    output [16:0]LargeWindowShifted ;

    wire RegisterPEN, RegisterPDin_16, RegisterPDin_15, RegisterPDin_14, 
         RegisterPDin_13, RegisterPDin_12, RegisterPDin_11, RegisterPDin_10, 
         RegisterPDin_9, RegisterPDin_8, RegisterPDin_7, RegisterPDin_6, 
         RegisterPDin_5, RegisterPDin_4, RegisterPDin_3, RegisterPDin_2, 
         RegisterPDin_1, RegisterPDin_0, RegisterSDout_10, nx12, nx20, 
         RegisterADout_10, RegisterSDout_11, nx52, nx60, RegisterADout_11, 
         RegisterSDout_12, nx92, nx100, RegisterADout_12, RegisterSDout_13, 
         nx132, nx140, RegisterADout_13, RegisterSDout_14, nx172, nx180, 
         RegisterADout_14, RegisterSDout_15, nx212, nx220, RegisterADout_15, 
         RegisterSDout_16, nx246, RegisterADout_16, nx69, nx79, nx89, nx99, 
         nx109, nx119, nx129, nx139, nx149, nx159, nx169, nx179, nx189, nx199, 
         nx209, nx224, nx226, nx235, nx249, nx261, nx273, nx286, nx299, nx320, 
         nx322, nx324, nx326, nx328;
    wire [14:0] \$dummy ;




    assign BoothResult[7] = LargeWindowShifted[16] ;
    assign BoothResult[6] = LargeWindowShifted[16] ;
    assign BoothResult[5] = LargeWindowShifted[16] ;
    assign BoothResult[4] = LargeWindowShifted[16] ;
    assign BoothResult[3] = LargeWindowShifted[16] ;
    assign BoothResult[2] = LargeWindowShifted[16] ;
    assign BoothResult[1] = LargeWindowShifted[16] ;
    assign BoothResult[0] = LargeWindowShifted[16] ;
    assign BoothAddingOperand[8] = LargeWindowShifted[16] ;
    assign BoothAddingOperand[7] = LargeWindowShifted[16] ;
    assign BoothAddingOperand[6] = LargeWindowShifted[16] ;
    assign BoothAddingOperand[5] = LargeWindowShifted[16] ;
    assign BoothAddingOperand[4] = LargeWindowShifted[16] ;
    assign BoothAddingOperand[3] = LargeWindowShifted[16] ;
    assign BoothAddingOperand[2] = LargeWindowShifted[16] ;
    assign BoothAddingOperand[1] = LargeWindowShifted[16] ;
    assign BoothAddingOperand[0] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[15] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[14] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[13] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[12] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[11] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[10] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[9] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[8] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[7] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[6] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[5] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[4] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[3] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[2] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[1] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[0] = LargeWindowShifted[16] ;
    register_edge_17 REGISTER_P (.CLK (CLK), .RST (RST), .EN (RegisterPEN), .Din (
                     {RegisterPDin_16,RegisterPDin_15,RegisterPDin_14,
                     RegisterPDin_13,RegisterPDin_12,RegisterPDin_11,
                     RegisterPDin_10,RegisterPDin_9,RegisterPDin_8,
                     RegisterPDin_7,RegisterPDin_6,RegisterPDin_5,RegisterPDin_4
                     ,RegisterPDin_3,RegisterPDin_2,RegisterPDin_1,
                     RegisterPDin_0}), .Dout ({BoothP[16],BoothP[15],BoothP[14],
                     BoothP[13],BoothP[12],BoothP[11],BoothP[10],BoothP[9],
                     BoothP[8],BoothP[7],BoothP[6],BoothP[5],BoothP[4],BoothP[3]
                     ,BoothP[2],BoothP[1],BoothP[0]})) ;
    mux_4x1_17 P_INPUT_DATA_MUX (.A ({LargeWindowShifted[16],
               AdderBoothResult[15],AdderBoothResult[14],AdderBoothResult[13],
               AdderBoothResult[12],AdderBoothResult[11],AdderBoothResult[10],
               AdderBoothResult[9],AdderBoothResult[8],AdderBoothResult[7],
               AdderBoothResult[6],AdderBoothResult[5],AdderBoothResult[4],
               AdderBoothResult[3],AdderBoothResult[2],AdderBoothResult[1],
               AdderBoothResult[0]}), .B ({LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16]}), .C ({
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],Window[7],Window[6]
               ,Window[5],Window[4],Window[3],Window[2],Window[1],Window[0],
               LargeWindowShifted[16]}), .D ({LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16]}), .S ({Start,Instr
               }), .Dout ({RegisterPDin_16,RegisterPDin_15,RegisterPDin_14,
               RegisterPDin_13,RegisterPDin_12,RegisterPDin_11,RegisterPDin_10,
               RegisterPDin_9,RegisterPDin_8,RegisterPDin_7,RegisterPDin_6,
               RegisterPDin_5,RegisterPDin_4,RegisterPDin_3,RegisterPDin_2,
               RegisterPDin_1,RegisterPDin_0})) ;
    fake_gnd ix43 (.Y (LargeWindowShifted[16])) ;
    dff REGISTER_A_reg_Dout_9 (.Q (BoothAddingOperand[9]), .QB (\$dummy [0]), .D (
        nx209), .CLK (CLK)) ;
    ao32 ix210 (.Y (nx209), .A0 (nx324), .A1 (Filter[0]), .A2 (Start), .B0 (
         BoothAddingOperand[9]), .B1 (nx326)) ;
    inv01 ix225 (.Y (nx224), .A (RST)) ;
    nor02_2x ix227 (.Y (nx226), .A0 (Start), .A1 (RST)) ;
    or02 ix287 (.Y (RegisterPEN), .A0 (Start), .A1 (LoopingAndResultNotReady)) ;
    mux21_ni ix46 (.Y (BoothAddingOperand[10]), .A0 (RegisterSDout_10), .A1 (
             RegisterADout_10), .S0 (nx320)) ;
    dff REGISTER_S_reg_Dout_10 (.Q (RegisterSDout_10), .QB (\$dummy [1]), .D (
        nx69), .CLK (CLK)) ;
    mux21_ni ix70 (.Y (nx69), .A0 (nx20), .A1 (RegisterSDout_10), .S0 (nx326)) ;
    aoi21 ix21 (.Y (nx20), .A0 (Filter[1]), .A1 (Filter[0]), .B0 (nx235)) ;
    or02 ix236 (.Y (nx235), .A0 (RST), .A1 (nx12)) ;
    nor02_2x ix13 (.Y (nx12), .A0 (Filter[0]), .A1 (Filter[1])) ;
    dff REGISTER_A_reg_Dout_10 (.Q (RegisterADout_10), .QB (\$dummy [2]), .D (
        nx79), .CLK (CLK)) ;
    ao32 ix80 (.Y (nx79), .A0 (nx324), .A1 (Filter[1]), .A2 (Start), .B0 (
         RegisterADout_10), .B1 (nx326)) ;
    mux21_ni ix85 (.Y (BoothAddingOperand[11]), .A0 (RegisterSDout_11), .A1 (
             RegisterADout_11), .S0 (nx320)) ;
    dff REGISTER_S_reg_Dout_11 (.Q (RegisterSDout_11), .QB (\$dummy [3]), .D (
        nx89), .CLK (CLK)) ;
    mux21_ni ix90 (.Y (nx89), .A0 (nx60), .A1 (RegisterSDout_11), .S0 (nx326)) ;
    nor03_2x ix61 (.Y (nx60), .A0 (nx249), .A1 (RST), .A2 (nx52)) ;
    nor02ii ix250 (.Y (nx249), .A0 (nx12), .A1 (Filter[2])) ;
    nor03_2x ix53 (.Y (nx52), .A0 (Filter[2]), .A1 (Filter[0]), .A2 (Filter[1])
             ) ;
    dff REGISTER_A_reg_Dout_11 (.Q (RegisterADout_11), .QB (\$dummy [4]), .D (
        nx99), .CLK (CLK)) ;
    ao32 ix100 (.Y (nx99), .A0 (nx324), .A1 (Filter[2]), .A2 (Start), .B0 (
         RegisterADout_11), .B1 (nx326)) ;
    mux21_ni ix125 (.Y (BoothAddingOperand[12]), .A0 (RegisterSDout_12), .A1 (
             RegisterADout_12), .S0 (nx320)) ;
    dff REGISTER_S_reg_Dout_12 (.Q (RegisterSDout_12), .QB (\$dummy [5]), .D (
        nx109), .CLK (CLK)) ;
    mux21_ni ix110 (.Y (nx109), .A0 (nx100), .A1 (RegisterSDout_12), .S0 (nx326)
             ) ;
    nor03_2x ix101 (.Y (nx100), .A0 (nx261), .A1 (RST), .A2 (nx92)) ;
    nor02ii ix262 (.Y (nx261), .A0 (nx52), .A1 (Filter[3])) ;
    nor04 ix93 (.Y (nx92), .A0 (Filter[3]), .A1 (Filter[2]), .A2 (Filter[0]), .A3 (
          Filter[1])) ;
    dff REGISTER_A_reg_Dout_12 (.Q (RegisterADout_12), .QB (\$dummy [6]), .D (
        nx119), .CLK (CLK)) ;
    ao32 ix120 (.Y (nx119), .A0 (nx324), .A1 (Filter[3]), .A2 (Start), .B0 (
         RegisterADout_12), .B1 (nx326)) ;
    mux21_ni ix165 (.Y (BoothAddingOperand[13]), .A0 (RegisterSDout_13), .A1 (
             RegisterADout_13), .S0 (nx320)) ;
    dff REGISTER_S_reg_Dout_13 (.Q (RegisterSDout_13), .QB (\$dummy [7]), .D (
        nx129), .CLK (CLK)) ;
    mux21_ni ix130 (.Y (nx129), .A0 (nx140), .A1 (RegisterSDout_13), .S0 (nx328)
             ) ;
    nor03_2x ix141 (.Y (nx140), .A0 (nx273), .A1 (RST), .A2 (nx132)) ;
    nor02ii ix274 (.Y (nx273), .A0 (nx92), .A1 (Filter[4])) ;
    nor02ii ix133 (.Y (nx132), .A0 (Filter[4]), .A1 (nx92)) ;
    dff REGISTER_A_reg_Dout_13 (.Q (RegisterADout_13), .QB (\$dummy [8]), .D (
        nx139), .CLK (CLK)) ;
    ao32 ix140 (.Y (nx139), .A0 (nx324), .A1 (Filter[4]), .A2 (Start), .B0 (
         RegisterADout_13), .B1 (nx328)) ;
    mux21_ni ix205 (.Y (BoothAddingOperand[14]), .A0 (RegisterSDout_14), .A1 (
             RegisterADout_14), .S0 (nx320)) ;
    dff REGISTER_S_reg_Dout_14 (.Q (RegisterSDout_14), .QB (\$dummy [9]), .D (
        nx149), .CLK (CLK)) ;
    mux21_ni ix150 (.Y (nx149), .A0 (nx180), .A1 (RegisterSDout_14), .S0 (nx328)
             ) ;
    nor03_2x ix181 (.Y (nx180), .A0 (nx286), .A1 (RST), .A2 (nx172)) ;
    nor02ii ix288 (.Y (nx286), .A0 (nx132), .A1 (Filter[5])) ;
    nor02ii ix173 (.Y (nx172), .A0 (Filter[5]), .A1 (nx132)) ;
    dff REGISTER_A_reg_Dout_14 (.Q (RegisterADout_14), .QB (\$dummy [10]), .D (
        nx159), .CLK (CLK)) ;
    ao32 ix160 (.Y (nx159), .A0 (nx324), .A1 (Filter[5]), .A2 (Start), .B0 (
         RegisterADout_14), .B1 (nx328)) ;
    mux21_ni ix245 (.Y (BoothAddingOperand[15]), .A0 (RegisterSDout_15), .A1 (
             RegisterADout_15), .S0 (nx320)) ;
    dff REGISTER_S_reg_Dout_15 (.Q (RegisterSDout_15), .QB (\$dummy [11]), .D (
        nx169), .CLK (CLK)) ;
    mux21_ni ix170 (.Y (nx169), .A0 (nx220), .A1 (RegisterSDout_15), .S0 (nx328)
             ) ;
    nor03_2x ix221 (.Y (nx220), .A0 (nx299), .A1 (RST), .A2 (nx212)) ;
    nor02ii ix300 (.Y (nx299), .A0 (nx172), .A1 (Filter[6])) ;
    nor02ii ix213 (.Y (nx212), .A0 (Filter[6]), .A1 (nx172)) ;
    dff REGISTER_A_reg_Dout_15 (.Q (RegisterADout_15), .QB (\$dummy [12]), .D (
        nx179), .CLK (CLK)) ;
    ao32 ix180 (.Y (nx179), .A0 (nx324), .A1 (Filter[6]), .A2 (Start), .B0 (
         RegisterADout_15), .B1 (nx328)) ;
    mux21_ni ix275 (.Y (BoothAddingOperand[16]), .A0 (RegisterSDout_16), .A1 (
             RegisterADout_16), .S0 (nx320)) ;
    dff REGISTER_S_reg_Dout_16 (.Q (RegisterSDout_16), .QB (\$dummy [13]), .D (
        nx189), .CLK (CLK)) ;
    ao32 ix190 (.Y (nx189), .A0 (nx224), .A1 (nx246), .A2 (Start), .B0 (
         RegisterSDout_16), .B1 (nx328)) ;
    xnor2 ix247 (.Y (nx246), .A0 (Filter[7]), .A1 (nx212)) ;
    dff REGISTER_A_reg_Dout_16 (.Q (RegisterADout_16), .QB (\$dummy [14]), .D (
        nx199), .CLK (CLK)) ;
    ao32 ix200 (.Y (nx199), .A0 (nx224), .A1 (Filter[7]), .A2 (Start), .B0 (
         RegisterADout_16), .B1 (nx226)) ;
    xor2 ix289 (.Y (BoothXORCheck), .A0 (BoothP[1]), .A1 (nx322)) ;
    buf02 ix319 (.Y (nx320), .A (BoothP[0])) ;
    buf02 ix321 (.Y (nx322), .A (BoothP[0])) ;
    inv01 ix323 (.Y (nx324), .A (RST)) ;
    nor02_2x ix325 (.Y (nx326), .A0 (Start), .A1 (RST)) ;
    nor02_2x ix327 (.Y (nx328), .A0 (Start), .A1 (RST)) ;
endmodule


module mux_4x1_17 ( A, B, C, D, S, Dout ) ;

    input [16:0]A ;
    input [16:0]B ;
    input [16:0]C ;
    input [16:0]D ;
    input [1:0]S ;
    output [16:0]Dout ;

    wire nx28, nx46, nx131, nx136, nx139, nx142, nx145, nx148, nx151, nx166, 
         nx168, nx170, nx172, nx178, nx180;



    fake_gnd ix85 (.Y (Dout[16])) ;
    ao22 ix37 (.Y (Dout[0]), .A0 (A[0]), .A1 (nx170), .B0 (C[1]), .B1 (nx166)) ;
    and02 ix29 (.Y (nx28), .A0 (S[0]), .A1 (S[1])) ;
    inv01 ix53 (.Y (Dout[1]), .A (nx131)) ;
    aoi222 ix132 (.Y (nx131), .A0 (A[1]), .A1 (nx170), .B0 (C[1]), .B1 (nx178), 
           .C0 (C[2]), .C1 (nx166)) ;
    inv01 ix65 (.Y (Dout[2]), .A (nx136)) ;
    aoi222 ix137 (.Y (nx136), .A0 (A[2]), .A1 (nx170), .B0 (C[2]), .B1 (nx178), 
           .C0 (C[3]), .C1 (nx166)) ;
    inv01 ix77 (.Y (Dout[3]), .A (nx139)) ;
    aoi222 ix140 (.Y (nx139), .A0 (A[3]), .A1 (nx170), .B0 (C[3]), .B1 (nx178), 
           .C0 (C[4]), .C1 (nx166)) ;
    inv01 ix89 (.Y (Dout[4]), .A (nx142)) ;
    aoi222 ix143 (.Y (nx142), .A0 (A[4]), .A1 (nx170), .B0 (C[4]), .B1 (nx178), 
           .C0 (C[5]), .C1 (nx166)) ;
    inv01 ix101 (.Y (Dout[5]), .A (nx145)) ;
    aoi222 ix146 (.Y (nx145), .A0 (A[5]), .A1 (nx170), .B0 (C[5]), .B1 (nx178), 
           .C0 (C[6]), .C1 (nx166)) ;
    inv01 ix113 (.Y (Dout[6]), .A (nx148)) ;
    aoi222 ix149 (.Y (nx148), .A0 (A[6]), .A1 (nx172), .B0 (C[6]), .B1 (nx178), 
           .C0 (C[7]), .C1 (nx166)) ;
    inv01 ix125 (.Y (Dout[7]), .A (nx151)) ;
    aoi222 ix152 (.Y (nx151), .A0 (A[7]), .A1 (nx172), .B0 (C[7]), .B1 (nx178), 
           .C0 (C[8]), .C1 (nx168)) ;
    ao22 ix133 (.Y (Dout[8]), .A0 (nx172), .A1 (A[8]), .B0 (C[8]), .B1 (nx180)
         ) ;
    nor02ii ix3 (.Y (Dout[9]), .A0 (S[1]), .A1 (A[9])) ;
    nor02ii ix7 (.Y (Dout[10]), .A0 (S[1]), .A1 (A[10])) ;
    nor02ii ix11 (.Y (Dout[11]), .A0 (S[1]), .A1 (A[11])) ;
    nor02ii ix15 (.Y (Dout[12]), .A0 (S[1]), .A1 (A[12])) ;
    nor02ii ix19 (.Y (Dout[13]), .A0 (S[1]), .A1 (A[13])) ;
    nor02ii ix23 (.Y (Dout[14]), .A0 (S[1]), .A1 (A[14])) ;
    nor02ii ix27 (.Y (Dout[15]), .A0 (S[1]), .A1 (A[15])) ;
    buf02 ix165 (.Y (nx166), .A (nx28)) ;
    buf02 ix167 (.Y (nx168), .A (nx28)) ;
    inv02 ix169 (.Y (nx170), .A (S[1])) ;
    inv02 ix171 (.Y (nx172), .A (S[1])) ;
    nor02ii ix47 (.Y (nx46), .A0 (S[0]), .A1 (S[1])) ;
    buf02 ix177 (.Y (nx178), .A (nx46)) ;
    buf02 ix179 (.Y (nx180), .A (nx46)) ;
endmodule


module register_edge_17 ( CLK, RST, EN, Din, Dout ) ;

    input CLK ;
    input RST ;
    input EN ;
    input [16:0]Din ;
    output [16:0]Dout ;

    wire nx402, nx412, nx422, nx432, nx442, nx452, nx462, nx472, nx482, nx492, 
         nx502, nx512, nx522, nx532, nx542, nx552, nx562, nx574, nx576, nx632, 
         nx634, nx636, nx638, nx644, nx646, nx648, nx650;
    wire [16:0] \$dummy ;




    dff reg_Dout_0 (.Q (Dout[0]), .QB (\$dummy [0]), .D (nx402), .CLK (CLK)) ;
    ao32 ix403 (.Y (nx402), .A0 (Din[0]), .A1 (nx632), .A2 (nx646), .B0 (Dout[0]
         ), .B1 (nx636)) ;
    inv01 ix575 (.Y (nx574), .A (RST)) ;
    nor02_2x ix577 (.Y (nx576), .A0 (RST), .A1 (nx646)) ;
    dff reg_Dout_1 (.Q (Dout[1]), .QB (\$dummy [1]), .D (nx412), .CLK (CLK)) ;
    ao32 ix413 (.Y (nx412), .A0 (Din[1]), .A1 (nx632), .A2 (nx646), .B0 (Dout[1]
         ), .B1 (nx636)) ;
    dff reg_Dout_2 (.Q (Dout[2]), .QB (\$dummy [2]), .D (nx422), .CLK (CLK)) ;
    ao32 ix423 (.Y (nx422), .A0 (Din[2]), .A1 (nx632), .A2 (nx646), .B0 (Dout[2]
         ), .B1 (nx636)) ;
    dff reg_Dout_3 (.Q (Dout[3]), .QB (\$dummy [3]), .D (nx432), .CLK (CLK)) ;
    ao32 ix433 (.Y (nx432), .A0 (Din[3]), .A1 (nx632), .A2 (nx646), .B0 (Dout[3]
         ), .B1 (nx636)) ;
    dff reg_Dout_4 (.Q (Dout[4]), .QB (\$dummy [4]), .D (nx442), .CLK (CLK)) ;
    ao32 ix443 (.Y (nx442), .A0 (Din[4]), .A1 (nx632), .A2 (nx646), .B0 (Dout[4]
         ), .B1 (nx636)) ;
    dff reg_Dout_5 (.Q (Dout[5]), .QB (\$dummy [5]), .D (nx452), .CLK (CLK)) ;
    ao32 ix453 (.Y (nx452), .A0 (Din[5]), .A1 (nx632), .A2 (nx646), .B0 (Dout[5]
         ), .B1 (nx636)) ;
    dff reg_Dout_6 (.Q (Dout[6]), .QB (\$dummy [6]), .D (nx462), .CLK (CLK)) ;
    ao32 ix463 (.Y (nx462), .A0 (Din[6]), .A1 (nx634), .A2 (nx648), .B0 (Dout[6]
         ), .B1 (nx636)) ;
    dff reg_Dout_7 (.Q (Dout[7]), .QB (\$dummy [7]), .D (nx472), .CLK (CLK)) ;
    ao32 ix473 (.Y (nx472), .A0 (Din[7]), .A1 (nx634), .A2 (nx648), .B0 (Dout[7]
         ), .B1 (nx638)) ;
    dff reg_Dout_8 (.Q (Dout[8]), .QB (\$dummy [8]), .D (nx482), .CLK (CLK)) ;
    ao32 ix483 (.Y (nx482), .A0 (Din[8]), .A1 (nx634), .A2 (nx648), .B0 (Dout[8]
         ), .B1 (nx638)) ;
    dff reg_Dout_9 (.Q (Dout[9]), .QB (\$dummy [9]), .D (nx492), .CLK (CLK)) ;
    ao32 ix493 (.Y (nx492), .A0 (Din[9]), .A1 (nx634), .A2 (nx648), .B0 (Dout[9]
         ), .B1 (nx638)) ;
    dff reg_Dout_10 (.Q (Dout[10]), .QB (\$dummy [10]), .D (nx502), .CLK (CLK)
        ) ;
    ao32 ix503 (.Y (nx502), .A0 (Din[10]), .A1 (nx634), .A2 (nx648), .B0 (
         Dout[10]), .B1 (nx638)) ;
    dff reg_Dout_11 (.Q (Dout[11]), .QB (\$dummy [11]), .D (nx512), .CLK (CLK)
        ) ;
    ao32 ix513 (.Y (nx512), .A0 (Din[11]), .A1 (nx634), .A2 (nx648), .B0 (
         Dout[11]), .B1 (nx638)) ;
    dff reg_Dout_12 (.Q (Dout[12]), .QB (\$dummy [12]), .D (nx522), .CLK (CLK)
        ) ;
    ao32 ix523 (.Y (nx522), .A0 (Din[12]), .A1 (nx574), .A2 (nx648), .B0 (
         Dout[12]), .B1 (nx638)) ;
    dff reg_Dout_13 (.Q (Dout[13]), .QB (\$dummy [13]), .D (nx532), .CLK (CLK)
        ) ;
    ao32 ix533 (.Y (nx532), .A0 (Din[13]), .A1 (nx574), .A2 (nx650), .B0 (
         Dout[13]), .B1 (nx638)) ;
    dff reg_Dout_14 (.Q (Dout[14]), .QB (\$dummy [14]), .D (nx542), .CLK (CLK)
        ) ;
    ao32 ix543 (.Y (nx542), .A0 (Din[14]), .A1 (nx574), .A2 (nx650), .B0 (
         Dout[14]), .B1 (nx576)) ;
    dff reg_Dout_15 (.Q (Dout[15]), .QB (\$dummy [15]), .D (nx552), .CLK (CLK)
        ) ;
    ao32 ix553 (.Y (nx552), .A0 (Din[15]), .A1 (nx574), .A2 (nx650), .B0 (
         Dout[15]), .B1 (nx576)) ;
    dff reg_Dout_16 (.Q (Dout[16]), .QB (\$dummy [16]), .D (nx562), .CLK (CLK)
        ) ;
    ao32 ix563 (.Y (nx562), .A0 (Din[16]), .A1 (nx574), .A2 (nx650), .B0 (
         Dout[16]), .B1 (nx576)) ;
    inv01 ix631 (.Y (nx632), .A (RST)) ;
    inv01 ix633 (.Y (nx634), .A (RST)) ;
    nor02_2x ix635 (.Y (nx636), .A0 (RST), .A1 (nx650)) ;
    nor02_2x ix637 (.Y (nx638), .A0 (RST), .A1 (nx650)) ;
    inv01 ix643 (.Y (nx644), .A (EN)) ;
    inv02 ix645 (.Y (nx646), .A (nx644)) ;
    inv02 ix647 (.Y (nx648), .A (nx644)) ;
    inv02 ix649 (.Y (nx650), .A (nx644)) ;
endmodule


module booth_adder_17 ( AdderFirstOperand, AdderSecondOperand, BoothOperand, 
                        BoothP, SelOperand, Operation, AdderResult, 
                        AdderBoothResult ) ;

    input [16:0]AdderFirstOperand ;
    input [16:0]AdderSecondOperand ;
    input [16:0]BoothOperand ;
    input [16:0]BoothP ;
    input SelOperand ;
    input Operation ;
    output [16:0]AdderResult ;
    output [16:0]AdderBoothResult ;

    wire FirstOperand_16, FirstOperand_15, FirstOperand_14, FirstOperand_13, 
         FirstOperand_12, FirstOperand_11, FirstOperand_10, FirstOperand_9, 
         FirstOperand_8, FirstOperand_7, FirstOperand_6, FirstOperand_5, 
         FirstOperand_4, FirstOperand_3, FirstOperand_2, FirstOperand_1, 
         FirstOperand_0, SecondOperand_16, SecondOperand_15, SecondOperand_14, 
         SecondOperand_13, SecondOperand_12, SecondOperand_11, SecondOperand_10, 
         SecondOperand_9, SecondOperand_8, SecondOperand_7, SecondOperand_6, 
         SecondOperand_5, SecondOperand_4, SecondOperand_3, SecondOperand_2, 
         SecondOperand_1, SecondOperand_0, nx224, nx227, nx229, nx231, nx233, 
         nx235, nx237, nx239, nx241, nx243;
    wire [0:0] \$dummy ;




    adder_17 ADDER (.A ({FirstOperand_16,FirstOperand_15,FirstOperand_14,
             FirstOperand_13,FirstOperand_12,FirstOperand_11,FirstOperand_10,
             FirstOperand_9,FirstOperand_8,FirstOperand_7,FirstOperand_6,
             FirstOperand_5,FirstOperand_4,FirstOperand_3,FirstOperand_2,
             FirstOperand_1,FirstOperand_0}), .B ({SecondOperand_16,
             SecondOperand_15,SecondOperand_14,SecondOperand_13,SecondOperand_12
             ,SecondOperand_11,SecondOperand_10,SecondOperand_9,SecondOperand_8,
             SecondOperand_7,SecondOperand_6,SecondOperand_5,SecondOperand_4,
             SecondOperand_3,SecondOperand_2,SecondOperand_1,SecondOperand_0}), 
             .Cin (AdderBoothResult[16]), .Sum ({AdderResult[16],AdderResult[15]
             ,AdderResult[14],AdderResult[13],AdderResult[12],AdderResult[11],
             AdderResult[10],AdderResult[9],AdderResult[8],AdderResult[7],
             AdderResult[6],AdderResult[5],AdderResult[4],AdderResult[3],
             AdderResult[2],AdderResult[1],AdderResult[0]}), .Cout (\$dummy [0])
             ) ;
    fake_gnd ix47 (.Y (AdderBoothResult[16])) ;
    mux21_ni ix137 (.Y (SecondOperand_0), .A0 (AdderSecondOperand[0]), .A1 (
             BoothP[0]), .S0 (nx235)) ;
    mux21_ni ix145 (.Y (SecondOperand_1), .A0 (AdderSecondOperand[1]), .A1 (
             BoothP[1]), .S0 (nx235)) ;
    mux21_ni ix153 (.Y (SecondOperand_2), .A0 (AdderSecondOperand[2]), .A1 (
             BoothP[2]), .S0 (nx235)) ;
    mux21_ni ix161 (.Y (SecondOperand_3), .A0 (AdderSecondOperand[3]), .A1 (
             BoothP[3]), .S0 (nx235)) ;
    mux21_ni ix169 (.Y (SecondOperand_4), .A0 (AdderSecondOperand[4]), .A1 (
             BoothP[4]), .S0 (nx235)) ;
    mux21_ni ix177 (.Y (SecondOperand_5), .A0 (AdderSecondOperand[5]), .A1 (
             BoothP[5]), .S0 (nx235)) ;
    mux21_ni ix185 (.Y (SecondOperand_6), .A0 (AdderSecondOperand[6]), .A1 (
             BoothP[6]), .S0 (nx235)) ;
    mux21_ni ix193 (.Y (SecondOperand_7), .A0 (AdderSecondOperand[7]), .A1 (
             BoothP[7]), .S0 (nx237)) ;
    mux21_ni ix201 (.Y (SecondOperand_8), .A0 (AdderSecondOperand[8]), .A1 (
             BoothP[8]), .S0 (nx237)) ;
    mux21_ni ix209 (.Y (SecondOperand_9), .A0 (AdderSecondOperand[9]), .A1 (
             BoothP[9]), .S0 (nx237)) ;
    mux21_ni ix217 (.Y (SecondOperand_10), .A0 (AdderSecondOperand[10]), .A1 (
             BoothP[10]), .S0 (nx237)) ;
    mux21_ni ix225 (.Y (SecondOperand_11), .A0 (AdderSecondOperand[11]), .A1 (
             BoothP[11]), .S0 (nx237)) ;
    mux21_ni ix233 (.Y (SecondOperand_12), .A0 (AdderSecondOperand[12]), .A1 (
             BoothP[12]), .S0 (nx237)) ;
    mux21_ni ix241 (.Y (SecondOperand_13), .A0 (AdderSecondOperand[13]), .A1 (
             BoothP[13]), .S0 (nx237)) ;
    mux21_ni ix249 (.Y (SecondOperand_14), .A0 (AdderSecondOperand[14]), .A1 (
             BoothP[14]), .S0 (nx239)) ;
    mux21_ni ix257 (.Y (SecondOperand_15), .A0 (AdderSecondOperand[15]), .A1 (
             BoothP[15]), .S0 (nx239)) ;
    nor02ii ix261 (.Y (FirstOperand_0), .A0 (nx239), .A1 (AdderFirstOperand[0])
            ) ;
    nor02ii ix265 (.Y (FirstOperand_1), .A0 (nx239), .A1 (AdderFirstOperand[1])
            ) ;
    nor02ii ix269 (.Y (FirstOperand_2), .A0 (nx239), .A1 (AdderFirstOperand[2])
            ) ;
    nor02ii ix273 (.Y (FirstOperand_3), .A0 (nx239), .A1 (AdderFirstOperand[3])
            ) ;
    nor02ii ix277 (.Y (FirstOperand_4), .A0 (nx239), .A1 (AdderFirstOperand[4])
            ) ;
    nor02ii ix281 (.Y (FirstOperand_5), .A0 (nx241), .A1 (AdderFirstOperand[5])
            ) ;
    nor02ii ix285 (.Y (FirstOperand_6), .A0 (nx241), .A1 (AdderFirstOperand[6])
            ) ;
    nor02ii ix289 (.Y (FirstOperand_7), .A0 (nx241), .A1 (AdderFirstOperand[7])
            ) ;
    nor02ii ix293 (.Y (FirstOperand_8), .A0 (nx241), .A1 (AdderFirstOperand[8])
            ) ;
    mux21_ni ix303 (.Y (FirstOperand_9), .A0 (AdderFirstOperand[9]), .A1 (
             BoothOperand[9]), .S0 (nx241)) ;
    mux21_ni ix311 (.Y (FirstOperand_10), .A0 (AdderFirstOperand[10]), .A1 (
             BoothOperand[10]), .S0 (nx241)) ;
    mux21_ni ix319 (.Y (FirstOperand_11), .A0 (AdderFirstOperand[11]), .A1 (
             BoothOperand[11]), .S0 (nx241)) ;
    mux21_ni ix327 (.Y (FirstOperand_12), .A0 (AdderFirstOperand[12]), .A1 (
             BoothOperand[12]), .S0 (nx243)) ;
    mux21_ni ix335 (.Y (FirstOperand_13), .A0 (AdderFirstOperand[13]), .A1 (
             BoothOperand[13]), .S0 (nx243)) ;
    mux21_ni ix343 (.Y (FirstOperand_14), .A0 (AdderFirstOperand[14]), .A1 (
             BoothOperand[14]), .S0 (nx243)) ;
    mux21_ni ix351 (.Y (FirstOperand_15), .A0 (AdderFirstOperand[15]), .A1 (
             BoothOperand[15]), .S0 (nx243)) ;
    mux21_ni ix7 (.Y (AdderBoothResult[0]), .A0 (BoothP[1]), .A1 (AdderResult[1]
             ), .S0 (nx227)) ;
    mux21_ni ix15 (.Y (AdderBoothResult[1]), .A0 (BoothP[2]), .A1 (
             AdderResult[2]), .S0 (nx227)) ;
    mux21_ni ix23 (.Y (AdderBoothResult[2]), .A0 (BoothP[3]), .A1 (
             AdderResult[3]), .S0 (nx227)) ;
    mux21_ni ix31 (.Y (AdderBoothResult[3]), .A0 (BoothP[4]), .A1 (
             AdderResult[4]), .S0 (nx227)) ;
    mux21_ni ix39 (.Y (AdderBoothResult[4]), .A0 (BoothP[5]), .A1 (
             AdderResult[5]), .S0 (nx227)) ;
    mux21_ni ix49 (.Y (AdderBoothResult[5]), .A0 (BoothP[6]), .A1 (
             AdderResult[6]), .S0 (nx227)) ;
    mux21_ni ix55 (.Y (AdderBoothResult[6]), .A0 (BoothP[7]), .A1 (
             AdderResult[7]), .S0 (nx227)) ;
    mux21_ni ix63 (.Y (AdderBoothResult[7]), .A0 (BoothP[8]), .A1 (
             AdderResult[8]), .S0 (nx229)) ;
    mux21_ni ix71 (.Y (AdderBoothResult[8]), .A0 (BoothP[9]), .A1 (
             AdderResult[9]), .S0 (nx229)) ;
    mux21_ni ix79 (.Y (AdderBoothResult[9]), .A0 (BoothP[10]), .A1 (
             AdderResult[10]), .S0 (nx229)) ;
    mux21_ni ix87 (.Y (AdderBoothResult[10]), .A0 (BoothP[11]), .A1 (
             AdderResult[11]), .S0 (nx229)) ;
    mux21_ni ix95 (.Y (AdderBoothResult[11]), .A0 (BoothP[12]), .A1 (
             AdderResult[12]), .S0 (nx229)) ;
    mux21_ni ix103 (.Y (AdderBoothResult[12]), .A0 (BoothP[13]), .A1 (
             AdderResult[13]), .S0 (nx229)) ;
    mux21_ni ix111 (.Y (AdderBoothResult[13]), .A0 (BoothP[14]), .A1 (
             AdderResult[14]), .S0 (nx229)) ;
    mux21_ni ix119 (.Y (AdderBoothResult[14]), .A0 (BoothP[15]), .A1 (
             AdderResult[15]), .S0 (nx231)) ;
    mux21_ni ix127 (.Y (AdderBoothResult[15]), .A0 (BoothP[16]), .A1 (
             AdderResult[16]), .S0 (nx231)) ;
    and02 ix129 (.Y (SecondOperand_16), .A0 (nx243), .A1 (BoothP[16])) ;
    and02 ix295 (.Y (FirstOperand_16), .A0 (nx243), .A1 (BoothOperand[16])) ;
    inv01 ix223 (.Y (nx224), .A (Operation)) ;
    inv02 ix226 (.Y (nx227), .A (nx224)) ;
    inv02 ix228 (.Y (nx229), .A (nx224)) ;
    inv02 ix230 (.Y (nx231), .A (nx224)) ;
    inv01 ix232 (.Y (nx233), .A (SelOperand)) ;
    inv02 ix234 (.Y (nx235), .A (nx233)) ;
    inv02 ix236 (.Y (nx237), .A (nx233)) ;
    inv02 ix238 (.Y (nx239), .A (nx233)) ;
    inv02 ix240 (.Y (nx241), .A (nx233)) ;
    inv02 ix242 (.Y (nx243), .A (nx233)) ;
endmodule


module adder_17 ( A, B, Cin, Sum, Cout ) ;

    input [16:0]A ;
    input [16:0]B ;
    input Cin ;
    output [16:0]Sum ;
    output Cout ;

    wire nx2, nx16, nx18, nx32, nx34, nx48, nx50, nx64, nx66, nx80, nx82, nx96, 
         nx98, nx112, nx114, nx122, nx105, nx107, nx111, nx115, nx121, nx123, 
         nx127, nx131, nx137, nx139, nx143, nx147, nx153, nx155, nx159, nx163, 
         nx167, nx169, nx172, nx175, nx179, nx181, nx184, nx187, nx191, nx193, 
         nx196, nx199, nx203, nx205, nx208;



    fake_gnd ix58 (.Y (Cout)) ;
    xor2 ix161 (.Y (Sum[0]), .A0 (B[0]), .A1 (A[0])) ;
    xor2 ix155 (.Y (Sum[1]), .A0 (nx105), .A1 (nx107)) ;
    nand02 ix106 (.Y (nx105), .A0 (B[0]), .A1 (A[0])) ;
    xnor2 ix108 (.Y (nx107), .A0 (A[1]), .A1 (B[1])) ;
    xor2 ix153 (.Y (Sum[2]), .A0 (nx111), .A1 (nx115)) ;
    aoi32 ix112 (.Y (nx111), .A0 (B[0]), .A1 (A[0]), .A2 (nx2), .B0 (B[1]), .B1 (
          A[1])) ;
    xnor2 ix116 (.Y (nx115), .A0 (A[2]), .A1 (B[2])) ;
    xnor2 ix151 (.Y (Sum[3]), .A0 (nx16), .A1 (nx123)) ;
    oai21 ix17 (.Y (nx16), .A0 (nx111), .A1 (nx115), .B0 (nx121)) ;
    nand02 ix122 (.Y (nx121), .A0 (B[2]), .A1 (A[2])) ;
    xnor2 ix124 (.Y (nx123), .A0 (A[3]), .A1 (B[3])) ;
    xor2 ix149 (.Y (Sum[4]), .A0 (nx127), .A1 (nx131)) ;
    aoi22 ix128 (.Y (nx127), .A0 (B[3]), .A1 (A[3]), .B0 (nx16), .B1 (nx18)) ;
    xnor2 ix132 (.Y (nx131), .A0 (A[4]), .A1 (B[4])) ;
    xnor2 ix147 (.Y (Sum[5]), .A0 (nx32), .A1 (nx139)) ;
    oai21 ix33 (.Y (nx32), .A0 (nx127), .A1 (nx131), .B0 (nx137)) ;
    nand02 ix138 (.Y (nx137), .A0 (B[4]), .A1 (A[4])) ;
    xnor2 ix140 (.Y (nx139), .A0 (A[5]), .A1 (B[5])) ;
    xor2 ix145 (.Y (Sum[6]), .A0 (nx143), .A1 (nx147)) ;
    aoi22 ix144 (.Y (nx143), .A0 (B[5]), .A1 (A[5]), .B0 (nx32), .B1 (nx34)) ;
    xnor2 ix148 (.Y (nx147), .A0 (A[6]), .A1 (B[6])) ;
    xnor2 ix143 (.Y (Sum[7]), .A0 (nx48), .A1 (nx155)) ;
    oai21 ix49 (.Y (nx48), .A0 (nx143), .A1 (nx147), .B0 (nx153)) ;
    nand02 ix154 (.Y (nx153), .A0 (B[6]), .A1 (A[6])) ;
    xnor2 ix156 (.Y (nx155), .A0 (A[7]), .A1 (B[7])) ;
    xor2 ix141 (.Y (Sum[8]), .A0 (nx159), .A1 (nx163)) ;
    aoi22 ix160 (.Y (nx159), .A0 (B[7]), .A1 (A[7]), .B0 (nx48), .B1 (nx50)) ;
    xnor2 ix164 (.Y (nx163), .A0 (A[8]), .A1 (B[8])) ;
    xnor2 ix139 (.Y (Sum[9]), .A0 (nx64), .A1 (nx169)) ;
    oai21 ix65 (.Y (nx64), .A0 (nx159), .A1 (nx163), .B0 (nx167)) ;
    nand02 ix168 (.Y (nx167), .A0 (B[8]), .A1 (A[8])) ;
    xnor2 ix170 (.Y (nx169), .A0 (A[9]), .A1 (B[9])) ;
    xor2 ix137 (.Y (Sum[10]), .A0 (nx172), .A1 (nx175)) ;
    aoi22 ix173 (.Y (nx172), .A0 (B[9]), .A1 (A[9]), .B0 (nx64), .B1 (nx66)) ;
    xnor2 ix176 (.Y (nx175), .A0 (A[10]), .A1 (B[10])) ;
    xnor2 ix135 (.Y (Sum[11]), .A0 (nx80), .A1 (nx181)) ;
    oai21 ix81 (.Y (nx80), .A0 (nx172), .A1 (nx175), .B0 (nx179)) ;
    nand02 ix180 (.Y (nx179), .A0 (B[10]), .A1 (A[10])) ;
    xnor2 ix182 (.Y (nx181), .A0 (A[11]), .A1 (B[11])) ;
    xor2 ix133 (.Y (Sum[12]), .A0 (nx184), .A1 (nx187)) ;
    aoi22 ix185 (.Y (nx184), .A0 (B[11]), .A1 (A[11]), .B0 (nx80), .B1 (nx82)) ;
    xnor2 ix188 (.Y (nx187), .A0 (A[12]), .A1 (B[12])) ;
    xnor2 ix131 (.Y (Sum[13]), .A0 (nx96), .A1 (nx193)) ;
    oai21 ix97 (.Y (nx96), .A0 (nx184), .A1 (nx187), .B0 (nx191)) ;
    nand02 ix192 (.Y (nx191), .A0 (B[12]), .A1 (A[12])) ;
    xnor2 ix194 (.Y (nx193), .A0 (A[13]), .A1 (B[13])) ;
    xor2 ix129 (.Y (Sum[14]), .A0 (nx196), .A1 (nx199)) ;
    aoi22 ix197 (.Y (nx196), .A0 (B[13]), .A1 (A[13]), .B0 (nx96), .B1 (nx98)) ;
    xnor2 ix200 (.Y (nx199), .A0 (A[14]), .A1 (B[14])) ;
    xnor2 ix127 (.Y (Sum[15]), .A0 (nx112), .A1 (nx205)) ;
    oai21 ix113 (.Y (nx112), .A0 (nx196), .A1 (nx199), .B0 (nx203)) ;
    nand02 ix204 (.Y (nx203), .A0 (B[14]), .A1 (A[14])) ;
    xnor2 ix206 (.Y (nx205), .A0 (A[15]), .A1 (B[15])) ;
    xnor2 ix125 (.Y (Sum[16]), .A0 (nx208), .A1 (nx122)) ;
    aoi22 ix209 (.Y (nx208), .A0 (B[15]), .A1 (A[15]), .B0 (nx112), .B1 (nx114)
          ) ;
    xor2 ix123 (.Y (nx122), .A0 (A[16]), .A1 (B[16])) ;
    inv01 ix115 (.Y (nx114), .A (nx205)) ;
    inv01 ix99 (.Y (nx98), .A (nx193)) ;
    inv01 ix83 (.Y (nx82), .A (nx181)) ;
    inv01 ix67 (.Y (nx66), .A (nx169)) ;
    inv01 ix51 (.Y (nx50), .A (nx155)) ;
    inv01 ix35 (.Y (nx34), .A (nx139)) ;
    inv01 ix19 (.Y (nx18), .A (nx123)) ;
    inv01 ix3 (.Y (nx2), .A (nx107)) ;
endmodule

