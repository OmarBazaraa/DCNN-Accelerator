//
// Verilog description for cell cache, 
// Wed May  9 07:36:08 2018
//
// LeonardoSpectrum Level 3, 2017a.2 
//


module cache ( CLK, RST, FilterSize, FilterWR, WindowWR, Din, FilterDout_0__0__7, 
               FilterDout_0__0__6, FilterDout_0__0__5, FilterDout_0__0__4, 
               FilterDout_0__0__3, FilterDout_0__0__2, FilterDout_0__0__1, 
               FilterDout_0__0__0, FilterDout_0__1__7, FilterDout_0__1__6, 
               FilterDout_0__1__5, FilterDout_0__1__4, FilterDout_0__1__3, 
               FilterDout_0__1__2, FilterDout_0__1__1, FilterDout_0__1__0, 
               FilterDout_0__2__7, FilterDout_0__2__6, FilterDout_0__2__5, 
               FilterDout_0__2__4, FilterDout_0__2__3, FilterDout_0__2__2, 
               FilterDout_0__2__1, FilterDout_0__2__0, FilterDout_0__3__7, 
               FilterDout_0__3__6, FilterDout_0__3__5, FilterDout_0__3__4, 
               FilterDout_0__3__3, FilterDout_0__3__2, FilterDout_0__3__1, 
               FilterDout_0__3__0, FilterDout_0__4__7, FilterDout_0__4__6, 
               FilterDout_0__4__5, FilterDout_0__4__4, FilterDout_0__4__3, 
               FilterDout_0__4__2, FilterDout_0__4__1, FilterDout_0__4__0, 
               FilterDout_1__0__7, FilterDout_1__0__6, FilterDout_1__0__5, 
               FilterDout_1__0__4, FilterDout_1__0__3, FilterDout_1__0__2, 
               FilterDout_1__0__1, FilterDout_1__0__0, FilterDout_1__1__7, 
               FilterDout_1__1__6, FilterDout_1__1__5, FilterDout_1__1__4, 
               FilterDout_1__1__3, FilterDout_1__1__2, FilterDout_1__1__1, 
               FilterDout_1__1__0, FilterDout_1__2__7, FilterDout_1__2__6, 
               FilterDout_1__2__5, FilterDout_1__2__4, FilterDout_1__2__3, 
               FilterDout_1__2__2, FilterDout_1__2__1, FilterDout_1__2__0, 
               FilterDout_1__3__7, FilterDout_1__3__6, FilterDout_1__3__5, 
               FilterDout_1__3__4, FilterDout_1__3__3, FilterDout_1__3__2, 
               FilterDout_1__3__1, FilterDout_1__3__0, FilterDout_1__4__7, 
               FilterDout_1__4__6, FilterDout_1__4__5, FilterDout_1__4__4, 
               FilterDout_1__4__3, FilterDout_1__4__2, FilterDout_1__4__1, 
               FilterDout_1__4__0, FilterDout_2__0__7, FilterDout_2__0__6, 
               FilterDout_2__0__5, FilterDout_2__0__4, FilterDout_2__0__3, 
               FilterDout_2__0__2, FilterDout_2__0__1, FilterDout_2__0__0, 
               FilterDout_2__1__7, FilterDout_2__1__6, FilterDout_2__1__5, 
               FilterDout_2__1__4, FilterDout_2__1__3, FilterDout_2__1__2, 
               FilterDout_2__1__1, FilterDout_2__1__0, FilterDout_2__2__7, 
               FilterDout_2__2__6, FilterDout_2__2__5, FilterDout_2__2__4, 
               FilterDout_2__2__3, FilterDout_2__2__2, FilterDout_2__2__1, 
               FilterDout_2__2__0, FilterDout_2__3__7, FilterDout_2__3__6, 
               FilterDout_2__3__5, FilterDout_2__3__4, FilterDout_2__3__3, 
               FilterDout_2__3__2, FilterDout_2__3__1, FilterDout_2__3__0, 
               FilterDout_2__4__7, FilterDout_2__4__6, FilterDout_2__4__5, 
               FilterDout_2__4__4, FilterDout_2__4__3, FilterDout_2__4__2, 
               FilterDout_2__4__1, FilterDout_2__4__0, FilterDout_3__0__7, 
               FilterDout_3__0__6, FilterDout_3__0__5, FilterDout_3__0__4, 
               FilterDout_3__0__3, FilterDout_3__0__2, FilterDout_3__0__1, 
               FilterDout_3__0__0, FilterDout_3__1__7, FilterDout_3__1__6, 
               FilterDout_3__1__5, FilterDout_3__1__4, FilterDout_3__1__3, 
               FilterDout_3__1__2, FilterDout_3__1__1, FilterDout_3__1__0, 
               FilterDout_3__2__7, FilterDout_3__2__6, FilterDout_3__2__5, 
               FilterDout_3__2__4, FilterDout_3__2__3, FilterDout_3__2__2, 
               FilterDout_3__2__1, FilterDout_3__2__0, FilterDout_3__3__7, 
               FilterDout_3__3__6, FilterDout_3__3__5, FilterDout_3__3__4, 
               FilterDout_3__3__3, FilterDout_3__3__2, FilterDout_3__3__1, 
               FilterDout_3__3__0, FilterDout_3__4__7, FilterDout_3__4__6, 
               FilterDout_3__4__5, FilterDout_3__4__4, FilterDout_3__4__3, 
               FilterDout_3__4__2, FilterDout_3__4__1, FilterDout_3__4__0, 
               FilterDout_4__0__7, FilterDout_4__0__6, FilterDout_4__0__5, 
               FilterDout_4__0__4, FilterDout_4__0__3, FilterDout_4__0__2, 
               FilterDout_4__0__1, FilterDout_4__0__0, FilterDout_4__1__7, 
               FilterDout_4__1__6, FilterDout_4__1__5, FilterDout_4__1__4, 
               FilterDout_4__1__3, FilterDout_4__1__2, FilterDout_4__1__1, 
               FilterDout_4__1__0, FilterDout_4__2__7, FilterDout_4__2__6, 
               FilterDout_4__2__5, FilterDout_4__2__4, FilterDout_4__2__3, 
               FilterDout_4__2__2, FilterDout_4__2__1, FilterDout_4__2__0, 
               FilterDout_4__3__7, FilterDout_4__3__6, FilterDout_4__3__5, 
               FilterDout_4__3__4, FilterDout_4__3__3, FilterDout_4__3__2, 
               FilterDout_4__3__1, FilterDout_4__3__0, FilterDout_4__4__7, 
               FilterDout_4__4__6, FilterDout_4__4__5, FilterDout_4__4__4, 
               FilterDout_4__4__3, FilterDout_4__4__2, FilterDout_4__4__1, 
               FilterDout_4__4__0, WindowDout_0__0__7, WindowDout_0__0__6, 
               WindowDout_0__0__5, WindowDout_0__0__4, WindowDout_0__0__3, 
               WindowDout_0__0__2, WindowDout_0__0__1, WindowDout_0__0__0, 
               WindowDout_0__1__7, WindowDout_0__1__6, WindowDout_0__1__5, 
               WindowDout_0__1__4, WindowDout_0__1__3, WindowDout_0__1__2, 
               WindowDout_0__1__1, WindowDout_0__1__0, WindowDout_0__2__7, 
               WindowDout_0__2__6, WindowDout_0__2__5, WindowDout_0__2__4, 
               WindowDout_0__2__3, WindowDout_0__2__2, WindowDout_0__2__1, 
               WindowDout_0__2__0, WindowDout_0__3__7, WindowDout_0__3__6, 
               WindowDout_0__3__5, WindowDout_0__3__4, WindowDout_0__3__3, 
               WindowDout_0__3__2, WindowDout_0__3__1, WindowDout_0__3__0, 
               WindowDout_0__4__7, WindowDout_0__4__6, WindowDout_0__4__5, 
               WindowDout_0__4__4, WindowDout_0__4__3, WindowDout_0__4__2, 
               WindowDout_0__4__1, WindowDout_0__4__0, WindowDout_1__0__7, 
               WindowDout_1__0__6, WindowDout_1__0__5, WindowDout_1__0__4, 
               WindowDout_1__0__3, WindowDout_1__0__2, WindowDout_1__0__1, 
               WindowDout_1__0__0, WindowDout_1__1__7, WindowDout_1__1__6, 
               WindowDout_1__1__5, WindowDout_1__1__4, WindowDout_1__1__3, 
               WindowDout_1__1__2, WindowDout_1__1__1, WindowDout_1__1__0, 
               WindowDout_1__2__7, WindowDout_1__2__6, WindowDout_1__2__5, 
               WindowDout_1__2__4, WindowDout_1__2__3, WindowDout_1__2__2, 
               WindowDout_1__2__1, WindowDout_1__2__0, WindowDout_1__3__7, 
               WindowDout_1__3__6, WindowDout_1__3__5, WindowDout_1__3__4, 
               WindowDout_1__3__3, WindowDout_1__3__2, WindowDout_1__3__1, 
               WindowDout_1__3__0, WindowDout_1__4__7, WindowDout_1__4__6, 
               WindowDout_1__4__5, WindowDout_1__4__4, WindowDout_1__4__3, 
               WindowDout_1__4__2, WindowDout_1__4__1, WindowDout_1__4__0, 
               WindowDout_2__0__7, WindowDout_2__0__6, WindowDout_2__0__5, 
               WindowDout_2__0__4, WindowDout_2__0__3, WindowDout_2__0__2, 
               WindowDout_2__0__1, WindowDout_2__0__0, WindowDout_2__1__7, 
               WindowDout_2__1__6, WindowDout_2__1__5, WindowDout_2__1__4, 
               WindowDout_2__1__3, WindowDout_2__1__2, WindowDout_2__1__1, 
               WindowDout_2__1__0, WindowDout_2__2__7, WindowDout_2__2__6, 
               WindowDout_2__2__5, WindowDout_2__2__4, WindowDout_2__2__3, 
               WindowDout_2__2__2, WindowDout_2__2__1, WindowDout_2__2__0, 
               WindowDout_2__3__7, WindowDout_2__3__6, WindowDout_2__3__5, 
               WindowDout_2__3__4, WindowDout_2__3__3, WindowDout_2__3__2, 
               WindowDout_2__3__1, WindowDout_2__3__0, WindowDout_2__4__7, 
               WindowDout_2__4__6, WindowDout_2__4__5, WindowDout_2__4__4, 
               WindowDout_2__4__3, WindowDout_2__4__2, WindowDout_2__4__1, 
               WindowDout_2__4__0, WindowDout_3__0__7, WindowDout_3__0__6, 
               WindowDout_3__0__5, WindowDout_3__0__4, WindowDout_3__0__3, 
               WindowDout_3__0__2, WindowDout_3__0__1, WindowDout_3__0__0, 
               WindowDout_3__1__7, WindowDout_3__1__6, WindowDout_3__1__5, 
               WindowDout_3__1__4, WindowDout_3__1__3, WindowDout_3__1__2, 
               WindowDout_3__1__1, WindowDout_3__1__0, WindowDout_3__2__7, 
               WindowDout_3__2__6, WindowDout_3__2__5, WindowDout_3__2__4, 
               WindowDout_3__2__3, WindowDout_3__2__2, WindowDout_3__2__1, 
               WindowDout_3__2__0, WindowDout_3__3__7, WindowDout_3__3__6, 
               WindowDout_3__3__5, WindowDout_3__3__4, WindowDout_3__3__3, 
               WindowDout_3__3__2, WindowDout_3__3__1, WindowDout_3__3__0, 
               WindowDout_3__4__7, WindowDout_3__4__6, WindowDout_3__4__5, 
               WindowDout_3__4__4, WindowDout_3__4__3, WindowDout_3__4__2, 
               WindowDout_3__4__1, WindowDout_3__4__0, WindowDout_4__0__7, 
               WindowDout_4__0__6, WindowDout_4__0__5, WindowDout_4__0__4, 
               WindowDout_4__0__3, WindowDout_4__0__2, WindowDout_4__0__1, 
               WindowDout_4__0__0, WindowDout_4__1__7, WindowDout_4__1__6, 
               WindowDout_4__1__5, WindowDout_4__1__4, WindowDout_4__1__3, 
               WindowDout_4__1__2, WindowDout_4__1__1, WindowDout_4__1__0, 
               WindowDout_4__2__7, WindowDout_4__2__6, WindowDout_4__2__5, 
               WindowDout_4__2__4, WindowDout_4__2__3, WindowDout_4__2__2, 
               WindowDout_4__2__1, WindowDout_4__2__0, WindowDout_4__3__7, 
               WindowDout_4__3__6, WindowDout_4__3__5, WindowDout_4__3__4, 
               WindowDout_4__3__3, WindowDout_4__3__2, WindowDout_4__3__1, 
               WindowDout_4__3__0, WindowDout_4__4__7, WindowDout_4__4__6, 
               WindowDout_4__4__5, WindowDout_4__4__4, WindowDout_4__4__3, 
               WindowDout_4__4__2, WindowDout_4__4__1, WindowDout_4__4__0, 
               ResultWR, ResultDin, ResultDout ) ;

    input CLK ;
    input RST ;
    input FilterSize ;
    input FilterWR ;
    input WindowWR ;
    input [39:0]Din ;
    output FilterDout_0__0__7 ;
    output FilterDout_0__0__6 ;
    output FilterDout_0__0__5 ;
    output FilterDout_0__0__4 ;
    output FilterDout_0__0__3 ;
    output FilterDout_0__0__2 ;
    output FilterDout_0__0__1 ;
    output FilterDout_0__0__0 ;
    output FilterDout_0__1__7 ;
    output FilterDout_0__1__6 ;
    output FilterDout_0__1__5 ;
    output FilterDout_0__1__4 ;
    output FilterDout_0__1__3 ;
    output FilterDout_0__1__2 ;
    output FilterDout_0__1__1 ;
    output FilterDout_0__1__0 ;
    output FilterDout_0__2__7 ;
    output FilterDout_0__2__6 ;
    output FilterDout_0__2__5 ;
    output FilterDout_0__2__4 ;
    output FilterDout_0__2__3 ;
    output FilterDout_0__2__2 ;
    output FilterDout_0__2__1 ;
    output FilterDout_0__2__0 ;
    output FilterDout_0__3__7 ;
    output FilterDout_0__3__6 ;
    output FilterDout_0__3__5 ;
    output FilterDout_0__3__4 ;
    output FilterDout_0__3__3 ;
    output FilterDout_0__3__2 ;
    output FilterDout_0__3__1 ;
    output FilterDout_0__3__0 ;
    output FilterDout_0__4__7 ;
    output FilterDout_0__4__6 ;
    output FilterDout_0__4__5 ;
    output FilterDout_0__4__4 ;
    output FilterDout_0__4__3 ;
    output FilterDout_0__4__2 ;
    output FilterDout_0__4__1 ;
    output FilterDout_0__4__0 ;
    output FilterDout_1__0__7 ;
    output FilterDout_1__0__6 ;
    output FilterDout_1__0__5 ;
    output FilterDout_1__0__4 ;
    output FilterDout_1__0__3 ;
    output FilterDout_1__0__2 ;
    output FilterDout_1__0__1 ;
    output FilterDout_1__0__0 ;
    output FilterDout_1__1__7 ;
    output FilterDout_1__1__6 ;
    output FilterDout_1__1__5 ;
    output FilterDout_1__1__4 ;
    output FilterDout_1__1__3 ;
    output FilterDout_1__1__2 ;
    output FilterDout_1__1__1 ;
    output FilterDout_1__1__0 ;
    output FilterDout_1__2__7 ;
    output FilterDout_1__2__6 ;
    output FilterDout_1__2__5 ;
    output FilterDout_1__2__4 ;
    output FilterDout_1__2__3 ;
    output FilterDout_1__2__2 ;
    output FilterDout_1__2__1 ;
    output FilterDout_1__2__0 ;
    output FilterDout_1__3__7 ;
    output FilterDout_1__3__6 ;
    output FilterDout_1__3__5 ;
    output FilterDout_1__3__4 ;
    output FilterDout_1__3__3 ;
    output FilterDout_1__3__2 ;
    output FilterDout_1__3__1 ;
    output FilterDout_1__3__0 ;
    output FilterDout_1__4__7 ;
    output FilterDout_1__4__6 ;
    output FilterDout_1__4__5 ;
    output FilterDout_1__4__4 ;
    output FilterDout_1__4__3 ;
    output FilterDout_1__4__2 ;
    output FilterDout_1__4__1 ;
    output FilterDout_1__4__0 ;
    output FilterDout_2__0__7 ;
    output FilterDout_2__0__6 ;
    output FilterDout_2__0__5 ;
    output FilterDout_2__0__4 ;
    output FilterDout_2__0__3 ;
    output FilterDout_2__0__2 ;
    output FilterDout_2__0__1 ;
    output FilterDout_2__0__0 ;
    output FilterDout_2__1__7 ;
    output FilterDout_2__1__6 ;
    output FilterDout_2__1__5 ;
    output FilterDout_2__1__4 ;
    output FilterDout_2__1__3 ;
    output FilterDout_2__1__2 ;
    output FilterDout_2__1__1 ;
    output FilterDout_2__1__0 ;
    output FilterDout_2__2__7 ;
    output FilterDout_2__2__6 ;
    output FilterDout_2__2__5 ;
    output FilterDout_2__2__4 ;
    output FilterDout_2__2__3 ;
    output FilterDout_2__2__2 ;
    output FilterDout_2__2__1 ;
    output FilterDout_2__2__0 ;
    output FilterDout_2__3__7 ;
    output FilterDout_2__3__6 ;
    output FilterDout_2__3__5 ;
    output FilterDout_2__3__4 ;
    output FilterDout_2__3__3 ;
    output FilterDout_2__3__2 ;
    output FilterDout_2__3__1 ;
    output FilterDout_2__3__0 ;
    output FilterDout_2__4__7 ;
    output FilterDout_2__4__6 ;
    output FilterDout_2__4__5 ;
    output FilterDout_2__4__4 ;
    output FilterDout_2__4__3 ;
    output FilterDout_2__4__2 ;
    output FilterDout_2__4__1 ;
    output FilterDout_2__4__0 ;
    output FilterDout_3__0__7 ;
    output FilterDout_3__0__6 ;
    output FilterDout_3__0__5 ;
    output FilterDout_3__0__4 ;
    output FilterDout_3__0__3 ;
    output FilterDout_3__0__2 ;
    output FilterDout_3__0__1 ;
    output FilterDout_3__0__0 ;
    output FilterDout_3__1__7 ;
    output FilterDout_3__1__6 ;
    output FilterDout_3__1__5 ;
    output FilterDout_3__1__4 ;
    output FilterDout_3__1__3 ;
    output FilterDout_3__1__2 ;
    output FilterDout_3__1__1 ;
    output FilterDout_3__1__0 ;
    output FilterDout_3__2__7 ;
    output FilterDout_3__2__6 ;
    output FilterDout_3__2__5 ;
    output FilterDout_3__2__4 ;
    output FilterDout_3__2__3 ;
    output FilterDout_3__2__2 ;
    output FilterDout_3__2__1 ;
    output FilterDout_3__2__0 ;
    output FilterDout_3__3__7 ;
    output FilterDout_3__3__6 ;
    output FilterDout_3__3__5 ;
    output FilterDout_3__3__4 ;
    output FilterDout_3__3__3 ;
    output FilterDout_3__3__2 ;
    output FilterDout_3__3__1 ;
    output FilterDout_3__3__0 ;
    output FilterDout_3__4__7 ;
    output FilterDout_3__4__6 ;
    output FilterDout_3__4__5 ;
    output FilterDout_3__4__4 ;
    output FilterDout_3__4__3 ;
    output FilterDout_3__4__2 ;
    output FilterDout_3__4__1 ;
    output FilterDout_3__4__0 ;
    output FilterDout_4__0__7 ;
    output FilterDout_4__0__6 ;
    output FilterDout_4__0__5 ;
    output FilterDout_4__0__4 ;
    output FilterDout_4__0__3 ;
    output FilterDout_4__0__2 ;
    output FilterDout_4__0__1 ;
    output FilterDout_4__0__0 ;
    output FilterDout_4__1__7 ;
    output FilterDout_4__1__6 ;
    output FilterDout_4__1__5 ;
    output FilterDout_4__1__4 ;
    output FilterDout_4__1__3 ;
    output FilterDout_4__1__2 ;
    output FilterDout_4__1__1 ;
    output FilterDout_4__1__0 ;
    output FilterDout_4__2__7 ;
    output FilterDout_4__2__6 ;
    output FilterDout_4__2__5 ;
    output FilterDout_4__2__4 ;
    output FilterDout_4__2__3 ;
    output FilterDout_4__2__2 ;
    output FilterDout_4__2__1 ;
    output FilterDout_4__2__0 ;
    output FilterDout_4__3__7 ;
    output FilterDout_4__3__6 ;
    output FilterDout_4__3__5 ;
    output FilterDout_4__3__4 ;
    output FilterDout_4__3__3 ;
    output FilterDout_4__3__2 ;
    output FilterDout_4__3__1 ;
    output FilterDout_4__3__0 ;
    output FilterDout_4__4__7 ;
    output FilterDout_4__4__6 ;
    output FilterDout_4__4__5 ;
    output FilterDout_4__4__4 ;
    output FilterDout_4__4__3 ;
    output FilterDout_4__4__2 ;
    output FilterDout_4__4__1 ;
    output FilterDout_4__4__0 ;
    output WindowDout_0__0__7 ;
    output WindowDout_0__0__6 ;
    output WindowDout_0__0__5 ;
    output WindowDout_0__0__4 ;
    output WindowDout_0__0__3 ;
    output WindowDout_0__0__2 ;
    output WindowDout_0__0__1 ;
    output WindowDout_0__0__0 ;
    output WindowDout_0__1__7 ;
    output WindowDout_0__1__6 ;
    output WindowDout_0__1__5 ;
    output WindowDout_0__1__4 ;
    output WindowDout_0__1__3 ;
    output WindowDout_0__1__2 ;
    output WindowDout_0__1__1 ;
    output WindowDout_0__1__0 ;
    output WindowDout_0__2__7 ;
    output WindowDout_0__2__6 ;
    output WindowDout_0__2__5 ;
    output WindowDout_0__2__4 ;
    output WindowDout_0__2__3 ;
    output WindowDout_0__2__2 ;
    output WindowDout_0__2__1 ;
    output WindowDout_0__2__0 ;
    output WindowDout_0__3__7 ;
    output WindowDout_0__3__6 ;
    output WindowDout_0__3__5 ;
    output WindowDout_0__3__4 ;
    output WindowDout_0__3__3 ;
    output WindowDout_0__3__2 ;
    output WindowDout_0__3__1 ;
    output WindowDout_0__3__0 ;
    output WindowDout_0__4__7 ;
    output WindowDout_0__4__6 ;
    output WindowDout_0__4__5 ;
    output WindowDout_0__4__4 ;
    output WindowDout_0__4__3 ;
    output WindowDout_0__4__2 ;
    output WindowDout_0__4__1 ;
    output WindowDout_0__4__0 ;
    output WindowDout_1__0__7 ;
    output WindowDout_1__0__6 ;
    output WindowDout_1__0__5 ;
    output WindowDout_1__0__4 ;
    output WindowDout_1__0__3 ;
    output WindowDout_1__0__2 ;
    output WindowDout_1__0__1 ;
    output WindowDout_1__0__0 ;
    output WindowDout_1__1__7 ;
    output WindowDout_1__1__6 ;
    output WindowDout_1__1__5 ;
    output WindowDout_1__1__4 ;
    output WindowDout_1__1__3 ;
    output WindowDout_1__1__2 ;
    output WindowDout_1__1__1 ;
    output WindowDout_1__1__0 ;
    output WindowDout_1__2__7 ;
    output WindowDout_1__2__6 ;
    output WindowDout_1__2__5 ;
    output WindowDout_1__2__4 ;
    output WindowDout_1__2__3 ;
    output WindowDout_1__2__2 ;
    output WindowDout_1__2__1 ;
    output WindowDout_1__2__0 ;
    output WindowDout_1__3__7 ;
    output WindowDout_1__3__6 ;
    output WindowDout_1__3__5 ;
    output WindowDout_1__3__4 ;
    output WindowDout_1__3__3 ;
    output WindowDout_1__3__2 ;
    output WindowDout_1__3__1 ;
    output WindowDout_1__3__0 ;
    output WindowDout_1__4__7 ;
    output WindowDout_1__4__6 ;
    output WindowDout_1__4__5 ;
    output WindowDout_1__4__4 ;
    output WindowDout_1__4__3 ;
    output WindowDout_1__4__2 ;
    output WindowDout_1__4__1 ;
    output WindowDout_1__4__0 ;
    output WindowDout_2__0__7 ;
    output WindowDout_2__0__6 ;
    output WindowDout_2__0__5 ;
    output WindowDout_2__0__4 ;
    output WindowDout_2__0__3 ;
    output WindowDout_2__0__2 ;
    output WindowDout_2__0__1 ;
    output WindowDout_2__0__0 ;
    output WindowDout_2__1__7 ;
    output WindowDout_2__1__6 ;
    output WindowDout_2__1__5 ;
    output WindowDout_2__1__4 ;
    output WindowDout_2__1__3 ;
    output WindowDout_2__1__2 ;
    output WindowDout_2__1__1 ;
    output WindowDout_2__1__0 ;
    output WindowDout_2__2__7 ;
    output WindowDout_2__2__6 ;
    output WindowDout_2__2__5 ;
    output WindowDout_2__2__4 ;
    output WindowDout_2__2__3 ;
    output WindowDout_2__2__2 ;
    output WindowDout_2__2__1 ;
    output WindowDout_2__2__0 ;
    output WindowDout_2__3__7 ;
    output WindowDout_2__3__6 ;
    output WindowDout_2__3__5 ;
    output WindowDout_2__3__4 ;
    output WindowDout_2__3__3 ;
    output WindowDout_2__3__2 ;
    output WindowDout_2__3__1 ;
    output WindowDout_2__3__0 ;
    output WindowDout_2__4__7 ;
    output WindowDout_2__4__6 ;
    output WindowDout_2__4__5 ;
    output WindowDout_2__4__4 ;
    output WindowDout_2__4__3 ;
    output WindowDout_2__4__2 ;
    output WindowDout_2__4__1 ;
    output WindowDout_2__4__0 ;
    output WindowDout_3__0__7 ;
    output WindowDout_3__0__6 ;
    output WindowDout_3__0__5 ;
    output WindowDout_3__0__4 ;
    output WindowDout_3__0__3 ;
    output WindowDout_3__0__2 ;
    output WindowDout_3__0__1 ;
    output WindowDout_3__0__0 ;
    output WindowDout_3__1__7 ;
    output WindowDout_3__1__6 ;
    output WindowDout_3__1__5 ;
    output WindowDout_3__1__4 ;
    output WindowDout_3__1__3 ;
    output WindowDout_3__1__2 ;
    output WindowDout_3__1__1 ;
    output WindowDout_3__1__0 ;
    output WindowDout_3__2__7 ;
    output WindowDout_3__2__6 ;
    output WindowDout_3__2__5 ;
    output WindowDout_3__2__4 ;
    output WindowDout_3__2__3 ;
    output WindowDout_3__2__2 ;
    output WindowDout_3__2__1 ;
    output WindowDout_3__2__0 ;
    output WindowDout_3__3__7 ;
    output WindowDout_3__3__6 ;
    output WindowDout_3__3__5 ;
    output WindowDout_3__3__4 ;
    output WindowDout_3__3__3 ;
    output WindowDout_3__3__2 ;
    output WindowDout_3__3__1 ;
    output WindowDout_3__3__0 ;
    output WindowDout_3__4__7 ;
    output WindowDout_3__4__6 ;
    output WindowDout_3__4__5 ;
    output WindowDout_3__4__4 ;
    output WindowDout_3__4__3 ;
    output WindowDout_3__4__2 ;
    output WindowDout_3__4__1 ;
    output WindowDout_3__4__0 ;
    output WindowDout_4__0__7 ;
    output WindowDout_4__0__6 ;
    output WindowDout_4__0__5 ;
    output WindowDout_4__0__4 ;
    output WindowDout_4__0__3 ;
    output WindowDout_4__0__2 ;
    output WindowDout_4__0__1 ;
    output WindowDout_4__0__0 ;
    output WindowDout_4__1__7 ;
    output WindowDout_4__1__6 ;
    output WindowDout_4__1__5 ;
    output WindowDout_4__1__4 ;
    output WindowDout_4__1__3 ;
    output WindowDout_4__1__2 ;
    output WindowDout_4__1__1 ;
    output WindowDout_4__1__0 ;
    output WindowDout_4__2__7 ;
    output WindowDout_4__2__6 ;
    output WindowDout_4__2__5 ;
    output WindowDout_4__2__4 ;
    output WindowDout_4__2__3 ;
    output WindowDout_4__2__2 ;
    output WindowDout_4__2__1 ;
    output WindowDout_4__2__0 ;
    output WindowDout_4__3__7 ;
    output WindowDout_4__3__6 ;
    output WindowDout_4__3__5 ;
    output WindowDout_4__3__4 ;
    output WindowDout_4__3__3 ;
    output WindowDout_4__3__2 ;
    output WindowDout_4__3__1 ;
    output WindowDout_4__3__0 ;
    output WindowDout_4__4__7 ;
    output WindowDout_4__4__6 ;
    output WindowDout_4__4__5 ;
    output WindowDout_4__4__4 ;
    output WindowDout_4__4__3 ;
    output WindowDout_4__4__2 ;
    output WindowDout_4__4__1 ;
    output WindowDout_4__4__0 ;
    input ResultWR ;
    input [7:0]ResultDin ;
    output [7:0]ResultDout ;

    wire nx82, nx86, nx96, nx106, nx116, nx126, nx136, nx146, nx156, nx166, 
         nx218, nx228, nx238, nx248, nx258, nx268, nx278, nx288, nx1897, nx1907, 
         nx1917, nx1927, nx1937, nx1947, nx1957, nx1967, nx1981, nx1991, nx2001, 
         nx2011, nx2021, nx2031, nx2041, nx2051, nx2061, nx2071, nx2081, nx2091, 
         nx2101, nx2111, nx2121, nx2131, nx2141, nx2151, nx2161, nx2171, nx2181, 
         nx2191, nx2201, nx2211, nx2221, nx2231, nx2241, nx2251, nx2261, nx2271, 
         nx2281, nx2291, nx2301, nx2311, nx2321, nx2331, nx2341, nx2351, nx2361, 
         nx2371, nx2381, nx2391, nx2401, nx2411, nx2421, nx2431, nx2441, nx2451, 
         nx2461, nx2471, nx2481, nx2491, nx2501, nx2511, nx2521, nx2531, nx2541, 
         nx2551, nx2561, nx2571, nx2581, nx2591, nx2601, nx2611, nx2621, nx2631, 
         nx2641, nx2651, nx2661, nx2671, nx2681, nx2691, nx2701, nx2711, nx2721, 
         nx2731, nx2741, nx2751, nx2761, nx2771, nx2781, nx2791, nx2801, nx2811, 
         nx2821, nx2831, nx2841, nx2851, nx2861, nx2871, nx2881, nx2891, nx2901, 
         nx2911, nx2921, nx2931, nx2941, nx2951, nx2961, nx2971, nx2981, nx2991, 
         nx3001, nx3011, nx3021, nx3031, nx3041, nx3051, nx3061, nx3071, nx3081, 
         nx3091, nx3101, nx3111, nx3121, nx3131, nx3141, nx3151, nx3161, nx3171, 
         nx3181, nx3191, nx3201, nx3211, nx3221, nx3231, nx3241, nx3251, nx3261, 
         nx3271, nx3281, nx3291, nx3301, nx3311, nx3321, nx3331, nx3341, nx3351, 
         nx3361, nx3371, nx3381, nx3391, nx3401, nx3411, nx3421, nx3431, nx3441, 
         nx3451, nx3461, nx3471, nx3481, nx3491, nx3501, nx3511, nx3521, nx3531, 
         nx3541, nx3551, nx3561, nx3571, nx3581, nx3591, nx3601, nx3611, nx3621, 
         nx3631, nx3641, nx3651, nx3661, nx3671, nx3681, nx3691, nx3701, nx3711, 
         nx3721, nx3731, nx3741, nx3751, nx3761, nx3771, nx3781, nx3791, nx3801, 
         nx3811, nx3821, nx3831, nx3841, nx3851, nx3861, nx3871, nx3881, nx3891, 
         nx3901, nx3911, nx3921, nx3931, nx3941, nx3951, nx3961, nx3971, nx3981, 
         nx3991, nx4001, nx4011, nx4021, nx4031, nx4041, nx4051, nx4061, nx4071, 
         nx4081, nx4091, nx4101, nx4111, nx4121, nx4131, nx4141, nx4151, nx4161, 
         nx4171, nx4181, nx4191, nx4201, nx4211, nx4221, nx4231, nx4241, nx4251, 
         nx4261, nx4271, nx4281, nx4291, nx4301, nx4311, nx4321, nx4331, nx4341, 
         nx4351, nx4361, nx4371, nx4381, nx4391, nx4401, nx4411, nx4421, nx4431, 
         nx4441, nx4451, nx4461, nx4471, nx4481, nx4491, nx4501, nx4511, nx4521, 
         nx4531, nx4541, nx4551, nx4561, nx4571, nx4581, nx4591, nx4601, nx4611, 
         nx4621, nx4631, nx4641, nx4651, nx4661, nx4671, nx4681, nx4691, nx4701, 
         nx4711, nx4721, nx4731, nx4741, nx4751, nx4761, nx4771, nx4781, nx4791, 
         nx4801, nx4811, nx4821, nx4831, nx4841, nx4851, nx4861, nx4871, nx4881, 
         nx4891, nx4901, nx4911, nx4921, nx4931, nx4941, nx4951, nx4961, nx4971, 
         nx4981, nx4991, nx5001, nx5011, nx5021, nx5031, nx5041, nx5051, nx5061, 
         nx5071, nx5081, nx5091, nx5101, nx5111, nx5121, nx5131, nx5141, nx5151, 
         nx5161, nx5171, nx5181, nx5191, nx5201, nx5211, nx5221, nx5231, nx5241, 
         nx5251, nx5261, nx5271, nx5281, nx5291, nx5301, nx5311, nx5321, nx5331, 
         nx5341, nx5351, nx5361, nx5371, nx5381, nx5391, nx5401, nx5411, nx5421, 
         nx5431, nx5441, nx5451, nx5461, nx5471, nx5481, nx5491, nx5501, nx5511, 
         nx5521, nx5531, nx5541, nx5551, nx5561, nx5571, nx5581, nx5591, nx5601, 
         nx5611, nx5621, nx5631, nx5641, nx5651, nx5661, nx5671, nx5681, nx5691, 
         nx5701, nx5711, nx5721, nx5731, nx5741, nx5751, nx5761, nx5771, nx5781, 
         nx5791, nx5801, nx5811, nx5821, nx5831, nx5841, nx5851, nx5861, nx5871, 
         nx5881, nx5891, nx5901, nx5911, nx5921, nx5931, nx5941, nx5951, nx5961, 
         nx5971, nx6008, nx6075, nx6149, nx6152, nx6156, nx6158, nx6162, nx6164, 
         nx6168, nx6170, nx6174, nx6176, nx6180, nx6182, nx6186, nx6188, nx6192, 
         nx6194, nx6198, nx6200, nx6204, nx6206, nx6210, nx6212, nx6216, nx6218, 
         nx6222, nx6224, nx6228, nx6230, nx6234, nx6236, nx6240, nx6242, nx6318, 
         nx6320, nx6324, nx6326, nx6330, nx6332, nx6336, nx6338, nx6342, nx6344, 
         nx6348, nx6350, nx6354, nx6356, nx6360, nx6362, nx6366, nx6368, nx6372, 
         nx6374, nx6378, nx6380, nx6384, nx6386, nx6390, nx6392, nx6396, nx6398, 
         nx6402, nx6404, nx6408, nx6410, nx6486, nx6488, nx6492, nx6494, nx6498, 
         nx6500, nx6504, nx6506, nx6510, nx6512, nx6516, nx6518, nx6522, nx6524, 
         nx6528, nx6530, nx6534, nx6536, nx6540, nx6542, nx6546, nx6548, nx6552, 
         nx6554, nx6558, nx6560, nx6564, nx6566, nx6570, nx6572, nx6576, nx6578, 
         nx6582, nx6584, nx6588, nx6590, nx6594, nx6596, nx6600, nx6602, nx6606, 
         nx6608, nx6612, nx6614, nx6618, nx6620, nx6624, nx6626, nx6630, nx6632, 
         nx6636, nx6638, nx6642, nx6644, nx6648, nx6650, nx6654, nx6656, nx6660, 
         nx6662, nx6666, nx6668, nx6672, nx6674, nx6678, nx6680, nx6684, nx6686, 
         nx6690, nx6692, nx6696, nx6698, nx6702, nx6704, nx6708, nx6710, nx6714, 
         nx6716, nx6720, nx6722, nx6726, nx6728, nx6732, nx6734, nx6738, nx6740, 
         nx6744, nx6746, nx6750, nx6752, nx6756, nx6758, nx6762, nx6764, nx6768, 
         nx6770, nx6774, nx6776, nx6780, nx6782, nx6786, nx6788, nx6792, nx6794, 
         nx6798, nx6800, nx6804, nx6806, nx6810, nx6812, nx6816, nx6818, nx6822, 
         nx6824, nx6828, nx6830, nx6834, nx6836, nx6840, nx6842, nx6846, nx6848, 
         nx6852, nx6854, nx6858, nx6860, nx6864, nx6866, nx6870, nx6872, nx6876, 
         nx6878, nx6882, nx6884, nx6888, nx6890, nx6894, nx6896, nx6900, nx6902, 
         nx6906, nx6908, nx6912, nx6914, nx6918, nx6920, nx6924, nx6926, nx6930, 
         nx6932, nx6936, nx6938, nx6942, nx6944, nx6948, nx6950, nx6954, nx6956, 
         nx6960, nx6962, nx6966, nx7016, nx7090, nx7093, nx7097, nx7099, nx7103, 
         nx7105, nx7109, nx7111, nx7115, nx7117, nx7121, nx7123, nx7127, nx7129, 
         nx7133, nx7135, nx7139, nx7141, nx7145, nx7147, nx7151, nx7153, nx7157, 
         nx7159, nx7163, nx7165, nx7169, nx7171, nx7175, nx7177, nx7181, nx7183, 
         nx7259, nx7261, nx7265, nx7267, nx7271, nx7273, nx7277, nx7279, nx7283, 
         nx7285, nx7289, nx7291, nx7295, nx7297, nx7301, nx7303, nx7307, nx7309, 
         nx7313, nx7315, nx7319, nx7321, nx7325, nx7327, nx7331, nx7333, nx7337, 
         nx7339, nx7343, nx7345, nx7349, nx7351, nx7427, nx7429, nx7433, nx7435, 
         nx7439, nx7441, nx7445, nx7447, nx7451, nx7453, nx7457, nx7459, nx7463, 
         nx7465, nx7469, nx7471, nx7475, nx7477, nx7481, nx7483, nx7487, nx7489, 
         nx7493, nx7495, nx7499, nx7501, nx7505, nx7507, nx7511, nx7513, nx7517, 
         nx7519, nx7523, nx7525, nx7529, nx7531, nx7535, nx7537, nx7541, nx7543, 
         nx7547, nx7549, nx7553, nx7555, nx7559, nx7561, nx7565, nx7567, nx7571, 
         nx7573, nx7577, nx7579, nx7583, nx7585, nx7589, nx7591, nx7595, nx7597, 
         nx7601, nx7603, nx7607, nx7609, nx7613, nx7615, nx7619, nx7621, nx7625, 
         nx7627, nx7631, nx7633, nx7637, nx7639, nx7643, nx7645, nx7649, nx7651, 
         nx7655, nx7657, nx7661, nx7663, nx7667, nx7669, nx7673, nx7675, nx7679, 
         nx7681, nx7685, nx7687, nx7691, nx7693, nx7697, nx7699, nx7703, nx7705, 
         nx7709, nx7711, nx7715, nx7717, nx7721, nx7723, nx7727, nx7729, nx7733, 
         nx7735, nx7739, nx7741, nx7745, nx7747, nx7751, nx7753, nx7757, nx7759, 
         nx7763, nx7765, nx7769, nx7771, nx7775, nx7777, nx7781, nx7783, nx7787, 
         nx7789, nx7793, nx7795, nx7799, nx7801, nx7805, nx7807, nx7811, nx7813, 
         nx7817, nx7819, nx7823, nx7825, nx7829, nx7831, nx7835, nx7837, nx7841, 
         nx7843, nx7847, nx7849, nx7853, nx7855, nx7859, nx7861, nx7865, nx7867, 
         nx7871, nx7873, nx7877, nx7879, nx7883, nx7885, nx7889, nx7891, nx7895, 
         nx7897, nx7901, nx7903, nx7910, nx7912, nx7914, nx7916, nx7918, nx7920, 
         nx7922, nx7924, nx7926, nx7928, nx7930, nx7932, nx7934, nx7936, nx7938, 
         nx7940, nx7942, nx7944, nx7946, nx7948, nx7950, nx7952, nx7954, nx7956, 
         nx7958, nx7960, nx7962, nx7964, nx7966, nx7968, nx7970, nx7972, nx7974, 
         nx7976, nx7978, nx7980, nx7982, nx7984, nx7986, nx7988, nx7990, nx7992, 
         nx7994, nx7996, nx7998, nx8000, nx8002, nx8004, nx8006, nx8008, nx8010, 
         nx8012, nx8014, nx8016, nx8018, nx8020, nx8022, nx8024, nx8026, nx8028, 
         nx8030, nx8032, nx8034, nx8036, nx8042, nx8044, nx8046, nx8048, nx8050, 
         nx8052, nx8054, nx8056, nx8058, nx8060, nx8062, nx8064, nx8066, nx8068, 
         nx8070, nx8074, nx8076, nx8078, nx8080, nx8086, nx8088, nx8090, nx8092, 
         nx8104, nx8106, nx8108, nx8110, nx8112, nx8114, nx8116, nx8118, nx8120, 
         nx8122, nx8126, nx8128, nx8130, nx8132, nx8134, nx8138, nx8140, nx8142, 
         nx8144, nx8160, nx8162, nx8164, nx8166, nx8168, nx8170, nx8172, nx8174, 
         nx8176, nx8178, nx8180, nx8186, nx8188, nx8190, nx8192, nx8194, nx8198, 
         nx8200, nx8202, nx8204, nx8206, nx8208, nx8210, nx8212, nx8214, nx8216, 
         nx8218, nx8220, nx8222, nx8224, nx8226, nx8236, nx8238, nx8240, nx8242, 
         nx8244, nx8246, nx8248, nx8250, nx8252, nx8254, nx8256, nx8258, nx8260, 
         nx8262, nx8264, nx8266, nx8268, nx8270, nx8272, nx8274, nx8276, nx8278, 
         nx8280, nx8282, nx8284, nx8286, nx8288, nx8290, nx8292, nx8294, nx8300, 
         nx8302;
    wire [183:0] \$dummy ;




    dff RESULT_REG_reg_Dout_0 (.Q (ResultDout[0]), .QB (\$dummy [0]), .D (nx1897
        ), .CLK (CLK)) ;
    nor02ii ix1898 (.Y (nx1897), .A0 (RST), .A1 (ResultDout[0])) ;
    dff RESULT_REG_reg_Dout_1 (.Q (ResultDout[1]), .QB (\$dummy [1]), .D (nx1907
        ), .CLK (CLK)) ;
    nor02ii ix1908 (.Y (nx1907), .A0 (RST), .A1 (ResultDout[1])) ;
    dff RESULT_REG_reg_Dout_2 (.Q (ResultDout[2]), .QB (\$dummy [2]), .D (nx1917
        ), .CLK (CLK)) ;
    nor02ii ix1918 (.Y (nx1917), .A0 (RST), .A1 (ResultDout[2])) ;
    dff RESULT_REG_reg_Dout_3 (.Q (ResultDout[3]), .QB (\$dummy [3]), .D (nx1927
        ), .CLK (CLK)) ;
    nor02ii ix1928 (.Y (nx1927), .A0 (RST), .A1 (ResultDout[3])) ;
    dff RESULT_REG_reg_Dout_4 (.Q (ResultDout[4]), .QB (\$dummy [4]), .D (nx1937
        ), .CLK (CLK)) ;
    nor02ii ix1938 (.Y (nx1937), .A0 (RST), .A1 (ResultDout[4])) ;
    dff RESULT_REG_reg_Dout_5 (.Q (ResultDout[5]), .QB (\$dummy [5]), .D (nx1947
        ), .CLK (CLK)) ;
    nor02ii ix1948 (.Y (nx1947), .A0 (RST), .A1 (ResultDout[5])) ;
    dff RESULT_REG_reg_Dout_6 (.Q (ResultDout[6]), .QB (\$dummy [6]), .D (nx1957
        ), .CLK (CLK)) ;
    nor02ii ix1958 (.Y (nx1957), .A0 (RST), .A1 (ResultDout[6])) ;
    dff RESULT_REG_reg_Dout_7 (.Q (ResultDout[7]), .QB (\$dummy [7]), .D (nx1967
        ), .CLK (CLK)) ;
    nor02ii ix1968 (.Y (nx1967), .A0 (RST), .A1 (ResultDout[7])) ;
    dff L0_4_L1_4_Wij_reg_Dout_0 (.Q (WindowDout_4__4__0), .QB (\$dummy [8]), .D (
        nx1981), .CLK (CLK)) ;
    nor02ii ix87 (.Y (nx86), .A0 (RST), .A1 (Din[32])) ;
    aoi21 ix6009 (.Y (nx6008), .A0 (WindowWR), .A1 (FilterSize), .B0 (RST)) ;
    dff L0_4_L1_4_Wij_reg_Dout_1 (.Q (WindowDout_4__4__1), .QB (\$dummy [9]), .D (
        nx1991), .CLK (CLK)) ;
    nor02ii ix97 (.Y (nx96), .A0 (RST), .A1 (Din[33])) ;
    dff L0_4_L1_4_Wij_reg_Dout_2 (.Q (WindowDout_4__4__2), .QB (\$dummy [10]), .D (
        nx2001), .CLK (CLK)) ;
    nor02ii ix107 (.Y (nx106), .A0 (RST), .A1 (Din[34])) ;
    dff L0_4_L1_4_Wij_reg_Dout_3 (.Q (WindowDout_4__4__3), .QB (\$dummy [11]), .D (
        nx2011), .CLK (CLK)) ;
    nor02ii ix117 (.Y (nx116), .A0 (RST), .A1 (Din[35])) ;
    dff L0_4_L1_4_Wij_reg_Dout_4 (.Q (WindowDout_4__4__4), .QB (\$dummy [12]), .D (
        nx2021), .CLK (CLK)) ;
    nor02ii ix127 (.Y (nx126), .A0 (RST), .A1 (Din[36])) ;
    dff L0_4_L1_4_Wij_reg_Dout_5 (.Q (WindowDout_4__4__5), .QB (\$dummy [13]), .D (
        nx2031), .CLK (CLK)) ;
    nor02ii ix137 (.Y (nx136), .A0 (RST), .A1 (Din[37])) ;
    dff L0_4_L1_4_Wij_reg_Dout_6 (.Q (WindowDout_4__4__6), .QB (\$dummy [14]), .D (
        nx2041), .CLK (CLK)) ;
    nor02ii ix147 (.Y (nx146), .A0 (RST), .A1 (Din[38])) ;
    dff L0_4_L1_4_Wij_reg_Dout_7 (.Q (WindowDout_4__4__7), .QB (\$dummy [15]), .D (
        nx2051), .CLK (CLK)) ;
    nor02ii ix157 (.Y (nx156), .A0 (RST), .A1 (Din[39])) ;
    dff L0_4_L1_3_Wij_reg_Dout_0 (.Q (WindowDout_4__3__0), .QB (\$dummy [16]), .D (
        nx2141), .CLK (CLK)) ;
    nor02ii ix219 (.Y (nx218), .A0 (RST), .A1 (Din[24])) ;
    dff L0_4_L1_3_Wij_reg_Dout_1 (.Q (WindowDout_4__3__1), .QB (\$dummy [17]), .D (
        nx2151), .CLK (CLK)) ;
    nor02ii ix229 (.Y (nx228), .A0 (RST), .A1 (Din[25])) ;
    dff L0_4_L1_3_Wij_reg_Dout_2 (.Q (WindowDout_4__3__2), .QB (\$dummy [18]), .D (
        nx2161), .CLK (CLK)) ;
    nor02ii ix239 (.Y (nx238), .A0 (RST), .A1 (Din[26])) ;
    dff L0_4_L1_3_Wij_reg_Dout_3 (.Q (WindowDout_4__3__3), .QB (\$dummy [19]), .D (
        nx2171), .CLK (CLK)) ;
    nor02ii ix249 (.Y (nx248), .A0 (RST), .A1 (Din[27])) ;
    dff L0_4_L1_3_Wij_reg_Dout_4 (.Q (WindowDout_4__3__4), .QB (\$dummy [20]), .D (
        nx2181), .CLK (CLK)) ;
    nor02ii ix259 (.Y (nx258), .A0 (RST), .A1 (Din[28])) ;
    dff L0_4_L1_3_Wij_reg_Dout_5 (.Q (WindowDout_4__3__5), .QB (\$dummy [21]), .D (
        nx2191), .CLK (CLK)) ;
    nor02ii ix269 (.Y (nx268), .A0 (RST), .A1 (Din[29])) ;
    dff L0_4_L1_3_Wij_reg_Dout_6 (.Q (WindowDout_4__3__6), .QB (\$dummy [22]), .D (
        nx2201), .CLK (CLK)) ;
    nor02ii ix279 (.Y (nx278), .A0 (RST), .A1 (Din[30])) ;
    dff L0_4_L1_3_Wij_reg_Dout_7 (.Q (WindowDout_4__3__7), .QB (\$dummy [23]), .D (
        nx2211), .CLK (CLK)) ;
    nor02ii ix289 (.Y (nx288), .A0 (RST), .A1 (Din[31])) ;
    dff L0_4_L1_2_Wij_reg_Dout_0 (.Q (WindowDout_4__2__0), .QB (\$dummy [24]), .D (
        nx2301), .CLK (CLK)) ;
    ao32 ix2302 (.Y (nx2301), .A0 (Din[16]), .A1 (nx8052), .A2 (WindowWR), .B0 (
         WindowDout_4__2__0), .B1 (nx8160)) ;
    nor02_2x ix6076 (.Y (nx6075), .A0 (WindowWR), .A1 (RST)) ;
    dff L0_4_L1_2_Wij_reg_Dout_1 (.Q (WindowDout_4__2__1), .QB (\$dummy [25]), .D (
        nx2311), .CLK (CLK)) ;
    ao32 ix2312 (.Y (nx2311), .A0 (Din[17]), .A1 (nx8052), .A2 (WindowWR), .B0 (
         WindowDout_4__2__1), .B1 (nx8160)) ;
    dff L0_4_L1_2_Wij_reg_Dout_2 (.Q (WindowDout_4__2__2), .QB (\$dummy [26]), .D (
        nx2321), .CLK (CLK)) ;
    ao32 ix2322 (.Y (nx2321), .A0 (Din[18]), .A1 (nx8052), .A2 (WindowWR), .B0 (
         WindowDout_4__2__2), .B1 (nx8160)) ;
    dff L0_4_L1_2_Wij_reg_Dout_3 (.Q (WindowDout_4__2__3), .QB (\$dummy [27]), .D (
        nx2331), .CLK (CLK)) ;
    ao32 ix2332 (.Y (nx2331), .A0 (Din[19]), .A1 (nx8052), .A2 (WindowWR), .B0 (
         WindowDout_4__2__3), .B1 (nx8160)) ;
    dff L0_4_L1_2_Wij_reg_Dout_4 (.Q (WindowDout_4__2__4), .QB (\$dummy [28]), .D (
        nx2341), .CLK (CLK)) ;
    ao32 ix2342 (.Y (nx2341), .A0 (Din[20]), .A1 (nx8052), .A2 (WindowWR), .B0 (
         WindowDout_4__2__4), .B1 (nx8160)) ;
    dff L0_4_L1_2_Wij_reg_Dout_5 (.Q (WindowDout_4__2__5), .QB (\$dummy [29]), .D (
        nx2351), .CLK (CLK)) ;
    ao32 ix2352 (.Y (nx2351), .A0 (Din[21]), .A1 (nx8052), .A2 (WindowWR), .B0 (
         WindowDout_4__2__5), .B1 (nx8160)) ;
    dff L0_4_L1_2_Wij_reg_Dout_6 (.Q (WindowDout_4__2__6), .QB (\$dummy [30]), .D (
        nx2361), .CLK (CLK)) ;
    ao32 ix2362 (.Y (nx2361), .A0 (Din[22]), .A1 (nx8052), .A2 (WindowWR), .B0 (
         WindowDout_4__2__6), .B1 (nx8160)) ;
    dff L0_4_L1_2_Wij_reg_Dout_7 (.Q (WindowDout_4__2__7), .QB (\$dummy [31]), .D (
        nx2371), .CLK (CLK)) ;
    ao32 ix2372 (.Y (nx2371), .A0 (Din[23]), .A1 (nx8054), .A2 (WindowWR), .B0 (
         WindowDout_4__2__7), .B1 (nx8162)) ;
    dff L0_4_L1_1_Wij_reg_Dout_0 (.Q (WindowDout_4__1__0), .QB (\$dummy [32]), .D (
        nx2461), .CLK (CLK)) ;
    ao32 ix2462 (.Y (nx2461), .A0 (Din[8]), .A1 (nx8054), .A2 (WindowWR), .B0 (
         WindowDout_4__1__0), .B1 (nx8162)) ;
    dff L0_4_L1_1_Wij_reg_Dout_1 (.Q (WindowDout_4__1__1), .QB (\$dummy [33]), .D (
        nx2471), .CLK (CLK)) ;
    ao32 ix2472 (.Y (nx2471), .A0 (Din[9]), .A1 (nx8054), .A2 (WindowWR), .B0 (
         WindowDout_4__1__1), .B1 (nx8162)) ;
    dff L0_4_L1_1_Wij_reg_Dout_2 (.Q (WindowDout_4__1__2), .QB (\$dummy [34]), .D (
        nx2481), .CLK (CLK)) ;
    ao32 ix2482 (.Y (nx2481), .A0 (Din[10]), .A1 (nx8054), .A2 (WindowWR), .B0 (
         WindowDout_4__1__2), .B1 (nx8162)) ;
    dff L0_4_L1_1_Wij_reg_Dout_3 (.Q (WindowDout_4__1__3), .QB (\$dummy [35]), .D (
        nx2491), .CLK (CLK)) ;
    ao32 ix2492 (.Y (nx2491), .A0 (Din[11]), .A1 (nx8054), .A2 (WindowWR), .B0 (
         WindowDout_4__1__3), .B1 (nx8162)) ;
    dff L0_4_L1_1_Wij_reg_Dout_4 (.Q (WindowDout_4__1__4), .QB (\$dummy [36]), .D (
        nx2501), .CLK (CLK)) ;
    ao32 ix2502 (.Y (nx2501), .A0 (Din[12]), .A1 (nx8054), .A2 (WindowWR), .B0 (
         WindowDout_4__1__4), .B1 (nx8162)) ;
    dff L0_4_L1_1_Wij_reg_Dout_5 (.Q (WindowDout_4__1__5), .QB (\$dummy [37]), .D (
        nx2511), .CLK (CLK)) ;
    ao32 ix2512 (.Y (nx2511), .A0 (Din[13]), .A1 (nx8054), .A2 (WindowWR), .B0 (
         WindowDout_4__1__5), .B1 (nx8162)) ;
    dff L0_4_L1_1_Wij_reg_Dout_6 (.Q (WindowDout_4__1__6), .QB (\$dummy [38]), .D (
        nx2521), .CLK (CLK)) ;
    ao32 ix2522 (.Y (nx2521), .A0 (Din[14]), .A1 (nx8056), .A2 (WindowWR), .B0 (
         WindowDout_4__1__6), .B1 (nx8164)) ;
    dff L0_4_L1_1_Wij_reg_Dout_7 (.Q (WindowDout_4__1__7), .QB (\$dummy [39]), .D (
        nx2531), .CLK (CLK)) ;
    ao32 ix2532 (.Y (nx2531), .A0 (Din[15]), .A1 (nx8056), .A2 (WindowWR), .B0 (
         WindowDout_4__1__7), .B1 (nx8164)) ;
    dff L0_4_L1_0_Wij_reg_Dout_0 (.Q (WindowDout_4__0__0), .QB (\$dummy [40]), .D (
        nx2621), .CLK (CLK)) ;
    ao32 ix2622 (.Y (nx2621), .A0 (Din[0]), .A1 (nx8056), .A2 (WindowWR), .B0 (
         WindowDout_4__0__0), .B1 (nx8164)) ;
    dff L0_4_L1_0_Wij_reg_Dout_1 (.Q (WindowDout_4__0__1), .QB (\$dummy [41]), .D (
        nx2631), .CLK (CLK)) ;
    ao32 ix2632 (.Y (nx2631), .A0 (Din[1]), .A1 (nx8056), .A2 (WindowWR), .B0 (
         WindowDout_4__0__1), .B1 (nx8164)) ;
    dff L0_4_L1_0_Wij_reg_Dout_2 (.Q (WindowDout_4__0__2), .QB (\$dummy [42]), .D (
        nx2641), .CLK (CLK)) ;
    ao32 ix2642 (.Y (nx2641), .A0 (Din[2]), .A1 (nx8056), .A2 (WindowWR), .B0 (
         WindowDout_4__0__2), .B1 (nx8164)) ;
    dff L0_4_L1_0_Wij_reg_Dout_3 (.Q (WindowDout_4__0__3), .QB (\$dummy [43]), .D (
        nx2651), .CLK (CLK)) ;
    ao32 ix2652 (.Y (nx2651), .A0 (Din[3]), .A1 (nx8056), .A2 (WindowWR), .B0 (
         WindowDout_4__0__3), .B1 (nx8164)) ;
    dff L0_4_L1_0_Wij_reg_Dout_4 (.Q (WindowDout_4__0__4), .QB (\$dummy [44]), .D (
        nx2661), .CLK (CLK)) ;
    ao32 ix2662 (.Y (nx2661), .A0 (Din[4]), .A1 (nx8056), .A2 (WindowWR), .B0 (
         WindowDout_4__0__4), .B1 (nx8164)) ;
    dff L0_4_L1_0_Wij_reg_Dout_5 (.Q (WindowDout_4__0__5), .QB (\$dummy [45]), .D (
        nx2671), .CLK (CLK)) ;
    ao32 ix2672 (.Y (nx2671), .A0 (Din[5]), .A1 (nx8058), .A2 (WindowWR), .B0 (
         WindowDout_4__0__5), .B1 (nx8166)) ;
    dff L0_4_L1_0_Wij_reg_Dout_6 (.Q (WindowDout_4__0__6), .QB (\$dummy [46]), .D (
        nx2681), .CLK (CLK)) ;
    ao32 ix2682 (.Y (nx2681), .A0 (Din[6]), .A1 (nx8058), .A2 (WindowWR), .B0 (
         WindowDout_4__0__6), .B1 (nx8166)) ;
    dff L0_4_L1_0_Wij_reg_Dout_7 (.Q (WindowDout_4__0__7), .QB (\$dummy [47]), .D (
        nx2691), .CLK (CLK)) ;
    ao32 ix2692 (.Y (nx2691), .A0 (Din[7]), .A1 (nx8058), .A2 (WindowWR), .B0 (
         WindowDout_4__0__7), .B1 (nx8166)) ;
    oai21 ix2782 (.Y (nx2781), .A0 (nx6149), .A1 (nx7910), .B0 (nx6152)) ;
    dff L0_3_L1_4_Wij_reg_Dout_0 (.Q (WindowDout_3__4__0), .QB (nx6149), .D (
        nx2781), .CLK (CLK)) ;
    nand03 ix6153 (.Y (nx6152), .A0 (nx8058), .A1 (WindowDout_4__4__0), .A2 (
           nx7910)) ;
    oai21 ix2792 (.Y (nx2791), .A0 (nx6156), .A1 (nx7910), .B0 (nx6158)) ;
    dff L0_3_L1_4_Wij_reg_Dout_1 (.Q (WindowDout_3__4__1), .QB (nx6156), .D (
        nx2791), .CLK (CLK)) ;
    nand03 ix6159 (.Y (nx6158), .A0 (nx8058), .A1 (WindowDout_4__4__1), .A2 (
           nx7910)) ;
    oai21 ix2802 (.Y (nx2801), .A0 (nx6162), .A1 (nx7910), .B0 (nx6164)) ;
    dff L0_3_L1_4_Wij_reg_Dout_2 (.Q (WindowDout_3__4__2), .QB (nx6162), .D (
        nx2801), .CLK (CLK)) ;
    nand03 ix6165 (.Y (nx6164), .A0 (nx8058), .A1 (WindowDout_4__4__2), .A2 (
           nx7910)) ;
    oai21 ix2812 (.Y (nx2811), .A0 (nx6168), .A1 (nx7910), .B0 (nx6170)) ;
    dff L0_3_L1_4_Wij_reg_Dout_3 (.Q (WindowDout_3__4__3), .QB (nx6168), .D (
        nx2811), .CLK (CLK)) ;
    nand03 ix6171 (.Y (nx6170), .A0 (nx8058), .A1 (WindowDout_4__4__3), .A2 (
           nx7912)) ;
    oai21 ix2822 (.Y (nx2821), .A0 (nx6174), .A1 (nx7912), .B0 (nx6176)) ;
    dff L0_3_L1_4_Wij_reg_Dout_4 (.Q (WindowDout_3__4__4), .QB (nx6174), .D (
        nx2821), .CLK (CLK)) ;
    nand03 ix6177 (.Y (nx6176), .A0 (nx8060), .A1 (WindowDout_4__4__4), .A2 (
           nx7912)) ;
    oai21 ix2832 (.Y (nx2831), .A0 (nx6180), .A1 (nx7912), .B0 (nx6182)) ;
    dff L0_3_L1_4_Wij_reg_Dout_5 (.Q (WindowDout_3__4__5), .QB (nx6180), .D (
        nx2831), .CLK (CLK)) ;
    nand03 ix6183 (.Y (nx6182), .A0 (nx8060), .A1 (WindowDout_4__4__5), .A2 (
           nx7912)) ;
    oai21 ix2842 (.Y (nx2841), .A0 (nx6186), .A1 (nx7912), .B0 (nx6188)) ;
    dff L0_3_L1_4_Wij_reg_Dout_6 (.Q (WindowDout_3__4__6), .QB (nx6186), .D (
        nx2841), .CLK (CLK)) ;
    nand03 ix6189 (.Y (nx6188), .A0 (nx8060), .A1 (WindowDout_4__4__6), .A2 (
           nx7912)) ;
    oai21 ix2852 (.Y (nx2851), .A0 (nx6192), .A1 (nx7914), .B0 (nx6194)) ;
    dff L0_3_L1_4_Wij_reg_Dout_7 (.Q (WindowDout_3__4__7), .QB (nx6192), .D (
        nx2851), .CLK (CLK)) ;
    nand03 ix6195 (.Y (nx6194), .A0 (nx8060), .A1 (WindowDout_4__4__7), .A2 (
           nx7914)) ;
    oai21 ix2942 (.Y (nx2941), .A0 (nx6198), .A1 (nx7914), .B0 (nx6200)) ;
    dff L0_3_L1_3_Wij_reg_Dout_0 (.Q (WindowDout_3__3__0), .QB (nx6198), .D (
        nx2941), .CLK (CLK)) ;
    nand03 ix6201 (.Y (nx6200), .A0 (nx8060), .A1 (WindowDout_4__3__0), .A2 (
           nx7914)) ;
    oai21 ix2952 (.Y (nx2951), .A0 (nx6204), .A1 (nx7914), .B0 (nx6206)) ;
    dff L0_3_L1_3_Wij_reg_Dout_1 (.Q (WindowDout_3__3__1), .QB (nx6204), .D (
        nx2951), .CLK (CLK)) ;
    nand03 ix6207 (.Y (nx6206), .A0 (nx8060), .A1 (WindowDout_4__3__1), .A2 (
           nx7914)) ;
    oai21 ix2962 (.Y (nx2961), .A0 (nx6210), .A1 (nx7914), .B0 (nx6212)) ;
    dff L0_3_L1_3_Wij_reg_Dout_2 (.Q (WindowDout_3__3__2), .QB (nx6210), .D (
        nx2961), .CLK (CLK)) ;
    nand03 ix6213 (.Y (nx6212), .A0 (nx8060), .A1 (WindowDout_4__3__2), .A2 (
           nx7916)) ;
    oai21 ix2972 (.Y (nx2971), .A0 (nx6216), .A1 (nx7916), .B0 (nx6218)) ;
    dff L0_3_L1_3_Wij_reg_Dout_3 (.Q (WindowDout_3__3__3), .QB (nx6216), .D (
        nx2971), .CLK (CLK)) ;
    nand03 ix6219 (.Y (nx6218), .A0 (nx8062), .A1 (WindowDout_4__3__3), .A2 (
           nx7916)) ;
    oai21 ix2982 (.Y (nx2981), .A0 (nx6222), .A1 (nx7916), .B0 (nx6224)) ;
    dff L0_3_L1_3_Wij_reg_Dout_4 (.Q (WindowDout_3__3__4), .QB (nx6222), .D (
        nx2981), .CLK (CLK)) ;
    nand03 ix6225 (.Y (nx6224), .A0 (nx8062), .A1 (WindowDout_4__3__4), .A2 (
           nx7916)) ;
    oai21 ix2992 (.Y (nx2991), .A0 (nx6228), .A1 (nx7916), .B0 (nx6230)) ;
    dff L0_3_L1_3_Wij_reg_Dout_5 (.Q (WindowDout_3__3__5), .QB (nx6228), .D (
        nx2991), .CLK (CLK)) ;
    nand03 ix6231 (.Y (nx6230), .A0 (nx8062), .A1 (WindowDout_4__3__5), .A2 (
           nx7916)) ;
    oai21 ix3002 (.Y (nx3001), .A0 (nx6234), .A1 (nx7918), .B0 (nx6236)) ;
    dff L0_3_L1_3_Wij_reg_Dout_6 (.Q (WindowDout_3__3__6), .QB (nx6234), .D (
        nx3001), .CLK (CLK)) ;
    nand03 ix6237 (.Y (nx6236), .A0 (nx8062), .A1 (WindowDout_4__3__6), .A2 (
           nx7918)) ;
    oai21 ix3012 (.Y (nx3011), .A0 (nx6240), .A1 (nx7918), .B0 (nx6242)) ;
    dff L0_3_L1_3_Wij_reg_Dout_7 (.Q (WindowDout_3__3__7), .QB (nx6240), .D (
        nx3011), .CLK (CLK)) ;
    nand03 ix6243 (.Y (nx6242), .A0 (nx8062), .A1 (WindowDout_4__3__7), .A2 (
           nx7918)) ;
    dff L0_3_L1_2_Wij_reg_Dout_0 (.Q (WindowDout_3__2__0), .QB (\$dummy [48]), .D (
        nx3101), .CLK (CLK)) ;
    ao32 ix3102 (.Y (nx3101), .A0 (nx8062), .A1 (WindowDout_4__2__0), .A2 (
         WindowWR), .B0 (WindowDout_3__2__0), .B1 (nx8166)) ;
    dff L0_3_L1_2_Wij_reg_Dout_1 (.Q (WindowDout_3__2__1), .QB (\$dummy [49]), .D (
        nx3111), .CLK (CLK)) ;
    ao32 ix3112 (.Y (nx3111), .A0 (nx8062), .A1 (WindowDout_4__2__1), .A2 (
         WindowWR), .B0 (WindowDout_3__2__1), .B1 (nx8166)) ;
    dff L0_3_L1_2_Wij_reg_Dout_2 (.Q (WindowDout_3__2__2), .QB (\$dummy [50]), .D (
        nx3121), .CLK (CLK)) ;
    ao32 ix3122 (.Y (nx3121), .A0 (nx8064), .A1 (WindowDout_4__2__2), .A2 (
         WindowWR), .B0 (WindowDout_3__2__2), .B1 (nx8166)) ;
    dff L0_3_L1_2_Wij_reg_Dout_3 (.Q (WindowDout_3__2__3), .QB (\$dummy [51]), .D (
        nx3131), .CLK (CLK)) ;
    ao32 ix3132 (.Y (nx3131), .A0 (nx8064), .A1 (WindowDout_4__2__3), .A2 (
         WindowWR), .B0 (WindowDout_3__2__3), .B1 (nx8166)) ;
    dff L0_3_L1_2_Wij_reg_Dout_4 (.Q (WindowDout_3__2__4), .QB (\$dummy [52]), .D (
        nx3141), .CLK (CLK)) ;
    ao32 ix3142 (.Y (nx3141), .A0 (nx8064), .A1 (WindowDout_4__2__4), .A2 (
         WindowWR), .B0 (WindowDout_3__2__4), .B1 (nx8168)) ;
    dff L0_3_L1_2_Wij_reg_Dout_5 (.Q (WindowDout_3__2__5), .QB (\$dummy [53]), .D (
        nx3151), .CLK (CLK)) ;
    ao32 ix3152 (.Y (nx3151), .A0 (nx8064), .A1 (WindowDout_4__2__5), .A2 (
         WindowWR), .B0 (WindowDout_3__2__5), .B1 (nx8168)) ;
    dff L0_3_L1_2_Wij_reg_Dout_6 (.Q (WindowDout_3__2__6), .QB (\$dummy [54]), .D (
        nx3161), .CLK (CLK)) ;
    ao32 ix3162 (.Y (nx3161), .A0 (nx8064), .A1 (WindowDout_4__2__6), .A2 (
         WindowWR), .B0 (WindowDout_3__2__6), .B1 (nx8168)) ;
    dff L0_3_L1_2_Wij_reg_Dout_7 (.Q (WindowDout_3__2__7), .QB (\$dummy [55]), .D (
        nx3171), .CLK (CLK)) ;
    ao32 ix3172 (.Y (nx3171), .A0 (nx8064), .A1 (WindowDout_4__2__7), .A2 (
         WindowWR), .B0 (WindowDout_3__2__7), .B1 (nx8168)) ;
    dff L0_3_L1_1_Wij_reg_Dout_0 (.Q (WindowDout_3__1__0), .QB (\$dummy [56]), .D (
        nx3261), .CLK (CLK)) ;
    ao32 ix3262 (.Y (nx3261), .A0 (nx8064), .A1 (WindowDout_4__1__0), .A2 (
         WindowWR), .B0 (WindowDout_3__1__0), .B1 (nx8168)) ;
    dff L0_3_L1_1_Wij_reg_Dout_1 (.Q (WindowDout_3__1__1), .QB (\$dummy [57]), .D (
        nx3271), .CLK (CLK)) ;
    ao32 ix3272 (.Y (nx3271), .A0 (nx8066), .A1 (WindowDout_4__1__1), .A2 (
         WindowWR), .B0 (WindowDout_3__1__1), .B1 (nx8168)) ;
    dff L0_3_L1_1_Wij_reg_Dout_2 (.Q (WindowDout_3__1__2), .QB (\$dummy [58]), .D (
        nx3281), .CLK (CLK)) ;
    ao32 ix3282 (.Y (nx3281), .A0 (nx8066), .A1 (WindowDout_4__1__2), .A2 (
         WindowWR), .B0 (WindowDout_3__1__2), .B1 (nx8168)) ;
    dff L0_3_L1_1_Wij_reg_Dout_3 (.Q (WindowDout_3__1__3), .QB (\$dummy [59]), .D (
        nx3291), .CLK (CLK)) ;
    ao32 ix3292 (.Y (nx3291), .A0 (nx8066), .A1 (WindowDout_4__1__3), .A2 (
         WindowWR), .B0 (WindowDout_3__1__3), .B1 (nx8170)) ;
    dff L0_3_L1_1_Wij_reg_Dout_4 (.Q (WindowDout_3__1__4), .QB (\$dummy [60]), .D (
        nx3301), .CLK (CLK)) ;
    ao32 ix3302 (.Y (nx3301), .A0 (nx8066), .A1 (WindowDout_4__1__4), .A2 (
         WindowWR), .B0 (WindowDout_3__1__4), .B1 (nx8170)) ;
    dff L0_3_L1_1_Wij_reg_Dout_5 (.Q (WindowDout_3__1__5), .QB (\$dummy [61]), .D (
        nx3311), .CLK (CLK)) ;
    ao32 ix3312 (.Y (nx3311), .A0 (nx8066), .A1 (WindowDout_4__1__5), .A2 (
         WindowWR), .B0 (WindowDout_3__1__5), .B1 (nx8170)) ;
    dff L0_3_L1_1_Wij_reg_Dout_6 (.Q (WindowDout_3__1__6), .QB (\$dummy [62]), .D (
        nx3321), .CLK (CLK)) ;
    ao32 ix3322 (.Y (nx3321), .A0 (nx8066), .A1 (WindowDout_4__1__6), .A2 (
         WindowWR), .B0 (WindowDout_3__1__6), .B1 (nx8170)) ;
    dff L0_3_L1_1_Wij_reg_Dout_7 (.Q (WindowDout_3__1__7), .QB (\$dummy [63]), .D (
        nx3331), .CLK (CLK)) ;
    ao32 ix3332 (.Y (nx3331), .A0 (nx8066), .A1 (WindowDout_4__1__7), .A2 (
         WindowWR), .B0 (WindowDout_3__1__7), .B1 (nx8170)) ;
    dff L0_3_L1_0_Wij_reg_Dout_0 (.Q (WindowDout_3__0__0), .QB (\$dummy [64]), .D (
        nx3421), .CLK (CLK)) ;
    ao32 ix3422 (.Y (nx3421), .A0 (nx8068), .A1 (WindowDout_4__0__0), .A2 (
         WindowWR), .B0 (WindowDout_3__0__0), .B1 (nx8170)) ;
    dff L0_3_L1_0_Wij_reg_Dout_1 (.Q (WindowDout_3__0__1), .QB (\$dummy [65]), .D (
        nx3431), .CLK (CLK)) ;
    ao32 ix3432 (.Y (nx3431), .A0 (nx8068), .A1 (WindowDout_4__0__1), .A2 (
         WindowWR), .B0 (WindowDout_3__0__1), .B1 (nx8170)) ;
    dff L0_3_L1_0_Wij_reg_Dout_2 (.Q (WindowDout_3__0__2), .QB (\$dummy [66]), .D (
        nx3441), .CLK (CLK)) ;
    ao32 ix3442 (.Y (nx3441), .A0 (nx8068), .A1 (WindowDout_4__0__2), .A2 (
         WindowWR), .B0 (WindowDout_3__0__2), .B1 (nx8172)) ;
    dff L0_3_L1_0_Wij_reg_Dout_3 (.Q (WindowDout_3__0__3), .QB (\$dummy [67]), .D (
        nx3451), .CLK (CLK)) ;
    ao32 ix3452 (.Y (nx3451), .A0 (nx8068), .A1 (WindowDout_4__0__3), .A2 (
         WindowWR), .B0 (WindowDout_3__0__3), .B1 (nx8172)) ;
    dff L0_3_L1_0_Wij_reg_Dout_4 (.Q (WindowDout_3__0__4), .QB (\$dummy [68]), .D (
        nx3461), .CLK (CLK)) ;
    ao32 ix3462 (.Y (nx3461), .A0 (nx8068), .A1 (WindowDout_4__0__4), .A2 (
         WindowWR), .B0 (WindowDout_3__0__4), .B1 (nx8172)) ;
    dff L0_3_L1_0_Wij_reg_Dout_5 (.Q (WindowDout_3__0__5), .QB (\$dummy [69]), .D (
        nx3471), .CLK (CLK)) ;
    ao32 ix3472 (.Y (nx3471), .A0 (nx8068), .A1 (WindowDout_4__0__5), .A2 (
         WindowWR), .B0 (WindowDout_3__0__5), .B1 (nx8172)) ;
    dff L0_3_L1_0_Wij_reg_Dout_6 (.Q (WindowDout_3__0__6), .QB (\$dummy [70]), .D (
        nx3481), .CLK (CLK)) ;
    ao32 ix3482 (.Y (nx3481), .A0 (nx8068), .A1 (WindowDout_4__0__6), .A2 (
         WindowWR), .B0 (WindowDout_3__0__6), .B1 (nx8172)) ;
    dff L0_3_L1_0_Wij_reg_Dout_7 (.Q (WindowDout_3__0__7), .QB (\$dummy [71]), .D (
        nx3491), .CLK (CLK)) ;
    ao32 ix3492 (.Y (nx3491), .A0 (nx8070), .A1 (WindowDout_4__0__7), .A2 (
         WindowWR), .B0 (WindowDout_3__0__7), .B1 (nx8172)) ;
    oai21 ix3582 (.Y (nx3581), .A0 (nx6318), .A1 (nx7918), .B0 (nx6320)) ;
    dff L0_2_L1_4_Wij_reg_Dout_0 (.Q (WindowDout_2__4__0), .QB (nx6318), .D (
        nx3581), .CLK (CLK)) ;
    oai21 ix3592 (.Y (nx3591), .A0 (nx6324), .A1 (nx7918), .B0 (nx6326)) ;
    dff L0_2_L1_4_Wij_reg_Dout_1 (.Q (WindowDout_2__4__1), .QB (nx6324), .D (
        nx3591), .CLK (CLK)) ;
    oai21 ix3602 (.Y (nx3601), .A0 (nx6330), .A1 (nx7920), .B0 (nx6332)) ;
    dff L0_2_L1_4_Wij_reg_Dout_2 (.Q (WindowDout_2__4__2), .QB (nx6330), .D (
        nx3601), .CLK (CLK)) ;
    oai21 ix3612 (.Y (nx3611), .A0 (nx6336), .A1 (nx7920), .B0 (nx6338)) ;
    dff L0_2_L1_4_Wij_reg_Dout_3 (.Q (WindowDout_2__4__3), .QB (nx6336), .D (
        nx3611), .CLK (CLK)) ;
    oai21 ix3622 (.Y (nx3621), .A0 (nx6342), .A1 (nx7920), .B0 (nx6344)) ;
    dff L0_2_L1_4_Wij_reg_Dout_4 (.Q (WindowDout_2__4__4), .QB (nx6342), .D (
        nx3621), .CLK (CLK)) ;
    oai21 ix3632 (.Y (nx3631), .A0 (nx6348), .A1 (nx7922), .B0 (nx6350)) ;
    dff L0_2_L1_4_Wij_reg_Dout_5 (.Q (WindowDout_2__4__5), .QB (nx6348), .D (
        nx3631), .CLK (CLK)) ;
    oai21 ix3642 (.Y (nx3641), .A0 (nx6354), .A1 (nx7922), .B0 (nx6356)) ;
    dff L0_2_L1_4_Wij_reg_Dout_6 (.Q (WindowDout_2__4__6), .QB (nx6354), .D (
        nx3641), .CLK (CLK)) ;
    oai21 ix3652 (.Y (nx3651), .A0 (nx6360), .A1 (nx7922), .B0 (nx6362)) ;
    dff L0_2_L1_4_Wij_reg_Dout_7 (.Q (WindowDout_2__4__7), .QB (nx6360), .D (
        nx3651), .CLK (CLK)) ;
    oai21 ix3742 (.Y (nx3741), .A0 (nx6366), .A1 (nx7922), .B0 (nx6368)) ;
    dff L0_2_L1_3_Wij_reg_Dout_0 (.Q (WindowDout_2__3__0), .QB (nx6366), .D (
        nx3741), .CLK (CLK)) ;
    oai21 ix3752 (.Y (nx3751), .A0 (nx6372), .A1 (nx7924), .B0 (nx6374)) ;
    dff L0_2_L1_3_Wij_reg_Dout_1 (.Q (WindowDout_2__3__1), .QB (nx6372), .D (
        nx3751), .CLK (CLK)) ;
    oai21 ix3762 (.Y (nx3761), .A0 (nx6378), .A1 (nx7924), .B0 (nx6380)) ;
    dff L0_2_L1_3_Wij_reg_Dout_2 (.Q (WindowDout_2__3__2), .QB (nx6378), .D (
        nx3761), .CLK (CLK)) ;
    oai21 ix3772 (.Y (nx3771), .A0 (nx6384), .A1 (nx7924), .B0 (nx6386)) ;
    dff L0_2_L1_3_Wij_reg_Dout_3 (.Q (WindowDout_2__3__3), .QB (nx6384), .D (
        nx3771), .CLK (CLK)) ;
    oai21 ix3782 (.Y (nx3781), .A0 (nx6390), .A1 (nx7926), .B0 (nx6392)) ;
    dff L0_2_L1_3_Wij_reg_Dout_4 (.Q (WindowDout_2__3__4), .QB (nx6390), .D (
        nx3781), .CLK (CLK)) ;
    oai21 ix3792 (.Y (nx3791), .A0 (nx6396), .A1 (nx7926), .B0 (nx6398)) ;
    dff L0_2_L1_3_Wij_reg_Dout_5 (.Q (WindowDout_2__3__5), .QB (nx6396), .D (
        nx3791), .CLK (CLK)) ;
    oai21 ix3802 (.Y (nx3801), .A0 (nx6402), .A1 (nx7926), .B0 (nx6404)) ;
    dff L0_2_L1_3_Wij_reg_Dout_6 (.Q (WindowDout_2__3__6), .QB (nx6402), .D (
        nx3801), .CLK (CLK)) ;
    oai21 ix3812 (.Y (nx3811), .A0 (nx6408), .A1 (nx7926), .B0 (nx6410)) ;
    dff L0_2_L1_3_Wij_reg_Dout_7 (.Q (WindowDout_2__3__7), .QB (nx6408), .D (
        nx3811), .CLK (CLK)) ;
    dff L0_2_L1_2_Wij_reg_Dout_0 (.Q (WindowDout_2__2__0), .QB (\$dummy [72]), .D (
        nx3901), .CLK (CLK)) ;
    ao32 ix3902 (.Y (nx3901), .A0 (nx8074), .A1 (WindowDout_3__2__0), .A2 (
         WindowWR), .B0 (WindowDout_2__2__0), .B1 (nx8172)) ;
    dff L0_2_L1_2_Wij_reg_Dout_1 (.Q (WindowDout_2__2__1), .QB (\$dummy [73]), .D (
        nx3911), .CLK (CLK)) ;
    ao32 ix3912 (.Y (nx3911), .A0 (nx8074), .A1 (WindowDout_3__2__1), .A2 (
         WindowWR), .B0 (WindowDout_2__2__1), .B1 (nx8174)) ;
    dff L0_2_L1_2_Wij_reg_Dout_2 (.Q (WindowDout_2__2__2), .QB (\$dummy [74]), .D (
        nx3921), .CLK (CLK)) ;
    ao32 ix3922 (.Y (nx3921), .A0 (nx8074), .A1 (WindowDout_3__2__2), .A2 (
         WindowWR), .B0 (WindowDout_2__2__2), .B1 (nx8174)) ;
    dff L0_2_L1_2_Wij_reg_Dout_3 (.Q (WindowDout_2__2__3), .QB (\$dummy [75]), .D (
        nx3931), .CLK (CLK)) ;
    ao32 ix3932 (.Y (nx3931), .A0 (nx8074), .A1 (WindowDout_3__2__3), .A2 (
         WindowWR), .B0 (WindowDout_2__2__3), .B1 (nx8174)) ;
    dff L0_2_L1_2_Wij_reg_Dout_4 (.Q (WindowDout_2__2__4), .QB (\$dummy [76]), .D (
        nx3941), .CLK (CLK)) ;
    ao32 ix3942 (.Y (nx3941), .A0 (nx8076), .A1 (WindowDout_3__2__4), .A2 (
         WindowWR), .B0 (WindowDout_2__2__4), .B1 (nx8174)) ;
    dff L0_2_L1_2_Wij_reg_Dout_5 (.Q (WindowDout_2__2__5), .QB (\$dummy [77]), .D (
        nx3951), .CLK (CLK)) ;
    ao32 ix3952 (.Y (nx3951), .A0 (nx8076), .A1 (WindowDout_3__2__5), .A2 (
         WindowWR), .B0 (WindowDout_2__2__5), .B1 (nx8174)) ;
    dff L0_2_L1_2_Wij_reg_Dout_6 (.Q (WindowDout_2__2__6), .QB (\$dummy [78]), .D (
        nx3961), .CLK (CLK)) ;
    ao32 ix3962 (.Y (nx3961), .A0 (nx8076), .A1 (WindowDout_3__2__6), .A2 (
         WindowWR), .B0 (WindowDout_2__2__6), .B1 (nx8174)) ;
    dff L0_2_L1_2_Wij_reg_Dout_7 (.Q (WindowDout_2__2__7), .QB (\$dummy [79]), .D (
        nx3971), .CLK (CLK)) ;
    ao32 ix3972 (.Y (nx3971), .A0 (nx8076), .A1 (WindowDout_3__2__7), .A2 (
         WindowWR), .B0 (WindowDout_2__2__7), .B1 (nx8174)) ;
    dff L0_2_L1_1_Wij_reg_Dout_0 (.Q (WindowDout_2__1__0), .QB (\$dummy [80]), .D (
        nx4061), .CLK (CLK)) ;
    ao32 ix4062 (.Y (nx4061), .A0 (nx8076), .A1 (WindowDout_3__1__0), .A2 (
         WindowWR), .B0 (WindowDout_2__1__0), .B1 (nx8176)) ;
    dff L0_2_L1_1_Wij_reg_Dout_1 (.Q (WindowDout_2__1__1), .QB (\$dummy [81]), .D (
        nx4071), .CLK (CLK)) ;
    ao32 ix4072 (.Y (nx4071), .A0 (nx8076), .A1 (WindowDout_3__1__1), .A2 (
         WindowWR), .B0 (WindowDout_2__1__1), .B1 (nx8176)) ;
    dff L0_2_L1_1_Wij_reg_Dout_2 (.Q (WindowDout_2__1__2), .QB (\$dummy [82]), .D (
        nx4081), .CLK (CLK)) ;
    ao32 ix4082 (.Y (nx4081), .A0 (nx8076), .A1 (WindowDout_3__1__2), .A2 (
         WindowWR), .B0 (WindowDout_2__1__2), .B1 (nx8176)) ;
    dff L0_2_L1_1_Wij_reg_Dout_3 (.Q (WindowDout_2__1__3), .QB (\$dummy [83]), .D (
        nx4091), .CLK (CLK)) ;
    ao32 ix4092 (.Y (nx4091), .A0 (nx8078), .A1 (WindowDout_3__1__3), .A2 (
         WindowWR), .B0 (WindowDout_2__1__3), .B1 (nx8176)) ;
    dff L0_2_L1_1_Wij_reg_Dout_4 (.Q (WindowDout_2__1__4), .QB (\$dummy [84]), .D (
        nx4101), .CLK (CLK)) ;
    ao32 ix4102 (.Y (nx4101), .A0 (nx8078), .A1 (WindowDout_3__1__4), .A2 (
         WindowWR), .B0 (WindowDout_2__1__4), .B1 (nx8176)) ;
    dff L0_2_L1_1_Wij_reg_Dout_5 (.Q (WindowDout_2__1__5), .QB (\$dummy [85]), .D (
        nx4111), .CLK (CLK)) ;
    ao32 ix4112 (.Y (nx4111), .A0 (nx8078), .A1 (WindowDout_3__1__5), .A2 (
         WindowWR), .B0 (WindowDout_2__1__5), .B1 (nx8176)) ;
    dff L0_2_L1_1_Wij_reg_Dout_6 (.Q (WindowDout_2__1__6), .QB (\$dummy [86]), .D (
        nx4121), .CLK (CLK)) ;
    ao32 ix4122 (.Y (nx4121), .A0 (nx8078), .A1 (WindowDout_3__1__6), .A2 (
         WindowWR), .B0 (WindowDout_2__1__6), .B1 (nx8176)) ;
    dff L0_2_L1_1_Wij_reg_Dout_7 (.Q (WindowDout_2__1__7), .QB (\$dummy [87]), .D (
        nx4131), .CLK (CLK)) ;
    ao32 ix4132 (.Y (nx4131), .A0 (nx8078), .A1 (WindowDout_3__1__7), .A2 (
         WindowWR), .B0 (WindowDout_2__1__7), .B1 (nx8178)) ;
    dff L0_2_L1_0_Wij_reg_Dout_0 (.Q (WindowDout_2__0__0), .QB (\$dummy [88]), .D (
        nx4221), .CLK (CLK)) ;
    ao32 ix4222 (.Y (nx4221), .A0 (nx8078), .A1 (WindowDout_3__0__0), .A2 (
         WindowWR), .B0 (WindowDout_2__0__0), .B1 (nx8178)) ;
    dff L0_2_L1_0_Wij_reg_Dout_1 (.Q (WindowDout_2__0__1), .QB (\$dummy [89]), .D (
        nx4231), .CLK (CLK)) ;
    ao32 ix4232 (.Y (nx4231), .A0 (nx8078), .A1 (WindowDout_3__0__1), .A2 (
         WindowWR), .B0 (WindowDout_2__0__1), .B1 (nx8178)) ;
    dff L0_2_L1_0_Wij_reg_Dout_2 (.Q (WindowDout_2__0__2), .QB (\$dummy [90]), .D (
        nx4241), .CLK (CLK)) ;
    ao32 ix4242 (.Y (nx4241), .A0 (nx8080), .A1 (WindowDout_3__0__2), .A2 (
         WindowWR), .B0 (WindowDout_2__0__2), .B1 (nx8178)) ;
    dff L0_2_L1_0_Wij_reg_Dout_3 (.Q (WindowDout_2__0__3), .QB (\$dummy [91]), .D (
        nx4251), .CLK (CLK)) ;
    ao32 ix4252 (.Y (nx4251), .A0 (nx8080), .A1 (WindowDout_3__0__3), .A2 (
         WindowWR), .B0 (WindowDout_2__0__3), .B1 (nx8178)) ;
    dff L0_2_L1_0_Wij_reg_Dout_4 (.Q (WindowDout_2__0__4), .QB (\$dummy [92]), .D (
        nx4261), .CLK (CLK)) ;
    ao32 ix4262 (.Y (nx4261), .A0 (nx8080), .A1 (WindowDout_3__0__4), .A2 (
         WindowWR), .B0 (WindowDout_2__0__4), .B1 (nx8178)) ;
    dff L0_2_L1_0_Wij_reg_Dout_5 (.Q (WindowDout_2__0__5), .QB (\$dummy [93]), .D (
        nx4271), .CLK (CLK)) ;
    ao32 ix4272 (.Y (nx4271), .A0 (nx8080), .A1 (WindowDout_3__0__5), .A2 (
         WindowWR), .B0 (WindowDout_2__0__5), .B1 (nx8178)) ;
    dff L0_2_L1_0_Wij_reg_Dout_6 (.Q (WindowDout_2__0__6), .QB (\$dummy [94]), .D (
        nx4281), .CLK (CLK)) ;
    ao32 ix4282 (.Y (nx4281), .A0 (nx8080), .A1 (WindowDout_3__0__6), .A2 (
         WindowWR), .B0 (WindowDout_2__0__6), .B1 (nx8180)) ;
    dff L0_2_L1_0_Wij_reg_Dout_7 (.Q (WindowDout_2__0__7), .QB (\$dummy [95]), .D (
        nx4291), .CLK (CLK)) ;
    ao32 ix4292 (.Y (nx4291), .A0 (nx8080), .A1 (WindowDout_3__0__7), .A2 (
         WindowWR), .B0 (WindowDout_2__0__7), .B1 (nx8180)) ;
    oai21 ix4382 (.Y (nx4381), .A0 (nx6486), .A1 (nx7928), .B0 (nx6488)) ;
    dff L0_1_L1_4_Wij_reg_Dout_0 (.Q (WindowDout_1__4__0), .QB (nx6486), .D (
        nx4381), .CLK (CLK)) ;
    oai21 ix4392 (.Y (nx4391), .A0 (nx6492), .A1 (nx7928), .B0 (nx6494)) ;
    dff L0_1_L1_4_Wij_reg_Dout_1 (.Q (WindowDout_1__4__1), .QB (nx6492), .D (
        nx4391), .CLK (CLK)) ;
    oai21 ix4402 (.Y (nx4401), .A0 (nx6498), .A1 (nx7928), .B0 (nx6500)) ;
    dff L0_1_L1_4_Wij_reg_Dout_2 (.Q (WindowDout_1__4__2), .QB (nx6498), .D (
        nx4401), .CLK (CLK)) ;
    oai21 ix4412 (.Y (nx4411), .A0 (nx6504), .A1 (nx7930), .B0 (nx6506)) ;
    dff L0_1_L1_4_Wij_reg_Dout_3 (.Q (WindowDout_1__4__3), .QB (nx6504), .D (
        nx4411), .CLK (CLK)) ;
    oai21 ix4422 (.Y (nx4421), .A0 (nx6510), .A1 (nx7930), .B0 (nx6512)) ;
    dff L0_1_L1_4_Wij_reg_Dout_4 (.Q (WindowDout_1__4__4), .QB (nx6510), .D (
        nx4421), .CLK (CLK)) ;
    oai21 ix4432 (.Y (nx4431), .A0 (nx6516), .A1 (nx7930), .B0 (nx6518)) ;
    dff L0_1_L1_4_Wij_reg_Dout_5 (.Q (WindowDout_1__4__5), .QB (nx6516), .D (
        nx4431), .CLK (CLK)) ;
    oai21 ix4442 (.Y (nx4441), .A0 (nx6522), .A1 (nx7930), .B0 (nx6524)) ;
    dff L0_1_L1_4_Wij_reg_Dout_6 (.Q (WindowDout_1__4__6), .QB (nx6522), .D (
        nx4441), .CLK (CLK)) ;
    oai21 ix4452 (.Y (nx4451), .A0 (nx6528), .A1 (nx7932), .B0 (nx6530)) ;
    dff L0_1_L1_4_Wij_reg_Dout_7 (.Q (WindowDout_1__4__7), .QB (nx6528), .D (
        nx4451), .CLK (CLK)) ;
    oai21 ix4702 (.Y (nx4701), .A0 (nx6534), .A1 (nx7932), .B0 (nx6536)) ;
    dff L0_1_L1_3_Wij_reg_Dout_0 (.Q (WindowDout_1__3__0), .QB (nx6534), .D (
        nx4701), .CLK (CLK)) ;
    oai21 ix4712 (.Y (nx4711), .A0 (nx6540), .A1 (nx7932), .B0 (nx6542)) ;
    dff L0_1_L1_3_Wij_reg_Dout_1 (.Q (WindowDout_1__3__1), .QB (nx6540), .D (
        nx4711), .CLK (CLK)) ;
    oai21 ix4722 (.Y (nx4721), .A0 (nx6546), .A1 (nx7934), .B0 (nx6548)) ;
    dff L0_1_L1_3_Wij_reg_Dout_2 (.Q (WindowDout_1__3__2), .QB (nx6546), .D (
        nx4721), .CLK (CLK)) ;
    oai21 ix4732 (.Y (nx4731), .A0 (nx6552), .A1 (nx7934), .B0 (nx6554)) ;
    dff L0_1_L1_3_Wij_reg_Dout_3 (.Q (WindowDout_1__3__3), .QB (nx6552), .D (
        nx4731), .CLK (CLK)) ;
    oai21 ix4742 (.Y (nx4741), .A0 (nx6558), .A1 (nx7934), .B0 (nx6560)) ;
    dff L0_1_L1_3_Wij_reg_Dout_4 (.Q (WindowDout_1__3__4), .QB (nx6558), .D (
        nx4741), .CLK (CLK)) ;
    oai21 ix4752 (.Y (nx4751), .A0 (nx6564), .A1 (nx7934), .B0 (nx6566)) ;
    dff L0_1_L1_3_Wij_reg_Dout_5 (.Q (WindowDout_1__3__5), .QB (nx6564), .D (
        nx4751), .CLK (CLK)) ;
    oai21 ix4762 (.Y (nx4761), .A0 (nx6570), .A1 (nx7936), .B0 (nx6572)) ;
    dff L0_1_L1_3_Wij_reg_Dout_6 (.Q (WindowDout_1__3__6), .QB (nx6570), .D (
        nx4761), .CLK (CLK)) ;
    oai21 ix4772 (.Y (nx4771), .A0 (nx6576), .A1 (nx7936), .B0 (nx6578)) ;
    dff L0_1_L1_3_Wij_reg_Dout_7 (.Q (WindowDout_1__3__7), .QB (nx6576), .D (
        nx4771), .CLK (CLK)) ;
    oai21 ix5022 (.Y (nx5021), .A0 (nx6582), .A1 (nx7936), .B0 (nx6584)) ;
    dff L0_1_L1_2_Wij_reg_Dout_0 (.Q (WindowDout_1__2__0), .QB (nx6582), .D (
        nx5021), .CLK (CLK)) ;
    nand03 ix6585 (.Y (nx6584), .A0 (nx8086), .A1 (WindowDout_2__2__0), .A2 (
           nx7936)) ;
    oai21 ix5032 (.Y (nx5031), .A0 (nx6588), .A1 (nx7938), .B0 (nx6590)) ;
    dff L0_1_L1_2_Wij_reg_Dout_1 (.Q (WindowDout_1__2__1), .QB (nx6588), .D (
        nx5031), .CLK (CLK)) ;
    nand03 ix6591 (.Y (nx6590), .A0 (nx8086), .A1 (WindowDout_2__2__1), .A2 (
           nx7938)) ;
    oai21 ix5042 (.Y (nx5041), .A0 (nx6594), .A1 (nx7938), .B0 (nx6596)) ;
    dff L0_1_L1_2_Wij_reg_Dout_2 (.Q (WindowDout_1__2__2), .QB (nx6594), .D (
        nx5041), .CLK (CLK)) ;
    nand03 ix6597 (.Y (nx6596), .A0 (nx8086), .A1 (WindowDout_2__2__2), .A2 (
           nx7938)) ;
    oai21 ix5052 (.Y (nx5051), .A0 (nx6600), .A1 (nx7938), .B0 (nx6602)) ;
    dff L0_1_L1_2_Wij_reg_Dout_3 (.Q (WindowDout_1__2__3), .QB (nx6600), .D (
        nx5051), .CLK (CLK)) ;
    nand03 ix6603 (.Y (nx6602), .A0 (nx8086), .A1 (WindowDout_2__2__3), .A2 (
           nx7938)) ;
    oai21 ix5062 (.Y (nx5061), .A0 (nx6606), .A1 (nx7938), .B0 (nx6608)) ;
    dff L0_1_L1_2_Wij_reg_Dout_4 (.Q (WindowDout_1__2__4), .QB (nx6606), .D (
        nx5061), .CLK (CLK)) ;
    nand03 ix6609 (.Y (nx6608), .A0 (nx8086), .A1 (WindowDout_2__2__4), .A2 (
           nx7940)) ;
    oai21 ix5072 (.Y (nx5071), .A0 (nx6612), .A1 (nx7940), .B0 (nx6614)) ;
    dff L0_1_L1_2_Wij_reg_Dout_5 (.Q (WindowDout_1__2__5), .QB (nx6612), .D (
        nx5071), .CLK (CLK)) ;
    nand03 ix6615 (.Y (nx6614), .A0 (nx8086), .A1 (WindowDout_2__2__5), .A2 (
           nx7940)) ;
    oai21 ix5082 (.Y (nx5081), .A0 (nx6618), .A1 (nx7940), .B0 (nx6620)) ;
    dff L0_1_L1_2_Wij_reg_Dout_6 (.Q (WindowDout_1__2__6), .QB (nx6618), .D (
        nx5081), .CLK (CLK)) ;
    nand03 ix6621 (.Y (nx6620), .A0 (nx8088), .A1 (WindowDout_2__2__6), .A2 (
           nx7940)) ;
    oai21 ix5092 (.Y (nx5091), .A0 (nx6624), .A1 (nx7940), .B0 (nx6626)) ;
    dff L0_1_L1_2_Wij_reg_Dout_7 (.Q (WindowDout_1__2__7), .QB (nx6624), .D (
        nx5091), .CLK (CLK)) ;
    nand03 ix6627 (.Y (nx6626), .A0 (nx8088), .A1 (WindowDout_2__2__7), .A2 (
           nx7940)) ;
    oai21 ix5342 (.Y (nx5341), .A0 (nx6630), .A1 (nx7942), .B0 (nx6632)) ;
    dff L0_1_L1_1_Wij_reg_Dout_0 (.Q (WindowDout_1__1__0), .QB (nx6630), .D (
        nx5341), .CLK (CLK)) ;
    nand03 ix6633 (.Y (nx6632), .A0 (nx8088), .A1 (WindowDout_2__1__0), .A2 (
           nx7942)) ;
    oai21 ix5352 (.Y (nx5351), .A0 (nx6636), .A1 (nx7942), .B0 (nx6638)) ;
    dff L0_1_L1_1_Wij_reg_Dout_1 (.Q (WindowDout_1__1__1), .QB (nx6636), .D (
        nx5351), .CLK (CLK)) ;
    nand03 ix6639 (.Y (nx6638), .A0 (nx8088), .A1 (WindowDout_2__1__1), .A2 (
           nx7942)) ;
    oai21 ix5362 (.Y (nx5361), .A0 (nx6642), .A1 (nx7942), .B0 (nx6644)) ;
    dff L0_1_L1_1_Wij_reg_Dout_2 (.Q (WindowDout_1__1__2), .QB (nx6642), .D (
        nx5361), .CLK (CLK)) ;
    nand03 ix6645 (.Y (nx6644), .A0 (nx8088), .A1 (WindowDout_2__1__2), .A2 (
           nx7942)) ;
    oai21 ix5372 (.Y (nx5371), .A0 (nx6648), .A1 (nx7942), .B0 (nx6650)) ;
    dff L0_1_L1_1_Wij_reg_Dout_3 (.Q (WindowDout_1__1__3), .QB (nx6648), .D (
        nx5371), .CLK (CLK)) ;
    nand03 ix6651 (.Y (nx6650), .A0 (nx8088), .A1 (WindowDout_2__1__3), .A2 (
           nx7944)) ;
    oai21 ix5382 (.Y (nx5381), .A0 (nx6654), .A1 (nx7944), .B0 (nx6656)) ;
    dff L0_1_L1_1_Wij_reg_Dout_4 (.Q (WindowDout_1__1__4), .QB (nx6654), .D (
        nx5381), .CLK (CLK)) ;
    nand03 ix6657 (.Y (nx6656), .A0 (nx8088), .A1 (WindowDout_2__1__4), .A2 (
           nx7944)) ;
    oai21 ix5392 (.Y (nx5391), .A0 (nx6660), .A1 (nx7944), .B0 (nx6662)) ;
    dff L0_1_L1_1_Wij_reg_Dout_5 (.Q (WindowDout_1__1__5), .QB (nx6660), .D (
        nx5391), .CLK (CLK)) ;
    nand03 ix6663 (.Y (nx6662), .A0 (nx8090), .A1 (WindowDout_2__1__5), .A2 (
           nx7944)) ;
    oai21 ix5402 (.Y (nx5401), .A0 (nx6666), .A1 (nx7944), .B0 (nx6668)) ;
    dff L0_1_L1_1_Wij_reg_Dout_6 (.Q (WindowDout_1__1__6), .QB (nx6666), .D (
        nx5401), .CLK (CLK)) ;
    nand03 ix6669 (.Y (nx6668), .A0 (nx8090), .A1 (WindowDout_2__1__6), .A2 (
           nx7944)) ;
    oai21 ix5412 (.Y (nx5411), .A0 (nx6672), .A1 (nx7946), .B0 (nx6674)) ;
    dff L0_1_L1_1_Wij_reg_Dout_7 (.Q (WindowDout_1__1__7), .QB (nx6672), .D (
        nx5411), .CLK (CLK)) ;
    nand03 ix6675 (.Y (nx6674), .A0 (nx8090), .A1 (WindowDout_2__1__7), .A2 (
           nx7946)) ;
    oai21 ix5662 (.Y (nx5661), .A0 (nx6678), .A1 (nx7946), .B0 (nx6680)) ;
    dff L0_1_L1_0_Wij_reg_Dout_0 (.Q (WindowDout_1__0__0), .QB (nx6678), .D (
        nx5661), .CLK (CLK)) ;
    nand03 ix6681 (.Y (nx6680), .A0 (nx8090), .A1 (WindowDout_2__0__0), .A2 (
           nx7946)) ;
    oai21 ix5672 (.Y (nx5671), .A0 (nx6684), .A1 (nx7946), .B0 (nx6686)) ;
    dff L0_1_L1_0_Wij_reg_Dout_1 (.Q (WindowDout_1__0__1), .QB (nx6684), .D (
        nx5671), .CLK (CLK)) ;
    nand03 ix6687 (.Y (nx6686), .A0 (nx8090), .A1 (WindowDout_2__0__1), .A2 (
           nx7946)) ;
    oai21 ix5682 (.Y (nx5681), .A0 (nx6690), .A1 (nx7946), .B0 (nx6692)) ;
    dff L0_1_L1_0_Wij_reg_Dout_2 (.Q (WindowDout_1__0__2), .QB (nx6690), .D (
        nx5681), .CLK (CLK)) ;
    nand03 ix6693 (.Y (nx6692), .A0 (nx8090), .A1 (WindowDout_2__0__2), .A2 (
           nx7948)) ;
    oai21 ix5692 (.Y (nx5691), .A0 (nx6696), .A1 (nx7948), .B0 (nx6698)) ;
    dff L0_1_L1_0_Wij_reg_Dout_3 (.Q (WindowDout_1__0__3), .QB (nx6696), .D (
        nx5691), .CLK (CLK)) ;
    nand03 ix6699 (.Y (nx6698), .A0 (nx8090), .A1 (WindowDout_2__0__3), .A2 (
           nx7948)) ;
    oai21 ix5702 (.Y (nx5701), .A0 (nx6702), .A1 (nx7948), .B0 (nx6704)) ;
    dff L0_1_L1_0_Wij_reg_Dout_4 (.Q (WindowDout_1__0__4), .QB (nx6702), .D (
        nx5701), .CLK (CLK)) ;
    nand03 ix6705 (.Y (nx6704), .A0 (nx8092), .A1 (WindowDout_2__0__4), .A2 (
           nx7948)) ;
    oai21 ix5712 (.Y (nx5711), .A0 (nx6708), .A1 (nx7948), .B0 (nx6710)) ;
    dff L0_1_L1_0_Wij_reg_Dout_5 (.Q (WindowDout_1__0__5), .QB (nx6708), .D (
        nx5711), .CLK (CLK)) ;
    nand03 ix6711 (.Y (nx6710), .A0 (nx8092), .A1 (WindowDout_2__0__5), .A2 (
           nx7948)) ;
    oai21 ix5722 (.Y (nx5721), .A0 (nx6714), .A1 (nx7950), .B0 (nx6716)) ;
    dff L0_1_L1_0_Wij_reg_Dout_6 (.Q (WindowDout_1__0__6), .QB (nx6714), .D (
        nx5721), .CLK (CLK)) ;
    nand03 ix6717 (.Y (nx6716), .A0 (nx8092), .A1 (WindowDout_2__0__6), .A2 (
           nx7950)) ;
    oai21 ix5732 (.Y (nx5731), .A0 (nx6720), .A1 (nx7950), .B0 (nx6722)) ;
    dff L0_1_L1_0_Wij_reg_Dout_7 (.Q (WindowDout_1__0__7), .QB (nx6720), .D (
        nx5731), .CLK (CLK)) ;
    nand03 ix6723 (.Y (nx6722), .A0 (nx8092), .A1 (WindowDout_2__0__7), .A2 (
           nx7950)) ;
    oai21 ix4462 (.Y (nx4461), .A0 (nx6726), .A1 (nx7950), .B0 (nx6728)) ;
    dff L0_0_L1_4_Wij_reg_Dout_0 (.Q (WindowDout_0__4__0), .QB (nx6726), .D (
        nx4461), .CLK (CLK)) ;
    oai21 ix4472 (.Y (nx4471), .A0 (nx6732), .A1 (nx7950), .B0 (nx6734)) ;
    dff L0_0_L1_4_Wij_reg_Dout_1 (.Q (WindowDout_0__4__1), .QB (nx6732), .D (
        nx4471), .CLK (CLK)) ;
    oai21 ix4482 (.Y (nx4481), .A0 (nx6738), .A1 (nx7952), .B0 (nx6740)) ;
    dff L0_0_L1_4_Wij_reg_Dout_2 (.Q (WindowDout_0__4__2), .QB (nx6738), .D (
        nx4481), .CLK (CLK)) ;
    oai21 ix4492 (.Y (nx4491), .A0 (nx6744), .A1 (nx7952), .B0 (nx6746)) ;
    dff L0_0_L1_4_Wij_reg_Dout_3 (.Q (WindowDout_0__4__3), .QB (nx6744), .D (
        nx4491), .CLK (CLK)) ;
    oai21 ix4502 (.Y (nx4501), .A0 (nx6750), .A1 (nx7952), .B0 (nx6752)) ;
    dff L0_0_L1_4_Wij_reg_Dout_4 (.Q (WindowDout_0__4__4), .QB (nx6750), .D (
        nx4501), .CLK (CLK)) ;
    oai21 ix4512 (.Y (nx4511), .A0 (nx6756), .A1 (nx7954), .B0 (nx6758)) ;
    dff L0_0_L1_4_Wij_reg_Dout_5 (.Q (WindowDout_0__4__5), .QB (nx6756), .D (
        nx4511), .CLK (CLK)) ;
    oai21 ix4522 (.Y (nx4521), .A0 (nx6762), .A1 (nx7954), .B0 (nx6764)) ;
    dff L0_0_L1_4_Wij_reg_Dout_6 (.Q (WindowDout_0__4__6), .QB (nx6762), .D (
        nx4521), .CLK (CLK)) ;
    oai21 ix4532 (.Y (nx4531), .A0 (nx6768), .A1 (nx7954), .B0 (nx6770)) ;
    dff L0_0_L1_4_Wij_reg_Dout_7 (.Q (WindowDout_0__4__7), .QB (nx6768), .D (
        nx4531), .CLK (CLK)) ;
    oai21 ix4782 (.Y (nx4781), .A0 (nx6774), .A1 (nx7954), .B0 (nx6776)) ;
    dff L0_0_L1_3_Wij_reg_Dout_0 (.Q (WindowDout_0__3__0), .QB (nx6774), .D (
        nx4781), .CLK (CLK)) ;
    oai21 ix4792 (.Y (nx4791), .A0 (nx6780), .A1 (nx7956), .B0 (nx6782)) ;
    dff L0_0_L1_3_Wij_reg_Dout_1 (.Q (WindowDout_0__3__1), .QB (nx6780), .D (
        nx4791), .CLK (CLK)) ;
    oai21 ix4802 (.Y (nx4801), .A0 (nx6786), .A1 (nx7956), .B0 (nx6788)) ;
    dff L0_0_L1_3_Wij_reg_Dout_2 (.Q (WindowDout_0__3__2), .QB (nx6786), .D (
        nx4801), .CLK (CLK)) ;
    oai21 ix4812 (.Y (nx4811), .A0 (nx6792), .A1 (nx7956), .B0 (nx6794)) ;
    dff L0_0_L1_3_Wij_reg_Dout_3 (.Q (WindowDout_0__3__3), .QB (nx6792), .D (
        nx4811), .CLK (CLK)) ;
    oai21 ix4822 (.Y (nx4821), .A0 (nx6798), .A1 (nx7958), .B0 (nx6800)) ;
    dff L0_0_L1_3_Wij_reg_Dout_4 (.Q (WindowDout_0__3__4), .QB (nx6798), .D (
        nx4821), .CLK (CLK)) ;
    oai21 ix4832 (.Y (nx4831), .A0 (nx6804), .A1 (nx7958), .B0 (nx6806)) ;
    dff L0_0_L1_3_Wij_reg_Dout_5 (.Q (WindowDout_0__3__5), .QB (nx6804), .D (
        nx4831), .CLK (CLK)) ;
    oai21 ix4842 (.Y (nx4841), .A0 (nx6810), .A1 (nx7958), .B0 (nx6812)) ;
    dff L0_0_L1_3_Wij_reg_Dout_6 (.Q (WindowDout_0__3__6), .QB (nx6810), .D (
        nx4841), .CLK (CLK)) ;
    oai21 ix4852 (.Y (nx4851), .A0 (nx6816), .A1 (nx7958), .B0 (nx6818)) ;
    dff L0_0_L1_3_Wij_reg_Dout_7 (.Q (WindowDout_0__3__7), .QB (nx6816), .D (
        nx4851), .CLK (CLK)) ;
    oai21 ix5102 (.Y (nx5101), .A0 (nx6822), .A1 (nx7960), .B0 (nx6824)) ;
    dff L0_0_L1_2_Wij_reg_Dout_0 (.Q (WindowDout_0__2__0), .QB (nx6822), .D (
        nx5101), .CLK (CLK)) ;
    oai21 ix5112 (.Y (nx5111), .A0 (nx6828), .A1 (nx7960), .B0 (nx6830)) ;
    dff L0_0_L1_2_Wij_reg_Dout_1 (.Q (WindowDout_0__2__1), .QB (nx6828), .D (
        nx5111), .CLK (CLK)) ;
    oai21 ix5122 (.Y (nx5121), .A0 (nx6834), .A1 (nx7960), .B0 (nx6836)) ;
    dff L0_0_L1_2_Wij_reg_Dout_2 (.Q (WindowDout_0__2__2), .QB (nx6834), .D (
        nx5121), .CLK (CLK)) ;
    oai21 ix5132 (.Y (nx5131), .A0 (nx6840), .A1 (nx7962), .B0 (nx6842)) ;
    dff L0_0_L1_2_Wij_reg_Dout_3 (.Q (WindowDout_0__2__3), .QB (nx6840), .D (
        nx5131), .CLK (CLK)) ;
    oai21 ix5142 (.Y (nx5141), .A0 (nx6846), .A1 (nx7962), .B0 (nx6848)) ;
    dff L0_0_L1_2_Wij_reg_Dout_4 (.Q (WindowDout_0__2__4), .QB (nx6846), .D (
        nx5141), .CLK (CLK)) ;
    oai21 ix5152 (.Y (nx5151), .A0 (nx6852), .A1 (nx7962), .B0 (nx6854)) ;
    dff L0_0_L1_2_Wij_reg_Dout_5 (.Q (WindowDout_0__2__5), .QB (nx6852), .D (
        nx5151), .CLK (CLK)) ;
    oai21 ix5162 (.Y (nx5161), .A0 (nx6858), .A1 (nx7962), .B0 (nx6860)) ;
    dff L0_0_L1_2_Wij_reg_Dout_6 (.Q (WindowDout_0__2__6), .QB (nx6858), .D (
        nx5161), .CLK (CLK)) ;
    oai21 ix5172 (.Y (nx5171), .A0 (nx6864), .A1 (nx7964), .B0 (nx6866)) ;
    dff L0_0_L1_2_Wij_reg_Dout_7 (.Q (WindowDout_0__2__7), .QB (nx6864), .D (
        nx5171), .CLK (CLK)) ;
    oai21 ix5422 (.Y (nx5421), .A0 (nx6870), .A1 (nx7964), .B0 (nx6872)) ;
    dff L0_0_L1_1_Wij_reg_Dout_0 (.Q (WindowDout_0__1__0), .QB (nx6870), .D (
        nx5421), .CLK (CLK)) ;
    oai21 ix5432 (.Y (nx5431), .A0 (nx6876), .A1 (nx7964), .B0 (nx6878)) ;
    dff L0_0_L1_1_Wij_reg_Dout_1 (.Q (WindowDout_0__1__1), .QB (nx6876), .D (
        nx5431), .CLK (CLK)) ;
    oai21 ix5442 (.Y (nx5441), .A0 (nx6882), .A1 (nx7966), .B0 (nx6884)) ;
    dff L0_0_L1_1_Wij_reg_Dout_2 (.Q (WindowDout_0__1__2), .QB (nx6882), .D (
        nx5441), .CLK (CLK)) ;
    oai21 ix5452 (.Y (nx5451), .A0 (nx6888), .A1 (nx7966), .B0 (nx6890)) ;
    dff L0_0_L1_1_Wij_reg_Dout_3 (.Q (WindowDout_0__1__3), .QB (nx6888), .D (
        nx5451), .CLK (CLK)) ;
    oai21 ix5462 (.Y (nx5461), .A0 (nx6894), .A1 (nx7966), .B0 (nx6896)) ;
    dff L0_0_L1_1_Wij_reg_Dout_4 (.Q (WindowDout_0__1__4), .QB (nx6894), .D (
        nx5461), .CLK (CLK)) ;
    oai21 ix5472 (.Y (nx5471), .A0 (nx6900), .A1 (nx7966), .B0 (nx6902)) ;
    dff L0_0_L1_1_Wij_reg_Dout_5 (.Q (WindowDout_0__1__5), .QB (nx6900), .D (
        nx5471), .CLK (CLK)) ;
    oai21 ix5482 (.Y (nx5481), .A0 (nx6906), .A1 (nx7968), .B0 (nx6908)) ;
    dff L0_0_L1_1_Wij_reg_Dout_6 (.Q (WindowDout_0__1__6), .QB (nx6906), .D (
        nx5481), .CLK (CLK)) ;
    oai21 ix5492 (.Y (nx5491), .A0 (nx6912), .A1 (nx7968), .B0 (nx6914)) ;
    dff L0_0_L1_1_Wij_reg_Dout_7 (.Q (WindowDout_0__1__7), .QB (nx6912), .D (
        nx5491), .CLK (CLK)) ;
    oai21 ix5742 (.Y (nx5741), .A0 (nx6918), .A1 (nx7968), .B0 (nx6920)) ;
    dff L0_0_L1_0_Wij_reg_Dout_0 (.Q (WindowDout_0__0__0), .QB (nx6918), .D (
        nx5741), .CLK (CLK)) ;
    oai21 ix5752 (.Y (nx5751), .A0 (nx6924), .A1 (nx7970), .B0 (nx6926)) ;
    dff L0_0_L1_0_Wij_reg_Dout_1 (.Q (WindowDout_0__0__1), .QB (nx6924), .D (
        nx5751), .CLK (CLK)) ;
    oai21 ix5762 (.Y (nx5761), .A0 (nx6930), .A1 (nx7970), .B0 (nx6932)) ;
    dff L0_0_L1_0_Wij_reg_Dout_2 (.Q (WindowDout_0__0__2), .QB (nx6930), .D (
        nx5761), .CLK (CLK)) ;
    oai21 ix5772 (.Y (nx5771), .A0 (nx6936), .A1 (nx7970), .B0 (nx6938)) ;
    dff L0_0_L1_0_Wij_reg_Dout_3 (.Q (WindowDout_0__0__3), .QB (nx6936), .D (
        nx5771), .CLK (CLK)) ;
    oai21 ix5782 (.Y (nx5781), .A0 (nx6942), .A1 (nx7970), .B0 (nx6944)) ;
    dff L0_0_L1_0_Wij_reg_Dout_4 (.Q (WindowDout_0__0__4), .QB (nx6942), .D (
        nx5781), .CLK (CLK)) ;
    oai21 ix5792 (.Y (nx5791), .A0 (nx6948), .A1 (nx7972), .B0 (nx6950)) ;
    dff L0_0_L1_0_Wij_reg_Dout_5 (.Q (WindowDout_0__0__5), .QB (nx6948), .D (
        nx5791), .CLK (CLK)) ;
    oai21 ix5802 (.Y (nx5801), .A0 (nx6954), .A1 (nx7972), .B0 (nx6956)) ;
    dff L0_0_L1_0_Wij_reg_Dout_6 (.Q (WindowDout_0__0__6), .QB (nx6954), .D (
        nx5801), .CLK (CLK)) ;
    oai21 ix5812 (.Y (nx5811), .A0 (nx6960), .A1 (nx7972), .B0 (nx6962)) ;
    dff L0_0_L1_0_Wij_reg_Dout_7 (.Q (WindowDout_0__0__7), .QB (nx6960), .D (
        nx5811), .CLK (CLK)) ;
    dff L0_4_L1_4_Fij_reg_Dout_0 (.Q (FilterDout_4__4__0), .QB (\$dummy [96]), .D (
        nx2061), .CLK (CLK)) ;
    aoi21 ix6967 (.Y (nx6966), .A0 (FilterSize), .A1 (FilterWR), .B0 (RST)) ;
    dff L0_4_L1_4_Fij_reg_Dout_1 (.Q (FilterDout_4__4__1), .QB (\$dummy [97]), .D (
        nx2071), .CLK (CLK)) ;
    dff L0_4_L1_4_Fij_reg_Dout_2 (.Q (FilterDout_4__4__2), .QB (\$dummy [98]), .D (
        nx2081), .CLK (CLK)) ;
    dff L0_4_L1_4_Fij_reg_Dout_3 (.Q (FilterDout_4__4__3), .QB (\$dummy [99]), .D (
        nx2091), .CLK (CLK)) ;
    dff L0_4_L1_4_Fij_reg_Dout_4 (.Q (FilterDout_4__4__4), .QB (\$dummy [100]), 
        .D (nx2101), .CLK (CLK)) ;
    dff L0_4_L1_4_Fij_reg_Dout_5 (.Q (FilterDout_4__4__5), .QB (\$dummy [101]), 
        .D (nx2111), .CLK (CLK)) ;
    dff L0_4_L1_4_Fij_reg_Dout_6 (.Q (FilterDout_4__4__6), .QB (\$dummy [102]), 
        .D (nx2121), .CLK (CLK)) ;
    dff L0_4_L1_4_Fij_reg_Dout_7 (.Q (FilterDout_4__4__7), .QB (\$dummy [103]), 
        .D (nx2131), .CLK (CLK)) ;
    dff L0_4_L1_3_Fij_reg_Dout_0 (.Q (FilterDout_4__3__0), .QB (\$dummy [104]), 
        .D (nx2221), .CLK (CLK)) ;
    dff L0_4_L1_3_Fij_reg_Dout_1 (.Q (FilterDout_4__3__1), .QB (\$dummy [105]), 
        .D (nx2231), .CLK (CLK)) ;
    dff L0_4_L1_3_Fij_reg_Dout_2 (.Q (FilterDout_4__3__2), .QB (\$dummy [106]), 
        .D (nx2241), .CLK (CLK)) ;
    dff L0_4_L1_3_Fij_reg_Dout_3 (.Q (FilterDout_4__3__3), .QB (\$dummy [107]), 
        .D (nx2251), .CLK (CLK)) ;
    dff L0_4_L1_3_Fij_reg_Dout_4 (.Q (FilterDout_4__3__4), .QB (\$dummy [108]), 
        .D (nx2261), .CLK (CLK)) ;
    dff L0_4_L1_3_Fij_reg_Dout_5 (.Q (FilterDout_4__3__5), .QB (\$dummy [109]), 
        .D (nx2271), .CLK (CLK)) ;
    dff L0_4_L1_3_Fij_reg_Dout_6 (.Q (FilterDout_4__3__6), .QB (\$dummy [110]), 
        .D (nx2281), .CLK (CLK)) ;
    dff L0_4_L1_3_Fij_reg_Dout_7 (.Q (FilterDout_4__3__7), .QB (\$dummy [111]), 
        .D (nx2291), .CLK (CLK)) ;
    dff L0_4_L1_2_Fij_reg_Dout_0 (.Q (FilterDout_4__2__0), .QB (\$dummy [112]), 
        .D (nx2381), .CLK (CLK)) ;
    ao32 ix2382 (.Y (nx2381), .A0 (Din[16]), .A1 (nx8104), .A2 (FilterWR), .B0 (
         FilterDout_4__2__0), .B1 (nx8198)) ;
    nor02_2x ix7017 (.Y (nx7016), .A0 (FilterWR), .A1 (RST)) ;
    dff L0_4_L1_2_Fij_reg_Dout_1 (.Q (FilterDout_4__2__1), .QB (\$dummy [113]), 
        .D (nx2391), .CLK (CLK)) ;
    ao32 ix2392 (.Y (nx2391), .A0 (Din[17]), .A1 (nx8104), .A2 (FilterWR), .B0 (
         FilterDout_4__2__1), .B1 (nx8198)) ;
    dff L0_4_L1_2_Fij_reg_Dout_2 (.Q (FilterDout_4__2__2), .QB (\$dummy [114]), 
        .D (nx2401), .CLK (CLK)) ;
    ao32 ix2402 (.Y (nx2401), .A0 (Din[18]), .A1 (nx8104), .A2 (FilterWR), .B0 (
         FilterDout_4__2__2), .B1 (nx8198)) ;
    dff L0_4_L1_2_Fij_reg_Dout_3 (.Q (FilterDout_4__2__3), .QB (\$dummy [115]), 
        .D (nx2411), .CLK (CLK)) ;
    ao32 ix2412 (.Y (nx2411), .A0 (Din[19]), .A1 (nx8104), .A2 (FilterWR), .B0 (
         FilterDout_4__2__3), .B1 (nx8198)) ;
    dff L0_4_L1_2_Fij_reg_Dout_4 (.Q (FilterDout_4__2__4), .QB (\$dummy [116]), 
        .D (nx2421), .CLK (CLK)) ;
    ao32 ix2422 (.Y (nx2421), .A0 (Din[20]), .A1 (nx8104), .A2 (FilterWR), .B0 (
         FilterDout_4__2__4), .B1 (nx8198)) ;
    dff L0_4_L1_2_Fij_reg_Dout_5 (.Q (FilterDout_4__2__5), .QB (\$dummy [117]), 
        .D (nx2431), .CLK (CLK)) ;
    ao32 ix2432 (.Y (nx2431), .A0 (Din[21]), .A1 (nx8106), .A2 (FilterWR), .B0 (
         FilterDout_4__2__5), .B1 (nx8198)) ;
    dff L0_4_L1_2_Fij_reg_Dout_6 (.Q (FilterDout_4__2__6), .QB (\$dummy [118]), 
        .D (nx2441), .CLK (CLK)) ;
    ao32 ix2442 (.Y (nx2441), .A0 (Din[22]), .A1 (nx8106), .A2 (FilterWR), .B0 (
         FilterDout_4__2__6), .B1 (nx8198)) ;
    dff L0_4_L1_2_Fij_reg_Dout_7 (.Q (FilterDout_4__2__7), .QB (\$dummy [119]), 
        .D (nx2451), .CLK (CLK)) ;
    ao32 ix2452 (.Y (nx2451), .A0 (Din[23]), .A1 (nx8106), .A2 (FilterWR), .B0 (
         FilterDout_4__2__7), .B1 (nx8200)) ;
    dff L0_4_L1_1_Fij_reg_Dout_0 (.Q (FilterDout_4__1__0), .QB (\$dummy [120]), 
        .D (nx2541), .CLK (CLK)) ;
    ao32 ix2542 (.Y (nx2541), .A0 (Din[8]), .A1 (nx8106), .A2 (FilterWR), .B0 (
         FilterDout_4__1__0), .B1 (nx8200)) ;
    dff L0_4_L1_1_Fij_reg_Dout_1 (.Q (FilterDout_4__1__1), .QB (\$dummy [121]), 
        .D (nx2551), .CLK (CLK)) ;
    ao32 ix2552 (.Y (nx2551), .A0 (Din[9]), .A1 (nx8106), .A2 (FilterWR), .B0 (
         FilterDout_4__1__1), .B1 (nx8200)) ;
    dff L0_4_L1_1_Fij_reg_Dout_2 (.Q (FilterDout_4__1__2), .QB (\$dummy [122]), 
        .D (nx2561), .CLK (CLK)) ;
    ao32 ix2562 (.Y (nx2561), .A0 (Din[10]), .A1 (nx8106), .A2 (FilterWR), .B0 (
         FilterDout_4__1__2), .B1 (nx8200)) ;
    dff L0_4_L1_1_Fij_reg_Dout_3 (.Q (FilterDout_4__1__3), .QB (\$dummy [123]), 
        .D (nx2571), .CLK (CLK)) ;
    ao32 ix2572 (.Y (nx2571), .A0 (Din[11]), .A1 (nx8106), .A2 (FilterWR), .B0 (
         FilterDout_4__1__3), .B1 (nx8200)) ;
    dff L0_4_L1_1_Fij_reg_Dout_4 (.Q (FilterDout_4__1__4), .QB (\$dummy [124]), 
        .D (nx2581), .CLK (CLK)) ;
    ao32 ix2582 (.Y (nx2581), .A0 (Din[12]), .A1 (nx8108), .A2 (FilterWR), .B0 (
         FilterDout_4__1__4), .B1 (nx8200)) ;
    dff L0_4_L1_1_Fij_reg_Dout_5 (.Q (FilterDout_4__1__5), .QB (\$dummy [125]), 
        .D (nx2591), .CLK (CLK)) ;
    ao32 ix2592 (.Y (nx2591), .A0 (Din[13]), .A1 (nx8108), .A2 (FilterWR), .B0 (
         FilterDout_4__1__5), .B1 (nx8200)) ;
    dff L0_4_L1_1_Fij_reg_Dout_6 (.Q (FilterDout_4__1__6), .QB (\$dummy [126]), 
        .D (nx2601), .CLK (CLK)) ;
    ao32 ix2602 (.Y (nx2601), .A0 (Din[14]), .A1 (nx8108), .A2 (FilterWR), .B0 (
         FilterDout_4__1__6), .B1 (nx8202)) ;
    dff L0_4_L1_1_Fij_reg_Dout_7 (.Q (FilterDout_4__1__7), .QB (\$dummy [127]), 
        .D (nx2611), .CLK (CLK)) ;
    ao32 ix2612 (.Y (nx2611), .A0 (Din[15]), .A1 (nx8108), .A2 (FilterWR), .B0 (
         FilterDout_4__1__7), .B1 (nx8202)) ;
    dff L0_4_L1_0_Fij_reg_Dout_0 (.Q (FilterDout_4__0__0), .QB (\$dummy [128]), 
        .D (nx2701), .CLK (CLK)) ;
    ao32 ix2702 (.Y (nx2701), .A0 (Din[0]), .A1 (nx8108), .A2 (FilterWR), .B0 (
         FilterDout_4__0__0), .B1 (nx8202)) ;
    dff L0_4_L1_0_Fij_reg_Dout_1 (.Q (FilterDout_4__0__1), .QB (\$dummy [129]), 
        .D (nx2711), .CLK (CLK)) ;
    ao32 ix2712 (.Y (nx2711), .A0 (Din[1]), .A1 (nx8108), .A2 (FilterWR), .B0 (
         FilterDout_4__0__1), .B1 (nx8202)) ;
    dff L0_4_L1_0_Fij_reg_Dout_2 (.Q (FilterDout_4__0__2), .QB (\$dummy [130]), 
        .D (nx2721), .CLK (CLK)) ;
    ao32 ix2722 (.Y (nx2721), .A0 (Din[2]), .A1 (nx8108), .A2 (FilterWR), .B0 (
         FilterDout_4__0__2), .B1 (nx8202)) ;
    dff L0_4_L1_0_Fij_reg_Dout_3 (.Q (FilterDout_4__0__3), .QB (\$dummy [131]), 
        .D (nx2731), .CLK (CLK)) ;
    ao32 ix2732 (.Y (nx2731), .A0 (Din[3]), .A1 (nx8110), .A2 (FilterWR), .B0 (
         FilterDout_4__0__3), .B1 (nx8202)) ;
    dff L0_4_L1_0_Fij_reg_Dout_4 (.Q (FilterDout_4__0__4), .QB (\$dummy [132]), 
        .D (nx2741), .CLK (CLK)) ;
    ao32 ix2742 (.Y (nx2741), .A0 (Din[4]), .A1 (nx8110), .A2 (FilterWR), .B0 (
         FilterDout_4__0__4), .B1 (nx8202)) ;
    dff L0_4_L1_0_Fij_reg_Dout_5 (.Q (FilterDout_4__0__5), .QB (\$dummy [133]), 
        .D (nx2751), .CLK (CLK)) ;
    ao32 ix2752 (.Y (nx2751), .A0 (Din[5]), .A1 (nx8110), .A2 (FilterWR), .B0 (
         FilterDout_4__0__5), .B1 (nx8204)) ;
    dff L0_4_L1_0_Fij_reg_Dout_6 (.Q (FilterDout_4__0__6), .QB (\$dummy [134]), 
        .D (nx2761), .CLK (CLK)) ;
    ao32 ix2762 (.Y (nx2761), .A0 (Din[6]), .A1 (nx8110), .A2 (FilterWR), .B0 (
         FilterDout_4__0__6), .B1 (nx8204)) ;
    dff L0_4_L1_0_Fij_reg_Dout_7 (.Q (FilterDout_4__0__7), .QB (\$dummy [135]), 
        .D (nx2771), .CLK (CLK)) ;
    ao32 ix2772 (.Y (nx2771), .A0 (Din[7]), .A1 (nx8110), .A2 (FilterWR), .B0 (
         FilterDout_4__0__7), .B1 (nx8204)) ;
    oai21 ix2862 (.Y (nx2861), .A0 (nx7090), .A1 (nx7974), .B0 (nx7093)) ;
    dff L0_3_L1_4_Fij_reg_Dout_0 (.Q (FilterDout_3__4__0), .QB (nx7090), .D (
        nx2861), .CLK (CLK)) ;
    nand03 ix7094 (.Y (nx7093), .A0 (nx8110), .A1 (FilterDout_4__4__0), .A2 (
           nx7974)) ;
    oai21 ix2872 (.Y (nx2871), .A0 (nx7097), .A1 (nx7974), .B0 (nx7099)) ;
    dff L0_3_L1_4_Fij_reg_Dout_1 (.Q (FilterDout_3__4__1), .QB (nx7097), .D (
        nx2871), .CLK (CLK)) ;
    nand03 ix7100 (.Y (nx7099), .A0 (nx8110), .A1 (FilterDout_4__4__1), .A2 (
           nx7974)) ;
    oai21 ix2882 (.Y (nx2881), .A0 (nx7103), .A1 (nx7974), .B0 (nx7105)) ;
    dff L0_3_L1_4_Fij_reg_Dout_2 (.Q (FilterDout_3__4__2), .QB (nx7103), .D (
        nx2881), .CLK (CLK)) ;
    nand03 ix7106 (.Y (nx7105), .A0 (nx8112), .A1 (FilterDout_4__4__2), .A2 (
           nx7974)) ;
    oai21 ix2892 (.Y (nx2891), .A0 (nx7109), .A1 (nx7974), .B0 (nx7111)) ;
    dff L0_3_L1_4_Fij_reg_Dout_3 (.Q (FilterDout_3__4__3), .QB (nx7109), .D (
        nx2891), .CLK (CLK)) ;
    nand03 ix7112 (.Y (nx7111), .A0 (nx8112), .A1 (FilterDout_4__4__3), .A2 (
           nx7976)) ;
    oai21 ix2902 (.Y (nx2901), .A0 (nx7115), .A1 (nx7976), .B0 (nx7117)) ;
    dff L0_3_L1_4_Fij_reg_Dout_4 (.Q (FilterDout_3__4__4), .QB (nx7115), .D (
        nx2901), .CLK (CLK)) ;
    nand03 ix7118 (.Y (nx7117), .A0 (nx8112), .A1 (FilterDout_4__4__4), .A2 (
           nx7976)) ;
    oai21 ix2912 (.Y (nx2911), .A0 (nx7121), .A1 (nx7976), .B0 (nx7123)) ;
    dff L0_3_L1_4_Fij_reg_Dout_5 (.Q (FilterDout_3__4__5), .QB (nx7121), .D (
        nx2911), .CLK (CLK)) ;
    nand03 ix7124 (.Y (nx7123), .A0 (nx8112), .A1 (FilterDout_4__4__5), .A2 (
           nx7976)) ;
    oai21 ix2922 (.Y (nx2921), .A0 (nx7127), .A1 (nx7976), .B0 (nx7129)) ;
    dff L0_3_L1_4_Fij_reg_Dout_6 (.Q (FilterDout_3__4__6), .QB (nx7127), .D (
        nx2921), .CLK (CLK)) ;
    nand03 ix7130 (.Y (nx7129), .A0 (nx8112), .A1 (FilterDout_4__4__6), .A2 (
           nx7976)) ;
    oai21 ix2932 (.Y (nx2931), .A0 (nx7133), .A1 (nx7978), .B0 (nx7135)) ;
    dff L0_3_L1_4_Fij_reg_Dout_7 (.Q (FilterDout_3__4__7), .QB (nx7133), .D (
        nx2931), .CLK (CLK)) ;
    nand03 ix7136 (.Y (nx7135), .A0 (nx8112), .A1 (FilterDout_4__4__7), .A2 (
           nx7978)) ;
    oai21 ix3022 (.Y (nx3021), .A0 (nx7139), .A1 (nx7978), .B0 (nx7141)) ;
    dff L0_3_L1_3_Fij_reg_Dout_0 (.Q (FilterDout_3__3__0), .QB (nx7139), .D (
        nx3021), .CLK (CLK)) ;
    nand03 ix7142 (.Y (nx7141), .A0 (nx8112), .A1 (FilterDout_4__3__0), .A2 (
           nx7978)) ;
    oai21 ix3032 (.Y (nx3031), .A0 (nx7145), .A1 (nx7978), .B0 (nx7147)) ;
    dff L0_3_L1_3_Fij_reg_Dout_1 (.Q (FilterDout_3__3__1), .QB (nx7145), .D (
        nx3031), .CLK (CLK)) ;
    nand03 ix7148 (.Y (nx7147), .A0 (nx8114), .A1 (FilterDout_4__3__1), .A2 (
           nx7978)) ;
    oai21 ix3042 (.Y (nx3041), .A0 (nx7151), .A1 (nx7978), .B0 (nx7153)) ;
    dff L0_3_L1_3_Fij_reg_Dout_2 (.Q (FilterDout_3__3__2), .QB (nx7151), .D (
        nx3041), .CLK (CLK)) ;
    nand03 ix7154 (.Y (nx7153), .A0 (nx8114), .A1 (FilterDout_4__3__2), .A2 (
           nx7980)) ;
    oai21 ix3052 (.Y (nx3051), .A0 (nx7157), .A1 (nx7980), .B0 (nx7159)) ;
    dff L0_3_L1_3_Fij_reg_Dout_3 (.Q (FilterDout_3__3__3), .QB (nx7157), .D (
        nx3051), .CLK (CLK)) ;
    nand03 ix7160 (.Y (nx7159), .A0 (nx8114), .A1 (FilterDout_4__3__3), .A2 (
           nx7980)) ;
    oai21 ix3062 (.Y (nx3061), .A0 (nx7163), .A1 (nx7980), .B0 (nx7165)) ;
    dff L0_3_L1_3_Fij_reg_Dout_4 (.Q (FilterDout_3__3__4), .QB (nx7163), .D (
        nx3061), .CLK (CLK)) ;
    nand03 ix7166 (.Y (nx7165), .A0 (nx8114), .A1 (FilterDout_4__3__4), .A2 (
           nx7980)) ;
    oai21 ix3072 (.Y (nx3071), .A0 (nx7169), .A1 (nx7980), .B0 (nx7171)) ;
    dff L0_3_L1_3_Fij_reg_Dout_5 (.Q (FilterDout_3__3__5), .QB (nx7169), .D (
        nx3071), .CLK (CLK)) ;
    nand03 ix7172 (.Y (nx7171), .A0 (nx8114), .A1 (FilterDout_4__3__5), .A2 (
           nx7980)) ;
    oai21 ix3082 (.Y (nx3081), .A0 (nx7175), .A1 (nx7982), .B0 (nx7177)) ;
    dff L0_3_L1_3_Fij_reg_Dout_6 (.Q (FilterDout_3__3__6), .QB (nx7175), .D (
        nx3081), .CLK (CLK)) ;
    nand03 ix7178 (.Y (nx7177), .A0 (nx8114), .A1 (FilterDout_4__3__6), .A2 (
           nx7982)) ;
    oai21 ix3092 (.Y (nx3091), .A0 (nx7181), .A1 (nx7982), .B0 (nx7183)) ;
    dff L0_3_L1_3_Fij_reg_Dout_7 (.Q (FilterDout_3__3__7), .QB (nx7181), .D (
        nx3091), .CLK (CLK)) ;
    nand03 ix7184 (.Y (nx7183), .A0 (nx8114), .A1 (FilterDout_4__3__7), .A2 (
           nx7982)) ;
    dff L0_3_L1_2_Fij_reg_Dout_0 (.Q (FilterDout_3__2__0), .QB (\$dummy [136]), 
        .D (nx3181), .CLK (CLK)) ;
    ao32 ix3182 (.Y (nx3181), .A0 (nx8116), .A1 (FilterDout_4__2__0), .A2 (
         FilterWR), .B0 (FilterDout_3__2__0), .B1 (nx8204)) ;
    dff L0_3_L1_2_Fij_reg_Dout_1 (.Q (FilterDout_3__2__1), .QB (\$dummy [137]), 
        .D (nx3191), .CLK (CLK)) ;
    ao32 ix3192 (.Y (nx3191), .A0 (nx8116), .A1 (FilterDout_4__2__1), .A2 (
         FilterWR), .B0 (FilterDout_3__2__1), .B1 (nx8204)) ;
    dff L0_3_L1_2_Fij_reg_Dout_2 (.Q (FilterDout_3__2__2), .QB (\$dummy [138]), 
        .D (nx3201), .CLK (CLK)) ;
    ao32 ix3202 (.Y (nx3201), .A0 (nx8116), .A1 (FilterDout_4__2__2), .A2 (
         FilterWR), .B0 (FilterDout_3__2__2), .B1 (nx8204)) ;
    dff L0_3_L1_2_Fij_reg_Dout_3 (.Q (FilterDout_3__2__3), .QB (\$dummy [139]), 
        .D (nx3211), .CLK (CLK)) ;
    ao32 ix3212 (.Y (nx3211), .A0 (nx8116), .A1 (FilterDout_4__2__3), .A2 (
         FilterWR), .B0 (FilterDout_3__2__3), .B1 (nx8204)) ;
    dff L0_3_L1_2_Fij_reg_Dout_4 (.Q (FilterDout_3__2__4), .QB (\$dummy [140]), 
        .D (nx3221), .CLK (CLK)) ;
    ao32 ix3222 (.Y (nx3221), .A0 (nx8116), .A1 (FilterDout_4__2__4), .A2 (
         FilterWR), .B0 (FilterDout_3__2__4), .B1 (nx8206)) ;
    dff L0_3_L1_2_Fij_reg_Dout_5 (.Q (FilterDout_3__2__5), .QB (\$dummy [141]), 
        .D (nx3231), .CLK (CLK)) ;
    ao32 ix3232 (.Y (nx3231), .A0 (nx8116), .A1 (FilterDout_4__2__5), .A2 (
         FilterWR), .B0 (FilterDout_3__2__5), .B1 (nx8206)) ;
    dff L0_3_L1_2_Fij_reg_Dout_6 (.Q (FilterDout_3__2__6), .QB (\$dummy [142]), 
        .D (nx3241), .CLK (CLK)) ;
    ao32 ix3242 (.Y (nx3241), .A0 (nx8116), .A1 (FilterDout_4__2__6), .A2 (
         FilterWR), .B0 (FilterDout_3__2__6), .B1 (nx8206)) ;
    dff L0_3_L1_2_Fij_reg_Dout_7 (.Q (FilterDout_3__2__7), .QB (\$dummy [143]), 
        .D (nx3251), .CLK (CLK)) ;
    ao32 ix3252 (.Y (nx3251), .A0 (nx8118), .A1 (FilterDout_4__2__7), .A2 (
         FilterWR), .B0 (FilterDout_3__2__7), .B1 (nx8206)) ;
    dff L0_3_L1_1_Fij_reg_Dout_0 (.Q (FilterDout_3__1__0), .QB (\$dummy [144]), 
        .D (nx3341), .CLK (CLK)) ;
    ao32 ix3342 (.Y (nx3341), .A0 (nx8118), .A1 (FilterDout_4__1__0), .A2 (
         FilterWR), .B0 (FilterDout_3__1__0), .B1 (nx8206)) ;
    dff L0_3_L1_1_Fij_reg_Dout_1 (.Q (FilterDout_3__1__1), .QB (\$dummy [145]), 
        .D (nx3351), .CLK (CLK)) ;
    ao32 ix3352 (.Y (nx3351), .A0 (nx8118), .A1 (FilterDout_4__1__1), .A2 (
         FilterWR), .B0 (FilterDout_3__1__1), .B1 (nx8206)) ;
    dff L0_3_L1_1_Fij_reg_Dout_2 (.Q (FilterDout_3__1__2), .QB (\$dummy [146]), 
        .D (nx3361), .CLK (CLK)) ;
    ao32 ix3362 (.Y (nx3361), .A0 (nx8118), .A1 (FilterDout_4__1__2), .A2 (
         FilterWR), .B0 (FilterDout_3__1__2), .B1 (nx8206)) ;
    dff L0_3_L1_1_Fij_reg_Dout_3 (.Q (FilterDout_3__1__3), .QB (\$dummy [147]), 
        .D (nx3371), .CLK (CLK)) ;
    ao32 ix3372 (.Y (nx3371), .A0 (nx8118), .A1 (FilterDout_4__1__3), .A2 (
         FilterWR), .B0 (FilterDout_3__1__3), .B1 (nx8208)) ;
    dff L0_3_L1_1_Fij_reg_Dout_4 (.Q (FilterDout_3__1__4), .QB (\$dummy [148]), 
        .D (nx3381), .CLK (CLK)) ;
    ao32 ix3382 (.Y (nx3381), .A0 (nx8118), .A1 (FilterDout_4__1__4), .A2 (
         FilterWR), .B0 (FilterDout_3__1__4), .B1 (nx8208)) ;
    dff L0_3_L1_1_Fij_reg_Dout_5 (.Q (FilterDout_3__1__5), .QB (\$dummy [149]), 
        .D (nx3391), .CLK (CLK)) ;
    ao32 ix3392 (.Y (nx3391), .A0 (nx8118), .A1 (FilterDout_4__1__5), .A2 (
         FilterWR), .B0 (FilterDout_3__1__5), .B1 (nx8208)) ;
    dff L0_3_L1_1_Fij_reg_Dout_6 (.Q (FilterDout_3__1__6), .QB (\$dummy [150]), 
        .D (nx3401), .CLK (CLK)) ;
    ao32 ix3402 (.Y (nx3401), .A0 (nx8120), .A1 (FilterDout_4__1__6), .A2 (
         FilterWR), .B0 (FilterDout_3__1__6), .B1 (nx8208)) ;
    dff L0_3_L1_1_Fij_reg_Dout_7 (.Q (FilterDout_3__1__7), .QB (\$dummy [151]), 
        .D (nx3411), .CLK (CLK)) ;
    ao32 ix3412 (.Y (nx3411), .A0 (nx8120), .A1 (FilterDout_4__1__7), .A2 (
         FilterWR), .B0 (FilterDout_3__1__7), .B1 (nx8208)) ;
    dff L0_3_L1_0_Fij_reg_Dout_0 (.Q (FilterDout_3__0__0), .QB (\$dummy [152]), 
        .D (nx3501), .CLK (CLK)) ;
    ao32 ix3502 (.Y (nx3501), .A0 (nx8120), .A1 (FilterDout_4__0__0), .A2 (
         FilterWR), .B0 (FilterDout_3__0__0), .B1 (nx8208)) ;
    dff L0_3_L1_0_Fij_reg_Dout_1 (.Q (FilterDout_3__0__1), .QB (\$dummy [153]), 
        .D (nx3511), .CLK (CLK)) ;
    ao32 ix3512 (.Y (nx3511), .A0 (nx8120), .A1 (FilterDout_4__0__1), .A2 (
         FilterWR), .B0 (FilterDout_3__0__1), .B1 (nx8208)) ;
    dff L0_3_L1_0_Fij_reg_Dout_2 (.Q (FilterDout_3__0__2), .QB (\$dummy [154]), 
        .D (nx3521), .CLK (CLK)) ;
    ao32 ix3522 (.Y (nx3521), .A0 (nx8120), .A1 (FilterDout_4__0__2), .A2 (
         FilterWR), .B0 (FilterDout_3__0__2), .B1 (nx8210)) ;
    dff L0_3_L1_0_Fij_reg_Dout_3 (.Q (FilterDout_3__0__3), .QB (\$dummy [155]), 
        .D (nx3531), .CLK (CLK)) ;
    ao32 ix3532 (.Y (nx3531), .A0 (nx8120), .A1 (FilterDout_4__0__3), .A2 (
         FilterWR), .B0 (FilterDout_3__0__3), .B1 (nx8210)) ;
    dff L0_3_L1_0_Fij_reg_Dout_4 (.Q (FilterDout_3__0__4), .QB (\$dummy [156]), 
        .D (nx3541), .CLK (CLK)) ;
    ao32 ix3542 (.Y (nx3541), .A0 (nx8120), .A1 (FilterDout_4__0__4), .A2 (
         FilterWR), .B0 (FilterDout_3__0__4), .B1 (nx8210)) ;
    dff L0_3_L1_0_Fij_reg_Dout_5 (.Q (FilterDout_3__0__5), .QB (\$dummy [157]), 
        .D (nx3551), .CLK (CLK)) ;
    ao32 ix3552 (.Y (nx3551), .A0 (nx8122), .A1 (FilterDout_4__0__5), .A2 (
         FilterWR), .B0 (FilterDout_3__0__5), .B1 (nx8210)) ;
    dff L0_3_L1_0_Fij_reg_Dout_6 (.Q (FilterDout_3__0__6), .QB (\$dummy [158]), 
        .D (nx3561), .CLK (CLK)) ;
    ao32 ix3562 (.Y (nx3561), .A0 (nx8122), .A1 (FilterDout_4__0__6), .A2 (
         FilterWR), .B0 (FilterDout_3__0__6), .B1 (nx8210)) ;
    dff L0_3_L1_0_Fij_reg_Dout_7 (.Q (FilterDout_3__0__7), .QB (\$dummy [159]), 
        .D (nx3571), .CLK (CLK)) ;
    ao32 ix3572 (.Y (nx3571), .A0 (nx8122), .A1 (FilterDout_4__0__7), .A2 (
         FilterWR), .B0 (FilterDout_3__0__7), .B1 (nx8210)) ;
    oai21 ix3662 (.Y (nx3661), .A0 (nx7259), .A1 (nx7982), .B0 (nx7261)) ;
    dff L0_2_L1_4_Fij_reg_Dout_0 (.Q (FilterDout_2__4__0), .QB (nx7259), .D (
        nx3661), .CLK (CLK)) ;
    oai21 ix3672 (.Y (nx3671), .A0 (nx7265), .A1 (nx7982), .B0 (nx7267)) ;
    dff L0_2_L1_4_Fij_reg_Dout_1 (.Q (FilterDout_2__4__1), .QB (nx7265), .D (
        nx3671), .CLK (CLK)) ;
    oai21 ix3682 (.Y (nx3681), .A0 (nx7271), .A1 (nx7984), .B0 (nx7273)) ;
    dff L0_2_L1_4_Fij_reg_Dout_2 (.Q (FilterDout_2__4__2), .QB (nx7271), .D (
        nx3681), .CLK (CLK)) ;
    oai21 ix3692 (.Y (nx3691), .A0 (nx7277), .A1 (nx7984), .B0 (nx7279)) ;
    dff L0_2_L1_4_Fij_reg_Dout_3 (.Q (FilterDout_2__4__3), .QB (nx7277), .D (
        nx3691), .CLK (CLK)) ;
    oai21 ix3702 (.Y (nx3701), .A0 (nx7283), .A1 (nx7984), .B0 (nx7285)) ;
    dff L0_2_L1_4_Fij_reg_Dout_4 (.Q (FilterDout_2__4__4), .QB (nx7283), .D (
        nx3701), .CLK (CLK)) ;
    oai21 ix3712 (.Y (nx3711), .A0 (nx7289), .A1 (nx7986), .B0 (nx7291)) ;
    dff L0_2_L1_4_Fij_reg_Dout_5 (.Q (FilterDout_2__4__5), .QB (nx7289), .D (
        nx3711), .CLK (CLK)) ;
    oai21 ix3722 (.Y (nx3721), .A0 (nx7295), .A1 (nx7986), .B0 (nx7297)) ;
    dff L0_2_L1_4_Fij_reg_Dout_6 (.Q (FilterDout_2__4__6), .QB (nx7295), .D (
        nx3721), .CLK (CLK)) ;
    oai21 ix3732 (.Y (nx3731), .A0 (nx7301), .A1 (nx7986), .B0 (nx7303)) ;
    dff L0_2_L1_4_Fij_reg_Dout_7 (.Q (FilterDout_2__4__7), .QB (nx7301), .D (
        nx3731), .CLK (CLK)) ;
    oai21 ix3822 (.Y (nx3821), .A0 (nx7307), .A1 (nx7986), .B0 (nx7309)) ;
    dff L0_2_L1_3_Fij_reg_Dout_0 (.Q (FilterDout_2__3__0), .QB (nx7307), .D (
        nx3821), .CLK (CLK)) ;
    oai21 ix3832 (.Y (nx3831), .A0 (nx7313), .A1 (nx7988), .B0 (nx7315)) ;
    dff L0_2_L1_3_Fij_reg_Dout_1 (.Q (FilterDout_2__3__1), .QB (nx7313), .D (
        nx3831), .CLK (CLK)) ;
    oai21 ix3842 (.Y (nx3841), .A0 (nx7319), .A1 (nx7988), .B0 (nx7321)) ;
    dff L0_2_L1_3_Fij_reg_Dout_2 (.Q (FilterDout_2__3__2), .QB (nx7319), .D (
        nx3841), .CLK (CLK)) ;
    oai21 ix3852 (.Y (nx3851), .A0 (nx7325), .A1 (nx7988), .B0 (nx7327)) ;
    dff L0_2_L1_3_Fij_reg_Dout_3 (.Q (FilterDout_2__3__3), .QB (nx7325), .D (
        nx3851), .CLK (CLK)) ;
    oai21 ix3862 (.Y (nx3861), .A0 (nx7331), .A1 (nx7990), .B0 (nx7333)) ;
    dff L0_2_L1_3_Fij_reg_Dout_4 (.Q (FilterDout_2__3__4), .QB (nx7331), .D (
        nx3861), .CLK (CLK)) ;
    oai21 ix3872 (.Y (nx3871), .A0 (nx7337), .A1 (nx7990), .B0 (nx7339)) ;
    dff L0_2_L1_3_Fij_reg_Dout_5 (.Q (FilterDout_2__3__5), .QB (nx7337), .D (
        nx3871), .CLK (CLK)) ;
    oai21 ix3882 (.Y (nx3881), .A0 (nx7343), .A1 (nx7990), .B0 (nx7345)) ;
    dff L0_2_L1_3_Fij_reg_Dout_6 (.Q (FilterDout_2__3__6), .QB (nx7343), .D (
        nx3881), .CLK (CLK)) ;
    oai21 ix3892 (.Y (nx3891), .A0 (nx7349), .A1 (nx7990), .B0 (nx7351)) ;
    dff L0_2_L1_3_Fij_reg_Dout_7 (.Q (FilterDout_2__3__7), .QB (nx7349), .D (
        nx3891), .CLK (CLK)) ;
    dff L0_2_L1_2_Fij_reg_Dout_0 (.Q (FilterDout_2__2__0), .QB (\$dummy [160]), 
        .D (nx3981), .CLK (CLK)) ;
    ao32 ix3982 (.Y (nx3981), .A0 (nx8126), .A1 (FilterDout_3__2__0), .A2 (
         FilterWR), .B0 (FilterDout_2__2__0), .B1 (nx8210)) ;
    dff L0_2_L1_2_Fij_reg_Dout_1 (.Q (FilterDout_2__2__1), .QB (\$dummy [161]), 
        .D (nx3991), .CLK (CLK)) ;
    ao32 ix3992 (.Y (nx3991), .A0 (nx8126), .A1 (FilterDout_3__2__1), .A2 (
         FilterWR), .B0 (FilterDout_2__2__1), .B1 (nx8212)) ;
    dff L0_2_L1_2_Fij_reg_Dout_2 (.Q (FilterDout_2__2__2), .QB (\$dummy [162]), 
        .D (nx4001), .CLK (CLK)) ;
    ao32 ix4002 (.Y (nx4001), .A0 (nx8128), .A1 (FilterDout_3__2__2), .A2 (
         FilterWR), .B0 (FilterDout_2__2__2), .B1 (nx8212)) ;
    dff L0_2_L1_2_Fij_reg_Dout_3 (.Q (FilterDout_2__2__3), .QB (\$dummy [163]), 
        .D (nx4011), .CLK (CLK)) ;
    ao32 ix4012 (.Y (nx4011), .A0 (nx8128), .A1 (FilterDout_3__2__3), .A2 (
         FilterWR), .B0 (FilterDout_2__2__3), .B1 (nx8212)) ;
    dff L0_2_L1_2_Fij_reg_Dout_4 (.Q (FilterDout_2__2__4), .QB (\$dummy [164]), 
        .D (nx4021), .CLK (CLK)) ;
    ao32 ix4022 (.Y (nx4021), .A0 (nx8128), .A1 (FilterDout_3__2__4), .A2 (
         FilterWR), .B0 (FilterDout_2__2__4), .B1 (nx8212)) ;
    dff L0_2_L1_2_Fij_reg_Dout_5 (.Q (FilterDout_2__2__5), .QB (\$dummy [165]), 
        .D (nx4031), .CLK (CLK)) ;
    ao32 ix4032 (.Y (nx4031), .A0 (nx8128), .A1 (FilterDout_3__2__5), .A2 (
         FilterWR), .B0 (FilterDout_2__2__5), .B1 (nx8212)) ;
    dff L0_2_L1_2_Fij_reg_Dout_6 (.Q (FilterDout_2__2__6), .QB (\$dummy [166]), 
        .D (nx4041), .CLK (CLK)) ;
    ao32 ix4042 (.Y (nx4041), .A0 (nx8128), .A1 (FilterDout_3__2__6), .A2 (
         FilterWR), .B0 (FilterDout_2__2__6), .B1 (nx8212)) ;
    dff L0_2_L1_2_Fij_reg_Dout_7 (.Q (FilterDout_2__2__7), .QB (\$dummy [167]), 
        .D (nx4051), .CLK (CLK)) ;
    ao32 ix4052 (.Y (nx4051), .A0 (nx8128), .A1 (FilterDout_3__2__7), .A2 (
         FilterWR), .B0 (FilterDout_2__2__7), .B1 (nx8212)) ;
    dff L0_2_L1_1_Fij_reg_Dout_0 (.Q (FilterDout_2__1__0), .QB (\$dummy [168]), 
        .D (nx4141), .CLK (CLK)) ;
    ao32 ix4142 (.Y (nx4141), .A0 (nx8128), .A1 (FilterDout_3__1__0), .A2 (
         FilterWR), .B0 (FilterDout_2__1__0), .B1 (nx8214)) ;
    dff L0_2_L1_1_Fij_reg_Dout_1 (.Q (FilterDout_2__1__1), .QB (\$dummy [169]), 
        .D (nx4151), .CLK (CLK)) ;
    ao32 ix4152 (.Y (nx4151), .A0 (nx8130), .A1 (FilterDout_3__1__1), .A2 (
         FilterWR), .B0 (FilterDout_2__1__1), .B1 (nx8214)) ;
    dff L0_2_L1_1_Fij_reg_Dout_2 (.Q (FilterDout_2__1__2), .QB (\$dummy [170]), 
        .D (nx4161), .CLK (CLK)) ;
    ao32 ix4162 (.Y (nx4161), .A0 (nx8130), .A1 (FilterDout_3__1__2), .A2 (
         FilterWR), .B0 (FilterDout_2__1__2), .B1 (nx8214)) ;
    dff L0_2_L1_1_Fij_reg_Dout_3 (.Q (FilterDout_2__1__3), .QB (\$dummy [171]), 
        .D (nx4171), .CLK (CLK)) ;
    ao32 ix4172 (.Y (nx4171), .A0 (nx8130), .A1 (FilterDout_3__1__3), .A2 (
         FilterWR), .B0 (FilterDout_2__1__3), .B1 (nx8214)) ;
    dff L0_2_L1_1_Fij_reg_Dout_4 (.Q (FilterDout_2__1__4), .QB (\$dummy [172]), 
        .D (nx4181), .CLK (CLK)) ;
    ao32 ix4182 (.Y (nx4181), .A0 (nx8130), .A1 (FilterDout_3__1__4), .A2 (
         FilterWR), .B0 (FilterDout_2__1__4), .B1 (nx8214)) ;
    dff L0_2_L1_1_Fij_reg_Dout_5 (.Q (FilterDout_2__1__5), .QB (\$dummy [173]), 
        .D (nx4191), .CLK (CLK)) ;
    ao32 ix4192 (.Y (nx4191), .A0 (nx8130), .A1 (FilterDout_3__1__5), .A2 (
         FilterWR), .B0 (FilterDout_2__1__5), .B1 (nx8214)) ;
    dff L0_2_L1_1_Fij_reg_Dout_6 (.Q (FilterDout_2__1__6), .QB (\$dummy [174]), 
        .D (nx4201), .CLK (CLK)) ;
    ao32 ix4202 (.Y (nx4201), .A0 (nx8130), .A1 (FilterDout_3__1__6), .A2 (
         FilterWR), .B0 (FilterDout_2__1__6), .B1 (nx8214)) ;
    dff L0_2_L1_1_Fij_reg_Dout_7 (.Q (FilterDout_2__1__7), .QB (\$dummy [175]), 
        .D (nx4211), .CLK (CLK)) ;
    ao32 ix4212 (.Y (nx4211), .A0 (nx8130), .A1 (FilterDout_3__1__7), .A2 (
         FilterWR), .B0 (FilterDout_2__1__7), .B1 (nx8216)) ;
    dff L0_2_L1_0_Fij_reg_Dout_0 (.Q (FilterDout_2__0__0), .QB (\$dummy [176]), 
        .D (nx4301), .CLK (CLK)) ;
    ao32 ix4302 (.Y (nx4301), .A0 (nx8132), .A1 (FilterDout_3__0__0), .A2 (
         FilterWR), .B0 (FilterDout_2__0__0), .B1 (nx8216)) ;
    dff L0_2_L1_0_Fij_reg_Dout_1 (.Q (FilterDout_2__0__1), .QB (\$dummy [177]), 
        .D (nx4311), .CLK (CLK)) ;
    ao32 ix4312 (.Y (nx4311), .A0 (nx8132), .A1 (FilterDout_3__0__1), .A2 (
         FilterWR), .B0 (FilterDout_2__0__1), .B1 (nx8216)) ;
    dff L0_2_L1_0_Fij_reg_Dout_2 (.Q (FilterDout_2__0__2), .QB (\$dummy [178]), 
        .D (nx4321), .CLK (CLK)) ;
    ao32 ix4322 (.Y (nx4321), .A0 (nx8132), .A1 (FilterDout_3__0__2), .A2 (
         FilterWR), .B0 (FilterDout_2__0__2), .B1 (nx8216)) ;
    dff L0_2_L1_0_Fij_reg_Dout_3 (.Q (FilterDout_2__0__3), .QB (\$dummy [179]), 
        .D (nx4331), .CLK (CLK)) ;
    ao32 ix4332 (.Y (nx4331), .A0 (nx8132), .A1 (FilterDout_3__0__3), .A2 (
         FilterWR), .B0 (FilterDout_2__0__3), .B1 (nx8216)) ;
    dff L0_2_L1_0_Fij_reg_Dout_4 (.Q (FilterDout_2__0__4), .QB (\$dummy [180]), 
        .D (nx4341), .CLK (CLK)) ;
    ao32 ix4342 (.Y (nx4341), .A0 (nx8132), .A1 (FilterDout_3__0__4), .A2 (
         FilterWR), .B0 (FilterDout_2__0__4), .B1 (nx8216)) ;
    dff L0_2_L1_0_Fij_reg_Dout_5 (.Q (FilterDout_2__0__5), .QB (\$dummy [181]), 
        .D (nx4351), .CLK (CLK)) ;
    ao32 ix4352 (.Y (nx4351), .A0 (nx8132), .A1 (FilterDout_3__0__5), .A2 (
         FilterWR), .B0 (FilterDout_2__0__5), .B1 (nx8216)) ;
    dff L0_2_L1_0_Fij_reg_Dout_6 (.Q (FilterDout_2__0__6), .QB (\$dummy [182]), 
        .D (nx4361), .CLK (CLK)) ;
    ao32 ix4362 (.Y (nx4361), .A0 (nx8132), .A1 (FilterDout_3__0__6), .A2 (
         FilterWR), .B0 (FilterDout_2__0__6), .B1 (nx8218)) ;
    dff L0_2_L1_0_Fij_reg_Dout_7 (.Q (FilterDout_2__0__7), .QB (\$dummy [183]), 
        .D (nx4371), .CLK (CLK)) ;
    ao32 ix4372 (.Y (nx4371), .A0 (nx8134), .A1 (FilterDout_3__0__7), .A2 (
         FilterWR), .B0 (FilterDout_2__0__7), .B1 (nx8218)) ;
    oai21 ix4542 (.Y (nx4541), .A0 (nx7427), .A1 (nx7992), .B0 (nx7429)) ;
    dff L0_1_L1_4_Fij_reg_Dout_0 (.Q (FilterDout_1__4__0), .QB (nx7427), .D (
        nx4541), .CLK (CLK)) ;
    oai21 ix4552 (.Y (nx4551), .A0 (nx7433), .A1 (nx7992), .B0 (nx7435)) ;
    dff L0_1_L1_4_Fij_reg_Dout_1 (.Q (FilterDout_1__4__1), .QB (nx7433), .D (
        nx4551), .CLK (CLK)) ;
    oai21 ix4562 (.Y (nx4561), .A0 (nx7439), .A1 (nx7992), .B0 (nx7441)) ;
    dff L0_1_L1_4_Fij_reg_Dout_2 (.Q (FilterDout_1__4__2), .QB (nx7439), .D (
        nx4561), .CLK (CLK)) ;
    oai21 ix4572 (.Y (nx4571), .A0 (nx7445), .A1 (nx7994), .B0 (nx7447)) ;
    dff L0_1_L1_4_Fij_reg_Dout_3 (.Q (FilterDout_1__4__3), .QB (nx7445), .D (
        nx4571), .CLK (CLK)) ;
    oai21 ix4582 (.Y (nx4581), .A0 (nx7451), .A1 (nx7994), .B0 (nx7453)) ;
    dff L0_1_L1_4_Fij_reg_Dout_4 (.Q (FilterDout_1__4__4), .QB (nx7451), .D (
        nx4581), .CLK (CLK)) ;
    oai21 ix4592 (.Y (nx4591), .A0 (nx7457), .A1 (nx7994), .B0 (nx7459)) ;
    dff L0_1_L1_4_Fij_reg_Dout_5 (.Q (FilterDout_1__4__5), .QB (nx7457), .D (
        nx4591), .CLK (CLK)) ;
    oai21 ix4602 (.Y (nx4601), .A0 (nx7463), .A1 (nx7994), .B0 (nx7465)) ;
    dff L0_1_L1_4_Fij_reg_Dout_6 (.Q (FilterDout_1__4__6), .QB (nx7463), .D (
        nx4601), .CLK (CLK)) ;
    oai21 ix4612 (.Y (nx4611), .A0 (nx7469), .A1 (nx7996), .B0 (nx7471)) ;
    dff L0_1_L1_4_Fij_reg_Dout_7 (.Q (FilterDout_1__4__7), .QB (nx7469), .D (
        nx4611), .CLK (CLK)) ;
    oai21 ix4862 (.Y (nx4861), .A0 (nx7475), .A1 (nx7996), .B0 (nx7477)) ;
    dff L0_1_L1_3_Fij_reg_Dout_0 (.Q (FilterDout_1__3__0), .QB (nx7475), .D (
        nx4861), .CLK (CLK)) ;
    oai21 ix4872 (.Y (nx4871), .A0 (nx7481), .A1 (nx7996), .B0 (nx7483)) ;
    dff L0_1_L1_3_Fij_reg_Dout_1 (.Q (FilterDout_1__3__1), .QB (nx7481), .D (
        nx4871), .CLK (CLK)) ;
    oai21 ix4882 (.Y (nx4881), .A0 (nx7487), .A1 (nx7998), .B0 (nx7489)) ;
    dff L0_1_L1_3_Fij_reg_Dout_2 (.Q (FilterDout_1__3__2), .QB (nx7487), .D (
        nx4881), .CLK (CLK)) ;
    oai21 ix4892 (.Y (nx4891), .A0 (nx7493), .A1 (nx7998), .B0 (nx7495)) ;
    dff L0_1_L1_3_Fij_reg_Dout_3 (.Q (FilterDout_1__3__3), .QB (nx7493), .D (
        nx4891), .CLK (CLK)) ;
    oai21 ix4902 (.Y (nx4901), .A0 (nx7499), .A1 (nx7998), .B0 (nx7501)) ;
    dff L0_1_L1_3_Fij_reg_Dout_4 (.Q (FilterDout_1__3__4), .QB (nx7499), .D (
        nx4901), .CLK (CLK)) ;
    oai21 ix4912 (.Y (nx4911), .A0 (nx7505), .A1 (nx7998), .B0 (nx7507)) ;
    dff L0_1_L1_3_Fij_reg_Dout_5 (.Q (FilterDout_1__3__5), .QB (nx7505), .D (
        nx4911), .CLK (CLK)) ;
    oai21 ix4922 (.Y (nx4921), .A0 (nx7511), .A1 (nx8000), .B0 (nx7513)) ;
    dff L0_1_L1_3_Fij_reg_Dout_6 (.Q (FilterDout_1__3__6), .QB (nx7511), .D (
        nx4921), .CLK (CLK)) ;
    oai21 ix4932 (.Y (nx4931), .A0 (nx7517), .A1 (nx8000), .B0 (nx7519)) ;
    dff L0_1_L1_3_Fij_reg_Dout_7 (.Q (FilterDout_1__3__7), .QB (nx7517), .D (
        nx4931), .CLK (CLK)) ;
    oai21 ix5182 (.Y (nx5181), .A0 (nx7523), .A1 (nx8000), .B0 (nx7525)) ;
    dff L0_1_L1_2_Fij_reg_Dout_0 (.Q (FilterDout_1__2__0), .QB (nx7523), .D (
        nx5181), .CLK (CLK)) ;
    nand03 ix7526 (.Y (nx7525), .A0 (nx8138), .A1 (FilterDout_2__2__0), .A2 (
           nx8000)) ;
    oai21 ix5192 (.Y (nx5191), .A0 (nx7529), .A1 (nx8002), .B0 (nx7531)) ;
    dff L0_1_L1_2_Fij_reg_Dout_1 (.Q (FilterDout_1__2__1), .QB (nx7529), .D (
        nx5191), .CLK (CLK)) ;
    nand03 ix7532 (.Y (nx7531), .A0 (nx8138), .A1 (FilterDout_2__2__1), .A2 (
           nx8002)) ;
    oai21 ix5202 (.Y (nx5201), .A0 (nx7535), .A1 (nx8002), .B0 (nx7537)) ;
    dff L0_1_L1_2_Fij_reg_Dout_2 (.Q (FilterDout_1__2__2), .QB (nx7535), .D (
        nx5201), .CLK (CLK)) ;
    nand03 ix7538 (.Y (nx7537), .A0 (nx8138), .A1 (FilterDout_2__2__2), .A2 (
           nx8002)) ;
    oai21 ix5212 (.Y (nx5211), .A0 (nx7541), .A1 (nx8002), .B0 (nx7543)) ;
    dff L0_1_L1_2_Fij_reg_Dout_3 (.Q (FilterDout_1__2__3), .QB (nx7541), .D (
        nx5211), .CLK (CLK)) ;
    nand03 ix7544 (.Y (nx7543), .A0 (nx8138), .A1 (FilterDout_2__2__3), .A2 (
           nx8002)) ;
    oai21 ix5222 (.Y (nx5221), .A0 (nx7547), .A1 (nx8002), .B0 (nx7549)) ;
    dff L0_1_L1_2_Fij_reg_Dout_4 (.Q (FilterDout_1__2__4), .QB (nx7547), .D (
        nx5221), .CLK (CLK)) ;
    nand03 ix7550 (.Y (nx7549), .A0 (nx8140), .A1 (FilterDout_2__2__4), .A2 (
           nx8004)) ;
    oai21 ix5232 (.Y (nx5231), .A0 (nx7553), .A1 (nx8004), .B0 (nx7555)) ;
    dff L0_1_L1_2_Fij_reg_Dout_5 (.Q (FilterDout_1__2__5), .QB (nx7553), .D (
        nx5231), .CLK (CLK)) ;
    nand03 ix7556 (.Y (nx7555), .A0 (nx8140), .A1 (FilterDout_2__2__5), .A2 (
           nx8004)) ;
    oai21 ix5242 (.Y (nx5241), .A0 (nx7559), .A1 (nx8004), .B0 (nx7561)) ;
    dff L0_1_L1_2_Fij_reg_Dout_6 (.Q (FilterDout_1__2__6), .QB (nx7559), .D (
        nx5241), .CLK (CLK)) ;
    nand03 ix7562 (.Y (nx7561), .A0 (nx8140), .A1 (FilterDout_2__2__6), .A2 (
           nx8004)) ;
    oai21 ix5252 (.Y (nx5251), .A0 (nx7565), .A1 (nx8004), .B0 (nx7567)) ;
    dff L0_1_L1_2_Fij_reg_Dout_7 (.Q (FilterDout_1__2__7), .QB (nx7565), .D (
        nx5251), .CLK (CLK)) ;
    nand03 ix7568 (.Y (nx7567), .A0 (nx8140), .A1 (FilterDout_2__2__7), .A2 (
           nx8004)) ;
    oai21 ix5502 (.Y (nx5501), .A0 (nx7571), .A1 (nx8006), .B0 (nx7573)) ;
    dff L0_1_L1_1_Fij_reg_Dout_0 (.Q (FilterDout_1__1__0), .QB (nx7571), .D (
        nx5501), .CLK (CLK)) ;
    nand03 ix7574 (.Y (nx7573), .A0 (nx8140), .A1 (FilterDout_2__1__0), .A2 (
           nx8006)) ;
    oai21 ix5512 (.Y (nx5511), .A0 (nx7577), .A1 (nx8006), .B0 (nx7579)) ;
    dff L0_1_L1_1_Fij_reg_Dout_1 (.Q (FilterDout_1__1__1), .QB (nx7577), .D (
        nx5511), .CLK (CLK)) ;
    nand03 ix7580 (.Y (nx7579), .A0 (nx8140), .A1 (FilterDout_2__1__1), .A2 (
           nx8006)) ;
    oai21 ix5522 (.Y (nx5521), .A0 (nx7583), .A1 (nx8006), .B0 (nx7585)) ;
    dff L0_1_L1_1_Fij_reg_Dout_2 (.Q (FilterDout_1__1__2), .QB (nx7583), .D (
        nx5521), .CLK (CLK)) ;
    nand03 ix7586 (.Y (nx7585), .A0 (nx8140), .A1 (FilterDout_2__1__2), .A2 (
           nx8006)) ;
    oai21 ix5532 (.Y (nx5531), .A0 (nx7589), .A1 (nx8006), .B0 (nx7591)) ;
    dff L0_1_L1_1_Fij_reg_Dout_3 (.Q (FilterDout_1__1__3), .QB (nx7589), .D (
        nx5531), .CLK (CLK)) ;
    nand03 ix7592 (.Y (nx7591), .A0 (nx8142), .A1 (FilterDout_2__1__3), .A2 (
           nx8008)) ;
    oai21 ix5542 (.Y (nx5541), .A0 (nx7595), .A1 (nx8008), .B0 (nx7597)) ;
    dff L0_1_L1_1_Fij_reg_Dout_4 (.Q (FilterDout_1__1__4), .QB (nx7595), .D (
        nx5541), .CLK (CLK)) ;
    nand03 ix7598 (.Y (nx7597), .A0 (nx8142), .A1 (FilterDout_2__1__4), .A2 (
           nx8008)) ;
    oai21 ix5552 (.Y (nx5551), .A0 (nx7601), .A1 (nx8008), .B0 (nx7603)) ;
    dff L0_1_L1_1_Fij_reg_Dout_5 (.Q (FilterDout_1__1__5), .QB (nx7601), .D (
        nx5551), .CLK (CLK)) ;
    nand03 ix7604 (.Y (nx7603), .A0 (nx8142), .A1 (FilterDout_2__1__5), .A2 (
           nx8008)) ;
    oai21 ix5562 (.Y (nx5561), .A0 (nx7607), .A1 (nx8008), .B0 (nx7609)) ;
    dff L0_1_L1_1_Fij_reg_Dout_6 (.Q (FilterDout_1__1__6), .QB (nx7607), .D (
        nx5561), .CLK (CLK)) ;
    nand03 ix7610 (.Y (nx7609), .A0 (nx8142), .A1 (FilterDout_2__1__6), .A2 (
           nx8008)) ;
    oai21 ix5572 (.Y (nx5571), .A0 (nx7613), .A1 (nx8010), .B0 (nx7615)) ;
    dff L0_1_L1_1_Fij_reg_Dout_7 (.Q (FilterDout_1__1__7), .QB (nx7613), .D (
        nx5571), .CLK (CLK)) ;
    nand03 ix7616 (.Y (nx7615), .A0 (nx8142), .A1 (FilterDout_2__1__7), .A2 (
           nx8010)) ;
    oai21 ix5822 (.Y (nx5821), .A0 (nx7619), .A1 (nx8010), .B0 (nx7621)) ;
    dff L0_1_L1_0_Fij_reg_Dout_0 (.Q (FilterDout_1__0__0), .QB (nx7619), .D (
        nx5821), .CLK (CLK)) ;
    nand03 ix7622 (.Y (nx7621), .A0 (nx8142), .A1 (FilterDout_2__0__0), .A2 (
           nx8010)) ;
    oai21 ix5832 (.Y (nx5831), .A0 (nx7625), .A1 (nx8010), .B0 (nx7627)) ;
    dff L0_1_L1_0_Fij_reg_Dout_1 (.Q (FilterDout_1__0__1), .QB (nx7625), .D (
        nx5831), .CLK (CLK)) ;
    nand03 ix7628 (.Y (nx7627), .A0 (nx8142), .A1 (FilterDout_2__0__1), .A2 (
           nx8010)) ;
    oai21 ix5842 (.Y (nx5841), .A0 (nx7631), .A1 (nx8010), .B0 (nx7633)) ;
    dff L0_1_L1_0_Fij_reg_Dout_2 (.Q (FilterDout_1__0__2), .QB (nx7631), .D (
        nx5841), .CLK (CLK)) ;
    nand03 ix7634 (.Y (nx7633), .A0 (nx8144), .A1 (FilterDout_2__0__2), .A2 (
           nx8012)) ;
    oai21 ix5852 (.Y (nx5851), .A0 (nx7637), .A1 (nx8012), .B0 (nx7639)) ;
    dff L0_1_L1_0_Fij_reg_Dout_3 (.Q (FilterDout_1__0__3), .QB (nx7637), .D (
        nx5851), .CLK (CLK)) ;
    nand03 ix7640 (.Y (nx7639), .A0 (nx8144), .A1 (FilterDout_2__0__3), .A2 (
           nx8012)) ;
    oai21 ix5862 (.Y (nx5861), .A0 (nx7643), .A1 (nx8012), .B0 (nx7645)) ;
    dff L0_1_L1_0_Fij_reg_Dout_4 (.Q (FilterDout_1__0__4), .QB (nx7643), .D (
        nx5861), .CLK (CLK)) ;
    nand03 ix7646 (.Y (nx7645), .A0 (nx8144), .A1 (FilterDout_2__0__4), .A2 (
           nx8012)) ;
    oai21 ix5872 (.Y (nx5871), .A0 (nx7649), .A1 (nx8012), .B0 (nx7651)) ;
    dff L0_1_L1_0_Fij_reg_Dout_5 (.Q (FilterDout_1__0__5), .QB (nx7649), .D (
        nx5871), .CLK (CLK)) ;
    nand03 ix7652 (.Y (nx7651), .A0 (nx8144), .A1 (FilterDout_2__0__5), .A2 (
           nx8012)) ;
    oai21 ix5882 (.Y (nx5881), .A0 (nx7655), .A1 (nx8014), .B0 (nx7657)) ;
    dff L0_1_L1_0_Fij_reg_Dout_6 (.Q (FilterDout_1__0__6), .QB (nx7655), .D (
        nx5881), .CLK (CLK)) ;
    nand03 ix7658 (.Y (nx7657), .A0 (nx8144), .A1 (FilterDout_2__0__6), .A2 (
           nx8014)) ;
    oai21 ix5892 (.Y (nx5891), .A0 (nx7661), .A1 (nx8014), .B0 (nx7663)) ;
    dff L0_1_L1_0_Fij_reg_Dout_7 (.Q (FilterDout_1__0__7), .QB (nx7661), .D (
        nx5891), .CLK (CLK)) ;
    nand03 ix7664 (.Y (nx7663), .A0 (nx8144), .A1 (FilterDout_2__0__7), .A2 (
           nx8014)) ;
    oai21 ix4622 (.Y (nx4621), .A0 (nx7667), .A1 (nx8014), .B0 (nx7669)) ;
    dff L0_0_L1_4_Fij_reg_Dout_0 (.Q (FilterDout_0__4__0), .QB (nx7667), .D (
        nx4621), .CLK (CLK)) ;
    oai21 ix4632 (.Y (nx4631), .A0 (nx7673), .A1 (nx8014), .B0 (nx7675)) ;
    dff L0_0_L1_4_Fij_reg_Dout_1 (.Q (FilterDout_0__4__1), .QB (nx7673), .D (
        nx4631), .CLK (CLK)) ;
    oai21 ix4642 (.Y (nx4641), .A0 (nx7679), .A1 (nx8016), .B0 (nx7681)) ;
    dff L0_0_L1_4_Fij_reg_Dout_2 (.Q (FilterDout_0__4__2), .QB (nx7679), .D (
        nx4641), .CLK (CLK)) ;
    oai21 ix4652 (.Y (nx4651), .A0 (nx7685), .A1 (nx8016), .B0 (nx7687)) ;
    dff L0_0_L1_4_Fij_reg_Dout_3 (.Q (FilterDout_0__4__3), .QB (nx7685), .D (
        nx4651), .CLK (CLK)) ;
    oai21 ix4662 (.Y (nx4661), .A0 (nx7691), .A1 (nx8016), .B0 (nx7693)) ;
    dff L0_0_L1_4_Fij_reg_Dout_4 (.Q (FilterDout_0__4__4), .QB (nx7691), .D (
        nx4661), .CLK (CLK)) ;
    oai21 ix4672 (.Y (nx4671), .A0 (nx7697), .A1 (nx8018), .B0 (nx7699)) ;
    dff L0_0_L1_4_Fij_reg_Dout_5 (.Q (FilterDout_0__4__5), .QB (nx7697), .D (
        nx4671), .CLK (CLK)) ;
    oai21 ix4682 (.Y (nx4681), .A0 (nx7703), .A1 (nx8018), .B0 (nx7705)) ;
    dff L0_0_L1_4_Fij_reg_Dout_6 (.Q (FilterDout_0__4__6), .QB (nx7703), .D (
        nx4681), .CLK (CLK)) ;
    oai21 ix4692 (.Y (nx4691), .A0 (nx7709), .A1 (nx8018), .B0 (nx7711)) ;
    dff L0_0_L1_4_Fij_reg_Dout_7 (.Q (FilterDout_0__4__7), .QB (nx7709), .D (
        nx4691), .CLK (CLK)) ;
    oai21 ix4942 (.Y (nx4941), .A0 (nx7715), .A1 (nx8018), .B0 (nx7717)) ;
    dff L0_0_L1_3_Fij_reg_Dout_0 (.Q (FilterDout_0__3__0), .QB (nx7715), .D (
        nx4941), .CLK (CLK)) ;
    oai21 ix4952 (.Y (nx4951), .A0 (nx7721), .A1 (nx8020), .B0 (nx7723)) ;
    dff L0_0_L1_3_Fij_reg_Dout_1 (.Q (FilterDout_0__3__1), .QB (nx7721), .D (
        nx4951), .CLK (CLK)) ;
    oai21 ix4962 (.Y (nx4961), .A0 (nx7727), .A1 (nx8020), .B0 (nx7729)) ;
    dff L0_0_L1_3_Fij_reg_Dout_2 (.Q (FilterDout_0__3__2), .QB (nx7727), .D (
        nx4961), .CLK (CLK)) ;
    oai21 ix4972 (.Y (nx4971), .A0 (nx7733), .A1 (nx8020), .B0 (nx7735)) ;
    dff L0_0_L1_3_Fij_reg_Dout_3 (.Q (FilterDout_0__3__3), .QB (nx7733), .D (
        nx4971), .CLK (CLK)) ;
    oai21 ix4982 (.Y (nx4981), .A0 (nx7739), .A1 (nx8022), .B0 (nx7741)) ;
    dff L0_0_L1_3_Fij_reg_Dout_4 (.Q (FilterDout_0__3__4), .QB (nx7739), .D (
        nx4981), .CLK (CLK)) ;
    oai21 ix4992 (.Y (nx4991), .A0 (nx7745), .A1 (nx8022), .B0 (nx7747)) ;
    dff L0_0_L1_3_Fij_reg_Dout_5 (.Q (FilterDout_0__3__5), .QB (nx7745), .D (
        nx4991), .CLK (CLK)) ;
    oai21 ix5002 (.Y (nx5001), .A0 (nx7751), .A1 (nx8022), .B0 (nx7753)) ;
    dff L0_0_L1_3_Fij_reg_Dout_6 (.Q (FilterDout_0__3__6), .QB (nx7751), .D (
        nx5001), .CLK (CLK)) ;
    oai21 ix5012 (.Y (nx5011), .A0 (nx7757), .A1 (nx8022), .B0 (nx7759)) ;
    dff L0_0_L1_3_Fij_reg_Dout_7 (.Q (FilterDout_0__3__7), .QB (nx7757), .D (
        nx5011), .CLK (CLK)) ;
    oai21 ix5262 (.Y (nx5261), .A0 (nx7763), .A1 (nx8024), .B0 (nx7765)) ;
    dff L0_0_L1_2_Fij_reg_Dout_0 (.Q (FilterDout_0__2__0), .QB (nx7763), .D (
        nx5261), .CLK (CLK)) ;
    oai21 ix5272 (.Y (nx5271), .A0 (nx7769), .A1 (nx8024), .B0 (nx7771)) ;
    dff L0_0_L1_2_Fij_reg_Dout_1 (.Q (FilterDout_0__2__1), .QB (nx7769), .D (
        nx5271), .CLK (CLK)) ;
    oai21 ix5282 (.Y (nx5281), .A0 (nx7775), .A1 (nx8024), .B0 (nx7777)) ;
    dff L0_0_L1_2_Fij_reg_Dout_2 (.Q (FilterDout_0__2__2), .QB (nx7775), .D (
        nx5281), .CLK (CLK)) ;
    oai21 ix5292 (.Y (nx5291), .A0 (nx7781), .A1 (nx8026), .B0 (nx7783)) ;
    dff L0_0_L1_2_Fij_reg_Dout_3 (.Q (FilterDout_0__2__3), .QB (nx7781), .D (
        nx5291), .CLK (CLK)) ;
    oai21 ix5302 (.Y (nx5301), .A0 (nx7787), .A1 (nx8026), .B0 (nx7789)) ;
    dff L0_0_L1_2_Fij_reg_Dout_4 (.Q (FilterDout_0__2__4), .QB (nx7787), .D (
        nx5301), .CLK (CLK)) ;
    oai21 ix5312 (.Y (nx5311), .A0 (nx7793), .A1 (nx8026), .B0 (nx7795)) ;
    dff L0_0_L1_2_Fij_reg_Dout_5 (.Q (FilterDout_0__2__5), .QB (nx7793), .D (
        nx5311), .CLK (CLK)) ;
    oai21 ix5322 (.Y (nx5321), .A0 (nx7799), .A1 (nx8026), .B0 (nx7801)) ;
    dff L0_0_L1_2_Fij_reg_Dout_6 (.Q (FilterDout_0__2__6), .QB (nx7799), .D (
        nx5321), .CLK (CLK)) ;
    oai21 ix5332 (.Y (nx5331), .A0 (nx7805), .A1 (nx8028), .B0 (nx7807)) ;
    dff L0_0_L1_2_Fij_reg_Dout_7 (.Q (FilterDout_0__2__7), .QB (nx7805), .D (
        nx5331), .CLK (CLK)) ;
    oai21 ix5582 (.Y (nx5581), .A0 (nx7811), .A1 (nx8028), .B0 (nx7813)) ;
    dff L0_0_L1_1_Fij_reg_Dout_0 (.Q (FilterDout_0__1__0), .QB (nx7811), .D (
        nx5581), .CLK (CLK)) ;
    oai21 ix5592 (.Y (nx5591), .A0 (nx7817), .A1 (nx8028), .B0 (nx7819)) ;
    dff L0_0_L1_1_Fij_reg_Dout_1 (.Q (FilterDout_0__1__1), .QB (nx7817), .D (
        nx5591), .CLK (CLK)) ;
    oai21 ix5602 (.Y (nx5601), .A0 (nx7823), .A1 (nx8030), .B0 (nx7825)) ;
    dff L0_0_L1_1_Fij_reg_Dout_2 (.Q (FilterDout_0__1__2), .QB (nx7823), .D (
        nx5601), .CLK (CLK)) ;
    oai21 ix5612 (.Y (nx5611), .A0 (nx7829), .A1 (nx8030), .B0 (nx7831)) ;
    dff L0_0_L1_1_Fij_reg_Dout_3 (.Q (FilterDout_0__1__3), .QB (nx7829), .D (
        nx5611), .CLK (CLK)) ;
    oai21 ix5622 (.Y (nx5621), .A0 (nx7835), .A1 (nx8030), .B0 (nx7837)) ;
    dff L0_0_L1_1_Fij_reg_Dout_4 (.Q (FilterDout_0__1__4), .QB (nx7835), .D (
        nx5621), .CLK (CLK)) ;
    oai21 ix5632 (.Y (nx5631), .A0 (nx7841), .A1 (nx8030), .B0 (nx7843)) ;
    dff L0_0_L1_1_Fij_reg_Dout_5 (.Q (FilterDout_0__1__5), .QB (nx7841), .D (
        nx5631), .CLK (CLK)) ;
    oai21 ix5642 (.Y (nx5641), .A0 (nx7847), .A1 (nx8032), .B0 (nx7849)) ;
    dff L0_0_L1_1_Fij_reg_Dout_6 (.Q (FilterDout_0__1__6), .QB (nx7847), .D (
        nx5641), .CLK (CLK)) ;
    oai21 ix5652 (.Y (nx5651), .A0 (nx7853), .A1 (nx8032), .B0 (nx7855)) ;
    dff L0_0_L1_1_Fij_reg_Dout_7 (.Q (FilterDout_0__1__7), .QB (nx7853), .D (
        nx5651), .CLK (CLK)) ;
    oai21 ix5902 (.Y (nx5901), .A0 (nx7859), .A1 (nx8032), .B0 (nx7861)) ;
    dff L0_0_L1_0_Fij_reg_Dout_0 (.Q (FilterDout_0__0__0), .QB (nx7859), .D (
        nx5901), .CLK (CLK)) ;
    oai21 ix5912 (.Y (nx5911), .A0 (nx7865), .A1 (nx8034), .B0 (nx7867)) ;
    dff L0_0_L1_0_Fij_reg_Dout_1 (.Q (FilterDout_0__0__1), .QB (nx7865), .D (
        nx5911), .CLK (CLK)) ;
    oai21 ix5922 (.Y (nx5921), .A0 (nx7871), .A1 (nx8034), .B0 (nx7873)) ;
    dff L0_0_L1_0_Fij_reg_Dout_2 (.Q (FilterDout_0__0__2), .QB (nx7871), .D (
        nx5921), .CLK (CLK)) ;
    oai21 ix5932 (.Y (nx5931), .A0 (nx7877), .A1 (nx8034), .B0 (nx7879)) ;
    dff L0_0_L1_0_Fij_reg_Dout_3 (.Q (FilterDout_0__0__3), .QB (nx7877), .D (
        nx5931), .CLK (CLK)) ;
    oai21 ix5942 (.Y (nx5941), .A0 (nx7883), .A1 (nx8034), .B0 (nx7885)) ;
    dff L0_0_L1_0_Fij_reg_Dout_4 (.Q (FilterDout_0__0__4), .QB (nx7883), .D (
        nx5941), .CLK (CLK)) ;
    oai21 ix5952 (.Y (nx5951), .A0 (nx7889), .A1 (nx8036), .B0 (nx7891)) ;
    dff L0_0_L1_0_Fij_reg_Dout_5 (.Q (FilterDout_0__0__5), .QB (nx7889), .D (
        nx5951), .CLK (CLK)) ;
    oai21 ix5962 (.Y (nx5961), .A0 (nx7895), .A1 (nx8036), .B0 (nx7897)) ;
    dff L0_0_L1_0_Fij_reg_Dout_6 (.Q (FilterDout_0__0__6), .QB (nx7895), .D (
        nx5961), .CLK (CLK)) ;
    oai21 ix5972 (.Y (nx5971), .A0 (nx7901), .A1 (nx8036), .B0 (nx7903)) ;
    dff L0_0_L1_0_Fij_reg_Dout_7 (.Q (FilterDout_0__0__7), .QB (nx7901), .D (
        nx5971), .CLK (CLK)) ;
    inv02 ix167 (.Y (nx166), .A (nx6966)) ;
    inv02 ix83 (.Y (nx82), .A (nx6008)) ;
    inv02 ix7909 (.Y (nx7910), .A (nx8042)) ;
    inv02 ix7911 (.Y (nx7912), .A (nx8042)) ;
    inv02 ix7913 (.Y (nx7914), .A (nx8042)) ;
    inv02 ix7915 (.Y (nx7916), .A (nx8042)) ;
    inv02 ix7917 (.Y (nx7918), .A (nx8042)) ;
    inv02 ix7919 (.Y (nx7920), .A (nx8244)) ;
    inv02 ix7921 (.Y (nx7922), .A (nx8244)) ;
    inv02 ix7923 (.Y (nx7924), .A (nx8244)) ;
    inv02 ix7925 (.Y (nx7926), .A (nx8244)) ;
    inv02 ix7927 (.Y (nx7928), .A (nx8244)) ;
    inv02 ix7929 (.Y (nx7930), .A (nx8244)) ;
    inv02 ix7931 (.Y (nx7932), .A (nx8244)) ;
    inv02 ix7933 (.Y (nx7934), .A (nx8252)) ;
    inv02 ix7935 (.Y (nx7936), .A (nx8252)) ;
    inv02 ix7937 (.Y (nx7938), .A (nx8252)) ;
    inv02 ix7939 (.Y (nx7940), .A (nx8252)) ;
    inv02 ix7941 (.Y (nx7942), .A (nx8252)) ;
    inv02 ix7943 (.Y (nx7944), .A (nx8252)) ;
    inv02 ix7945 (.Y (nx7946), .A (nx8252)) ;
    inv02 ix7947 (.Y (nx7948), .A (nx8254)) ;
    inv02 ix7949 (.Y (nx7950), .A (nx8254)) ;
    inv02 ix7951 (.Y (nx7952), .A (nx8254)) ;
    inv02 ix7953 (.Y (nx7954), .A (nx8254)) ;
    inv02 ix7955 (.Y (nx7956), .A (nx8254)) ;
    inv02 ix7957 (.Y (nx7958), .A (nx8254)) ;
    inv02 ix7959 (.Y (nx7960), .A (nx8254)) ;
    inv02 ix7961 (.Y (nx7962), .A (nx8260)) ;
    inv02 ix7963 (.Y (nx7964), .A (nx8260)) ;
    inv02 ix7965 (.Y (nx7966), .A (nx8260)) ;
    inv02 ix7967 (.Y (nx7968), .A (nx8260)) ;
    inv02 ix7969 (.Y (nx7970), .A (nx8260)) ;
    inv02 ix7971 (.Y (nx7972), .A (nx8260)) ;
    inv02 ix7973 (.Y (nx7974), .A (nx8186)) ;
    inv02 ix7975 (.Y (nx7976), .A (nx8186)) ;
    inv02 ix7977 (.Y (nx7978), .A (nx8186)) ;
    inv02 ix7979 (.Y (nx7980), .A (nx8186)) ;
    inv02 ix7981 (.Y (nx7982), .A (nx8186)) ;
    inv02 ix7983 (.Y (nx7984), .A (nx8266)) ;
    inv02 ix7985 (.Y (nx7986), .A (nx8266)) ;
    inv02 ix7987 (.Y (nx7988), .A (nx8266)) ;
    inv02 ix7989 (.Y (nx7990), .A (nx8266)) ;
    inv02 ix7991 (.Y (nx7992), .A (nx8266)) ;
    inv02 ix7993 (.Y (nx7994), .A (nx8266)) ;
    inv02 ix7995 (.Y (nx7996), .A (nx8266)) ;
    inv02 ix7997 (.Y (nx7998), .A (nx8274)) ;
    inv02 ix7999 (.Y (nx8000), .A (nx8274)) ;
    inv02 ix8001 (.Y (nx8002), .A (nx8274)) ;
    inv02 ix8003 (.Y (nx8004), .A (nx8274)) ;
    inv02 ix8005 (.Y (nx8006), .A (nx8274)) ;
    inv02 ix8007 (.Y (nx8008), .A (nx8274)) ;
    inv02 ix8009 (.Y (nx8010), .A (nx8274)) ;
    inv02 ix8011 (.Y (nx8012), .A (nx8276)) ;
    inv02 ix8013 (.Y (nx8014), .A (nx8276)) ;
    inv02 ix8015 (.Y (nx8016), .A (nx8276)) ;
    inv02 ix8017 (.Y (nx8018), .A (nx8276)) ;
    inv02 ix8019 (.Y (nx8020), .A (nx8276)) ;
    inv02 ix8021 (.Y (nx8022), .A (nx8276)) ;
    inv02 ix8023 (.Y (nx8024), .A (nx8276)) ;
    inv02 ix8025 (.Y (nx8026), .A (nx8282)) ;
    inv02 ix8027 (.Y (nx8028), .A (nx8282)) ;
    inv02 ix8029 (.Y (nx8030), .A (nx8282)) ;
    inv02 ix8031 (.Y (nx8032), .A (nx8282)) ;
    inv02 ix8033 (.Y (nx8034), .A (nx8282)) ;
    inv02 ix8035 (.Y (nx8036), .A (nx8282)) ;
    inv02 ix8041 (.Y (nx8042), .A (nx8288)) ;
    inv02 ix8043 (.Y (nx8044), .A (nx8288)) ;
    inv02 ix8045 (.Y (nx8046), .A (nx8288)) ;
    inv02 ix8047 (.Y (nx8048), .A (nx8288)) ;
    inv02 ix8049 (.Y (nx8050), .A (nx8288)) ;
    inv02 ix8051 (.Y (nx8052), .A (RST)) ;
    inv02 ix8053 (.Y (nx8054), .A (RST)) ;
    inv02 ix8055 (.Y (nx8056), .A (RST)) ;
    inv02 ix8057 (.Y (nx8058), .A (RST)) ;
    inv02 ix8059 (.Y (nx8060), .A (RST)) ;
    inv02 ix8061 (.Y (nx8062), .A (RST)) ;
    inv02 ix8063 (.Y (nx8064), .A (RST)) ;
    inv02 ix8065 (.Y (nx8066), .A (RST)) ;
    inv02 ix8067 (.Y (nx8068), .A (RST)) ;
    inv02 ix8069 (.Y (nx8070), .A (RST)) ;
    inv02 ix8073 (.Y (nx8074), .A (RST)) ;
    inv02 ix8075 (.Y (nx8076), .A (RST)) ;
    inv02 ix8077 (.Y (nx8078), .A (RST)) ;
    inv02 ix8079 (.Y (nx8080), .A (RST)) ;
    inv02 ix8085 (.Y (nx8086), .A (RST)) ;
    inv02 ix8087 (.Y (nx8088), .A (RST)) ;
    inv02 ix8089 (.Y (nx8090), .A (RST)) ;
    inv02 ix8091 (.Y (nx8092), .A (RST)) ;
    inv02 ix8103 (.Y (nx8104), .A (RST)) ;
    inv02 ix8105 (.Y (nx8106), .A (RST)) ;
    inv02 ix8107 (.Y (nx8108), .A (RST)) ;
    inv02 ix8109 (.Y (nx8110), .A (RST)) ;
    inv02 ix8111 (.Y (nx8112), .A (RST)) ;
    inv02 ix8113 (.Y (nx8114), .A (RST)) ;
    inv02 ix8115 (.Y (nx8116), .A (RST)) ;
    inv02 ix8117 (.Y (nx8118), .A (RST)) ;
    inv02 ix8119 (.Y (nx8120), .A (RST)) ;
    inv02 ix8121 (.Y (nx8122), .A (RST)) ;
    inv02 ix8125 (.Y (nx8126), .A (RST)) ;
    inv02 ix8127 (.Y (nx8128), .A (RST)) ;
    inv02 ix8129 (.Y (nx8130), .A (RST)) ;
    inv02 ix8131 (.Y (nx8132), .A (RST)) ;
    inv02 ix8133 (.Y (nx8134), .A (RST)) ;
    inv02 ix8137 (.Y (nx8138), .A (RST)) ;
    inv02 ix8139 (.Y (nx8140), .A (RST)) ;
    inv02 ix8141 (.Y (nx8142), .A (RST)) ;
    inv02 ix8143 (.Y (nx8144), .A (RST)) ;
    inv02 ix8159 (.Y (nx8160), .A (nx8220)) ;
    inv02 ix8161 (.Y (nx8162), .A (nx8220)) ;
    inv02 ix8163 (.Y (nx8164), .A (nx8220)) ;
    inv02 ix8165 (.Y (nx8166), .A (nx8220)) ;
    inv02 ix8167 (.Y (nx8168), .A (nx8220)) ;
    inv02 ix8169 (.Y (nx8170), .A (nx8220)) ;
    inv02 ix8171 (.Y (nx8172), .A (nx8220)) ;
    inv02 ix8173 (.Y (nx8174), .A (nx8222)) ;
    inv02 ix8175 (.Y (nx8176), .A (nx8222)) ;
    inv02 ix8177 (.Y (nx8178), .A (nx8222)) ;
    inv02 ix8179 (.Y (nx8180), .A (nx8222)) ;
    inv02 ix8185 (.Y (nx8186), .A (nx8292)) ;
    inv02 ix8187 (.Y (nx8188), .A (nx8292)) ;
    inv02 ix8189 (.Y (nx8190), .A (nx8292)) ;
    inv02 ix8191 (.Y (nx8192), .A (nx8292)) ;
    inv02 ix8193 (.Y (nx8194), .A (nx8292)) ;
    inv02 ix8197 (.Y (nx8198), .A (nx8224)) ;
    inv02 ix8199 (.Y (nx8200), .A (nx8224)) ;
    inv02 ix8201 (.Y (nx8202), .A (nx8224)) ;
    inv02 ix8203 (.Y (nx8204), .A (nx8224)) ;
    inv02 ix8205 (.Y (nx8206), .A (nx8224)) ;
    inv02 ix8207 (.Y (nx8208), .A (nx8224)) ;
    inv02 ix8209 (.Y (nx8210), .A (nx8224)) ;
    inv02 ix8211 (.Y (nx8212), .A (nx8226)) ;
    inv02 ix8213 (.Y (nx8214), .A (nx8226)) ;
    inv02 ix8215 (.Y (nx8216), .A (nx8226)) ;
    inv02 ix8217 (.Y (nx8218), .A (nx8226)) ;
    inv02 ix8219 (.Y (nx8220), .A (nx6075)) ;
    inv02 ix8221 (.Y (nx8222), .A (nx6075)) ;
    inv02 ix8223 (.Y (nx8224), .A (nx7016)) ;
    inv02 ix8225 (.Y (nx8226), .A (nx7016)) ;
    mux21_ni ix1982 (.Y (nx1981), .A0 (WindowDout_4__4__0), .A1 (nx86), .S0 (
             nx8288)) ;
    mux21_ni ix1992 (.Y (nx1991), .A0 (WindowDout_4__4__1), .A1 (nx96), .S0 (
             nx8288)) ;
    mux21_ni ix2002 (.Y (nx2001), .A0 (WindowDout_4__4__2), .A1 (nx106), .S0 (
             nx8238)) ;
    mux21_ni ix2012 (.Y (nx2011), .A0 (WindowDout_4__4__3), .A1 (nx116), .S0 (
             nx8238)) ;
    mux21_ni ix2022 (.Y (nx2021), .A0 (WindowDout_4__4__4), .A1 (nx126), .S0 (
             nx8238)) ;
    mux21_ni ix2032 (.Y (nx2031), .A0 (WindowDout_4__4__5), .A1 (nx136), .S0 (
             nx8238)) ;
    mux21_ni ix2042 (.Y (nx2041), .A0 (WindowDout_4__4__6), .A1 (nx146), .S0 (
             nx8238)) ;
    mux21_ni ix2052 (.Y (nx2051), .A0 (WindowDout_4__4__7), .A1 (nx156), .S0 (
             nx8238)) ;
    mux21_ni ix2142 (.Y (nx2141), .A0 (WindowDout_4__3__0), .A1 (nx218), .S0 (
             nx8238)) ;
    mux21_ni ix2152 (.Y (nx2151), .A0 (WindowDout_4__3__1), .A1 (nx228), .S0 (
             nx82)) ;
    mux21_ni ix2162 (.Y (nx2161), .A0 (WindowDout_4__3__2), .A1 (nx238), .S0 (
             nx82)) ;
    mux21_ni ix2172 (.Y (nx2171), .A0 (WindowDout_4__3__3), .A1 (nx248), .S0 (
             nx82)) ;
    mux21_ni ix2182 (.Y (nx2181), .A0 (WindowDout_4__3__4), .A1 (nx258), .S0 (
             nx82)) ;
    mux21_ni ix2192 (.Y (nx2191), .A0 (WindowDout_4__3__5), .A1 (nx268), .S0 (
             nx82)) ;
    mux21_ni ix2202 (.Y (nx2201), .A0 (WindowDout_4__3__6), .A1 (nx278), .S0 (
             nx82)) ;
    mux21_ni ix2212 (.Y (nx2211), .A0 (WindowDout_4__3__7), .A1 (nx288), .S0 (
             nx82)) ;
    or03 ix6321 (.Y (nx6320), .A0 (RST), .A1 (nx6149), .A2 (nx8042)) ;
    or03 ix6327 (.Y (nx6326), .A0 (RST), .A1 (nx6156), .A2 (nx8246)) ;
    or03 ix6333 (.Y (nx6332), .A0 (RST), .A1 (nx6162), .A2 (nx8246)) ;
    or03 ix6339 (.Y (nx6338), .A0 (RST), .A1 (nx6168), .A2 (nx8246)) ;
    or03 ix6345 (.Y (nx6344), .A0 (RST), .A1 (nx6174), .A2 (nx8246)) ;
    or03 ix6351 (.Y (nx6350), .A0 (RST), .A1 (nx6180), .A2 (nx8246)) ;
    or03 ix6357 (.Y (nx6356), .A0 (RST), .A1 (nx6186), .A2 (nx8246)) ;
    or03 ix6363 (.Y (nx6362), .A0 (RST), .A1 (nx6192), .A2 (nx8246)) ;
    or03 ix6369 (.Y (nx6368), .A0 (RST), .A1 (nx6198), .A2 (nx8248)) ;
    or03 ix6375 (.Y (nx6374), .A0 (RST), .A1 (nx6204), .A2 (nx8248)) ;
    or03 ix6381 (.Y (nx6380), .A0 (RST), .A1 (nx6210), .A2 (nx8248)) ;
    or03 ix6387 (.Y (nx6386), .A0 (RST), .A1 (nx6216), .A2 (nx8248)) ;
    or03 ix6393 (.Y (nx6392), .A0 (RST), .A1 (nx6222), .A2 (nx8248)) ;
    or03 ix6399 (.Y (nx6398), .A0 (RST), .A1 (nx6228), .A2 (nx8248)) ;
    or03 ix6405 (.Y (nx6404), .A0 (RST), .A1 (nx6234), .A2 (nx8248)) ;
    or03 ix6411 (.Y (nx6410), .A0 (RST), .A1 (nx6240), .A2 (nx8250)) ;
    or03 ix6489 (.Y (nx6488), .A0 (RST), .A1 (nx6318), .A2 (nx8250)) ;
    or03 ix6495 (.Y (nx6494), .A0 (RST), .A1 (nx6324), .A2 (nx8250)) ;
    or03 ix6501 (.Y (nx6500), .A0 (RST), .A1 (nx6330), .A2 (nx8250)) ;
    or03 ix6507 (.Y (nx6506), .A0 (RST), .A1 (nx6336), .A2 (nx8250)) ;
    or03 ix6513 (.Y (nx6512), .A0 (RST), .A1 (nx6342), .A2 (nx8250)) ;
    or03 ix6519 (.Y (nx6518), .A0 (RST), .A1 (nx6348), .A2 (nx8250)) ;
    or03 ix6525 (.Y (nx6524), .A0 (RST), .A1 (nx6354), .A2 (nx8044)) ;
    or03 ix6531 (.Y (nx6530), .A0 (RST), .A1 (nx6360), .A2 (nx8044)) ;
    or03 ix6537 (.Y (nx6536), .A0 (RST), .A1 (nx6366), .A2 (nx8044)) ;
    or03 ix6543 (.Y (nx6542), .A0 (RST), .A1 (nx6372), .A2 (nx8044)) ;
    or03 ix6549 (.Y (nx6548), .A0 (RST), .A1 (nx6378), .A2 (nx8046)) ;
    or03 ix6555 (.Y (nx6554), .A0 (RST), .A1 (nx6384), .A2 (nx8046)) ;
    or03 ix6561 (.Y (nx6560), .A0 (RST), .A1 (nx6390), .A2 (nx8046)) ;
    or03 ix6567 (.Y (nx6566), .A0 (RST), .A1 (nx6396), .A2 (nx8046)) ;
    or03 ix6573 (.Y (nx6572), .A0 (RST), .A1 (nx6402), .A2 (nx8046)) ;
    or03 ix6579 (.Y (nx6578), .A0 (RST), .A1 (nx6408), .A2 (nx8046)) ;
    or03 ix6729 (.Y (nx6728), .A0 (RST), .A1 (nx6486), .A2 (nx8256)) ;
    or03 ix6735 (.Y (nx6734), .A0 (RST), .A1 (nx6492), .A2 (nx8256)) ;
    or03 ix6741 (.Y (nx6740), .A0 (RST), .A1 (nx6498), .A2 (nx8256)) ;
    or03 ix6747 (.Y (nx6746), .A0 (RST), .A1 (nx6504), .A2 (nx8256)) ;
    or03 ix6753 (.Y (nx6752), .A0 (RST), .A1 (nx6510), .A2 (nx8256)) ;
    or03 ix6759 (.Y (nx6758), .A0 (RST), .A1 (nx6516), .A2 (nx8256)) ;
    or03 ix6765 (.Y (nx6764), .A0 (RST), .A1 (nx6522), .A2 (nx8256)) ;
    or03 ix6771 (.Y (nx6770), .A0 (RST), .A1 (nx6528), .A2 (nx8258)) ;
    or03 ix6777 (.Y (nx6776), .A0 (RST), .A1 (nx6534), .A2 (nx8258)) ;
    or03 ix6783 (.Y (nx6782), .A0 (RST), .A1 (nx6540), .A2 (nx8258)) ;
    or03 ix6789 (.Y (nx6788), .A0 (RST), .A1 (nx6546), .A2 (nx8258)) ;
    or03 ix6795 (.Y (nx6794), .A0 (RST), .A1 (nx6552), .A2 (nx8258)) ;
    or03 ix6801 (.Y (nx6800), .A0 (RST), .A1 (nx6558), .A2 (nx8258)) ;
    or03 ix6807 (.Y (nx6806), .A0 (RST), .A1 (nx6564), .A2 (nx8258)) ;
    or03 ix6813 (.Y (nx6812), .A0 (RST), .A1 (nx6570), .A2 (nx8048)) ;
    or03 ix6819 (.Y (nx6818), .A0 (RST), .A1 (nx6576), .A2 (nx8048)) ;
    or03 ix6825 (.Y (nx6824), .A0 (RST), .A1 (nx6582), .A2 (nx8048)) ;
    or03 ix6831 (.Y (nx6830), .A0 (RST), .A1 (nx6588), .A2 (nx8048)) ;
    or03 ix6837 (.Y (nx6836), .A0 (RST), .A1 (nx6594), .A2 (nx8048)) ;
    or03 ix6843 (.Y (nx6842), .A0 (RST), .A1 (nx6600), .A2 (nx8260)) ;
    or03 ix6849 (.Y (nx6848), .A0 (RST), .A1 (nx6606), .A2 (nx8262)) ;
    or03 ix6855 (.Y (nx6854), .A0 (RST), .A1 (nx6612), .A2 (nx8262)) ;
    or03 ix6861 (.Y (nx6860), .A0 (RST), .A1 (nx6618), .A2 (nx8262)) ;
    or03 ix6867 (.Y (nx6866), .A0 (RST), .A1 (nx6624), .A2 (nx8262)) ;
    or03 ix6873 (.Y (nx6872), .A0 (RST), .A1 (nx6630), .A2 (nx8262)) ;
    or03 ix6879 (.Y (nx6878), .A0 (RST), .A1 (nx6636), .A2 (nx8262)) ;
    or03 ix6885 (.Y (nx6884), .A0 (RST), .A1 (nx6642), .A2 (nx8262)) ;
    or03 ix6891 (.Y (nx6890), .A0 (RST), .A1 (nx6648), .A2 (nx8264)) ;
    or03 ix6897 (.Y (nx6896), .A0 (RST), .A1 (nx6654), .A2 (nx8264)) ;
    or03 ix6903 (.Y (nx6902), .A0 (RST), .A1 (nx6660), .A2 (nx8264)) ;
    or03 ix6909 (.Y (nx6908), .A0 (RST), .A1 (nx6666), .A2 (nx8264)) ;
    or03 ix6915 (.Y (nx6914), .A0 (RST), .A1 (nx6672), .A2 (nx8264)) ;
    or03 ix6921 (.Y (nx6920), .A0 (RST), .A1 (nx6678), .A2 (nx8264)) ;
    or03 ix6927 (.Y (nx6926), .A0 (RST), .A1 (nx6684), .A2 (nx8264)) ;
    or03 ix6933 (.Y (nx6932), .A0 (RST), .A1 (nx6690), .A2 (nx8050)) ;
    or03 ix6939 (.Y (nx6938), .A0 (RST), .A1 (nx6696), .A2 (nx8050)) ;
    or03 ix6945 (.Y (nx6944), .A0 (RST), .A1 (nx6702), .A2 (nx8050)) ;
    or03 ix6951 (.Y (nx6950), .A0 (RST), .A1 (nx6708), .A2 (nx8050)) ;
    or03 ix6957 (.Y (nx6956), .A0 (RST), .A1 (nx6714), .A2 (nx8050)) ;
    or03 ix6963 (.Y (nx6962), .A0 (RST), .A1 (nx6720), .A2 (nx8050)) ;
    mux21_ni ix2062 (.Y (nx2061), .A0 (FilterDout_4__4__0), .A1 (nx86), .S0 (
             nx8292)) ;
    mux21_ni ix2072 (.Y (nx2071), .A0 (FilterDout_4__4__1), .A1 (nx96), .S0 (
             nx8292)) ;
    mux21_ni ix2082 (.Y (nx2081), .A0 (FilterDout_4__4__2), .A1 (nx106), .S0 (
             nx8242)) ;
    mux21_ni ix2092 (.Y (nx2091), .A0 (FilterDout_4__4__3), .A1 (nx116), .S0 (
             nx8242)) ;
    mux21_ni ix2102 (.Y (nx2101), .A0 (FilterDout_4__4__4), .A1 (nx126), .S0 (
             nx8242)) ;
    mux21_ni ix2112 (.Y (nx2111), .A0 (FilterDout_4__4__5), .A1 (nx136), .S0 (
             nx8242)) ;
    mux21_ni ix2122 (.Y (nx2121), .A0 (FilterDout_4__4__6), .A1 (nx146), .S0 (
             nx8242)) ;
    mux21_ni ix2132 (.Y (nx2131), .A0 (FilterDout_4__4__7), .A1 (nx156), .S0 (
             nx8242)) ;
    mux21_ni ix2222 (.Y (nx2221), .A0 (FilterDout_4__3__0), .A1 (nx218), .S0 (
             nx8242)) ;
    mux21_ni ix2232 (.Y (nx2231), .A0 (FilterDout_4__3__1), .A1 (nx228), .S0 (
             nx166)) ;
    mux21_ni ix2242 (.Y (nx2241), .A0 (FilterDout_4__3__2), .A1 (nx238), .S0 (
             nx166)) ;
    mux21_ni ix2252 (.Y (nx2251), .A0 (FilterDout_4__3__3), .A1 (nx248), .S0 (
             nx166)) ;
    mux21_ni ix2262 (.Y (nx2261), .A0 (FilterDout_4__3__4), .A1 (nx258), .S0 (
             nx166)) ;
    mux21_ni ix2272 (.Y (nx2271), .A0 (FilterDout_4__3__5), .A1 (nx268), .S0 (
             nx166)) ;
    mux21_ni ix2282 (.Y (nx2281), .A0 (FilterDout_4__3__6), .A1 (nx278), .S0 (
             nx166)) ;
    mux21_ni ix2292 (.Y (nx2291), .A0 (FilterDout_4__3__7), .A1 (nx288), .S0 (
             nx166)) ;
    or03 ix7262 (.Y (nx7261), .A0 (RST), .A1 (nx7090), .A2 (nx8186)) ;
    or03 ix7268 (.Y (nx7267), .A0 (RST), .A1 (nx7097), .A2 (nx8268)) ;
    or03 ix7274 (.Y (nx7273), .A0 (RST), .A1 (nx7103), .A2 (nx8268)) ;
    or03 ix7280 (.Y (nx7279), .A0 (RST), .A1 (nx7109), .A2 (nx8268)) ;
    or03 ix7286 (.Y (nx7285), .A0 (RST), .A1 (nx7115), .A2 (nx8268)) ;
    or03 ix7292 (.Y (nx7291), .A0 (RST), .A1 (nx7121), .A2 (nx8268)) ;
    or03 ix7298 (.Y (nx7297), .A0 (RST), .A1 (nx7127), .A2 (nx8268)) ;
    or03 ix7304 (.Y (nx7303), .A0 (RST), .A1 (nx7133), .A2 (nx8268)) ;
    or03 ix7310 (.Y (nx7309), .A0 (RST), .A1 (nx7139), .A2 (nx8270)) ;
    or03 ix7316 (.Y (nx7315), .A0 (RST), .A1 (nx7145), .A2 (nx8270)) ;
    or03 ix7322 (.Y (nx7321), .A0 (RST), .A1 (nx7151), .A2 (nx8270)) ;
    or03 ix7328 (.Y (nx7327), .A0 (RST), .A1 (nx7157), .A2 (nx8270)) ;
    or03 ix7334 (.Y (nx7333), .A0 (RST), .A1 (nx7163), .A2 (nx8270)) ;
    or03 ix7340 (.Y (nx7339), .A0 (RST), .A1 (nx7169), .A2 (nx8270)) ;
    or03 ix7346 (.Y (nx7345), .A0 (RST), .A1 (nx7175), .A2 (nx8270)) ;
    or03 ix7352 (.Y (nx7351), .A0 (RST), .A1 (nx7181), .A2 (nx8272)) ;
    or03 ix7430 (.Y (nx7429), .A0 (RST), .A1 (nx7259), .A2 (nx8272)) ;
    or03 ix7436 (.Y (nx7435), .A0 (RST), .A1 (nx7265), .A2 (nx8272)) ;
    or03 ix7442 (.Y (nx7441), .A0 (RST), .A1 (nx7271), .A2 (nx8272)) ;
    or03 ix7448 (.Y (nx7447), .A0 (RST), .A1 (nx7277), .A2 (nx8272)) ;
    or03 ix7454 (.Y (nx7453), .A0 (RST), .A1 (nx7283), .A2 (nx8272)) ;
    or03 ix7460 (.Y (nx7459), .A0 (RST), .A1 (nx7289), .A2 (nx8272)) ;
    or03 ix7466 (.Y (nx7465), .A0 (RST), .A1 (nx7295), .A2 (nx8188)) ;
    or03 ix7472 (.Y (nx7471), .A0 (RST), .A1 (nx7301), .A2 (nx8188)) ;
    or03 ix7478 (.Y (nx7477), .A0 (RST), .A1 (nx7307), .A2 (nx8188)) ;
    or03 ix7484 (.Y (nx7483), .A0 (RST), .A1 (nx7313), .A2 (nx8188)) ;
    or03 ix7490 (.Y (nx7489), .A0 (RST), .A1 (nx7319), .A2 (nx8190)) ;
    or03 ix7496 (.Y (nx7495), .A0 (RST), .A1 (nx7325), .A2 (nx8190)) ;
    or03 ix7502 (.Y (nx7501), .A0 (RST), .A1 (nx7331), .A2 (nx8190)) ;
    or03 ix7508 (.Y (nx7507), .A0 (RST), .A1 (nx7337), .A2 (nx8190)) ;
    or03 ix7514 (.Y (nx7513), .A0 (RST), .A1 (nx7343), .A2 (nx8190)) ;
    or03 ix7520 (.Y (nx7519), .A0 (RST), .A1 (nx7349), .A2 (nx8190)) ;
    or03 ix7670 (.Y (nx7669), .A0 (RST), .A1 (nx7427), .A2 (nx8278)) ;
    or03 ix7676 (.Y (nx7675), .A0 (RST), .A1 (nx7433), .A2 (nx8278)) ;
    or03 ix7682 (.Y (nx7681), .A0 (RST), .A1 (nx7439), .A2 (nx8278)) ;
    or03 ix7688 (.Y (nx7687), .A0 (RST), .A1 (nx7445), .A2 (nx8278)) ;
    or03 ix7694 (.Y (nx7693), .A0 (RST), .A1 (nx7451), .A2 (nx8278)) ;
    or03 ix7700 (.Y (nx7699), .A0 (RST), .A1 (nx7457), .A2 (nx8278)) ;
    or03 ix7706 (.Y (nx7705), .A0 (RST), .A1 (nx7463), .A2 (nx8278)) ;
    or03 ix7712 (.Y (nx7711), .A0 (RST), .A1 (nx7469), .A2 (nx8280)) ;
    or03 ix7718 (.Y (nx7717), .A0 (RST), .A1 (nx7475), .A2 (nx8280)) ;
    or03 ix7724 (.Y (nx7723), .A0 (RST), .A1 (nx7481), .A2 (nx8280)) ;
    or03 ix7730 (.Y (nx7729), .A0 (RST), .A1 (nx7487), .A2 (nx8280)) ;
    or03 ix7736 (.Y (nx7735), .A0 (RST), .A1 (nx7493), .A2 (nx8280)) ;
    or03 ix7742 (.Y (nx7741), .A0 (RST), .A1 (nx7499), .A2 (nx8280)) ;
    or03 ix7748 (.Y (nx7747), .A0 (RST), .A1 (nx7505), .A2 (nx8280)) ;
    or03 ix7754 (.Y (nx7753), .A0 (RST), .A1 (nx7511), .A2 (nx8192)) ;
    or03 ix7760 (.Y (nx7759), .A0 (RST), .A1 (nx7517), .A2 (nx8192)) ;
    or03 ix7766 (.Y (nx7765), .A0 (RST), .A1 (nx7523), .A2 (nx8192)) ;
    or03 ix7772 (.Y (nx7771), .A0 (RST), .A1 (nx7529), .A2 (nx8192)) ;
    or03 ix7778 (.Y (nx7777), .A0 (RST), .A1 (nx7535), .A2 (nx8192)) ;
    or03 ix7784 (.Y (nx7783), .A0 (RST), .A1 (nx7541), .A2 (nx8282)) ;
    or03 ix7790 (.Y (nx7789), .A0 (RST), .A1 (nx7547), .A2 (nx8284)) ;
    or03 ix7796 (.Y (nx7795), .A0 (RST), .A1 (nx7553), .A2 (nx8284)) ;
    or03 ix7802 (.Y (nx7801), .A0 (RST), .A1 (nx7559), .A2 (nx8284)) ;
    or03 ix7808 (.Y (nx7807), .A0 (RST), .A1 (nx7565), .A2 (nx8284)) ;
    or03 ix7814 (.Y (nx7813), .A0 (RST), .A1 (nx7571), .A2 (nx8284)) ;
    or03 ix7820 (.Y (nx7819), .A0 (RST), .A1 (nx7577), .A2 (nx8284)) ;
    or03 ix7826 (.Y (nx7825), .A0 (RST), .A1 (nx7583), .A2 (nx8284)) ;
    or03 ix7832 (.Y (nx7831), .A0 (RST), .A1 (nx7589), .A2 (nx8286)) ;
    or03 ix7838 (.Y (nx7837), .A0 (RST), .A1 (nx7595), .A2 (nx8286)) ;
    or03 ix7844 (.Y (nx7843), .A0 (RST), .A1 (nx7601), .A2 (nx8286)) ;
    or03 ix7850 (.Y (nx7849), .A0 (RST), .A1 (nx7607), .A2 (nx8286)) ;
    or03 ix7856 (.Y (nx7855), .A0 (RST), .A1 (nx7613), .A2 (nx8286)) ;
    or03 ix7862 (.Y (nx7861), .A0 (RST), .A1 (nx7619), .A2 (nx8286)) ;
    or03 ix7868 (.Y (nx7867), .A0 (RST), .A1 (nx7625), .A2 (nx8286)) ;
    or03 ix7874 (.Y (nx7873), .A0 (RST), .A1 (nx7631), .A2 (nx8194)) ;
    or03 ix7880 (.Y (nx7879), .A0 (RST), .A1 (nx7637), .A2 (nx8194)) ;
    or03 ix7886 (.Y (nx7885), .A0 (RST), .A1 (nx7643), .A2 (nx8194)) ;
    or03 ix7892 (.Y (nx7891), .A0 (RST), .A1 (nx7649), .A2 (nx8194)) ;
    or03 ix7898 (.Y (nx7897), .A0 (RST), .A1 (nx7655), .A2 (nx8194)) ;
    or03 ix7904 (.Y (nx7903), .A0 (RST), .A1 (nx7661), .A2 (nx8194)) ;
    inv02 ix8235 (.Y (nx8236), .A (nx8300)) ;
    inv02 ix8237 (.Y (nx8238), .A (nx8300)) ;
    inv02 ix8239 (.Y (nx8240), .A (nx8302)) ;
    inv02 ix8241 (.Y (nx8242), .A (nx8302)) ;
    inv02 ix8243 (.Y (nx8244), .A (nx8290)) ;
    inv02 ix8245 (.Y (nx8246), .A (nx8290)) ;
    inv02 ix8247 (.Y (nx8248), .A (nx8290)) ;
    inv02 ix8249 (.Y (nx8250), .A (nx8290)) ;
    inv02 ix8251 (.Y (nx8252), .A (nx8290)) ;
    inv02 ix8253 (.Y (nx8254), .A (nx8290)) ;
    inv02 ix8255 (.Y (nx8256), .A (nx8290)) ;
    inv02 ix8257 (.Y (nx8258), .A (nx8236)) ;
    inv02 ix8259 (.Y (nx8260), .A (nx8236)) ;
    inv02 ix8261 (.Y (nx8262), .A (nx8236)) ;
    inv02 ix8263 (.Y (nx8264), .A (nx8236)) ;
    inv02 ix8265 (.Y (nx8266), .A (nx8294)) ;
    inv02 ix8267 (.Y (nx8268), .A (nx8294)) ;
    inv02 ix8269 (.Y (nx8270), .A (nx8294)) ;
    inv02 ix8271 (.Y (nx8272), .A (nx8294)) ;
    inv02 ix8273 (.Y (nx8274), .A (nx8294)) ;
    inv02 ix8275 (.Y (nx8276), .A (nx8294)) ;
    inv02 ix8277 (.Y (nx8278), .A (nx8294)) ;
    inv02 ix8279 (.Y (nx8280), .A (nx8240)) ;
    inv02 ix8281 (.Y (nx8282), .A (nx8240)) ;
    inv02 ix8283 (.Y (nx8284), .A (nx8240)) ;
    inv02 ix8285 (.Y (nx8286), .A (nx8240)) ;
    inv02 ix8287 (.Y (nx8288), .A (nx8300)) ;
    inv02 ix8289 (.Y (nx8290), .A (nx8300)) ;
    inv02 ix8291 (.Y (nx8292), .A (nx8302)) ;
    inv02 ix8293 (.Y (nx8294), .A (nx8302)) ;
    inv01 ix8299 (.Y (nx8300), .A (nx82)) ;
    inv01 ix8301 (.Y (nx8302), .A (nx166)) ;
endmodule

