//
// Verilog description for cell accelerator, 
// Sat May 12 15:09:56 2018
//
// LeonardoSpectrum Level 3, 2017a.2 
//


module accelerator ( CLK, RST, Start, FilterSize, Stride, Instr, Done, MemRD, 
                     MemWR, MemAddr, MemDin, MemDout ) ;

    input CLK ;
    input RST ;
    input Start ;
    input FilterSize ;
    input Stride ;
    input Instr ;
    output Done ;
    output MemRD ;
    output MemWR ;
    output [17:0]MemAddr ;
    output [7:0]MemDin ;
    input [39:0]MemDout ;

    wire FirstCycle, CacheRST, CacheFilterWR, CacheWindowWR, CacheFilter_0__0__7, 
         CacheFilter_0__0__6, CacheFilter_0__0__5, CacheFilter_0__0__4, 
         CacheFilter_0__0__3, CacheFilter_0__0__2, CacheFilter_0__0__1, 
         CacheFilter_0__0__0, CacheFilter_0__1__7, CacheFilter_0__1__6, 
         CacheFilter_0__1__5, CacheFilter_0__1__4, CacheFilter_0__1__3, 
         CacheFilter_0__1__2, CacheFilter_0__1__1, CacheFilter_0__1__0, 
         CacheFilter_0__2__7, CacheFilter_0__2__6, CacheFilter_0__2__5, 
         CacheFilter_0__2__4, CacheFilter_0__2__3, CacheFilter_0__2__2, 
         CacheFilter_0__2__1, CacheFilter_0__2__0, CacheFilter_0__3__7, 
         CacheFilter_0__3__6, CacheFilter_0__3__5, CacheFilter_0__3__4, 
         CacheFilter_0__3__3, CacheFilter_0__3__2, CacheFilter_0__3__1, 
         CacheFilter_0__3__0, CacheFilter_0__4__7, CacheFilter_0__4__6, 
         CacheFilter_0__4__5, CacheFilter_0__4__4, CacheFilter_0__4__3, 
         CacheFilter_0__4__2, CacheFilter_0__4__1, CacheFilter_0__4__0, 
         CacheFilter_1__0__7, CacheFilter_1__0__6, CacheFilter_1__0__5, 
         CacheFilter_1__0__4, CacheFilter_1__0__3, CacheFilter_1__0__2, 
         CacheFilter_1__0__1, CacheFilter_1__0__0, CacheFilter_1__1__7, 
         CacheFilter_1__1__6, CacheFilter_1__1__5, CacheFilter_1__1__4, 
         CacheFilter_1__1__3, CacheFilter_1__1__2, CacheFilter_1__1__1, 
         CacheFilter_1__1__0, CacheFilter_1__2__7, CacheFilter_1__2__6, 
         CacheFilter_1__2__5, CacheFilter_1__2__4, CacheFilter_1__2__3, 
         CacheFilter_1__2__2, CacheFilter_1__2__1, CacheFilter_1__2__0, 
         CacheFilter_1__3__7, CacheFilter_1__3__6, CacheFilter_1__3__5, 
         CacheFilter_1__3__4, CacheFilter_1__3__3, CacheFilter_1__3__2, 
         CacheFilter_1__3__1, CacheFilter_1__3__0, CacheFilter_1__4__7, 
         CacheFilter_1__4__6, CacheFilter_1__4__5, CacheFilter_1__4__4, 
         CacheFilter_1__4__3, CacheFilter_1__4__2, CacheFilter_1__4__1, 
         CacheFilter_1__4__0, CacheFilter_2__0__7, CacheFilter_2__0__6, 
         CacheFilter_2__0__5, CacheFilter_2__0__4, CacheFilter_2__0__3, 
         CacheFilter_2__0__2, CacheFilter_2__0__1, CacheFilter_2__0__0, 
         CacheFilter_2__1__7, CacheFilter_2__1__6, CacheFilter_2__1__5, 
         CacheFilter_2__1__4, CacheFilter_2__1__3, CacheFilter_2__1__2, 
         CacheFilter_2__1__1, CacheFilter_2__1__0, CacheFilter_2__2__7, 
         CacheFilter_2__2__6, CacheFilter_2__2__5, CacheFilter_2__2__4, 
         CacheFilter_2__2__3, CacheFilter_2__2__2, CacheFilter_2__2__1, 
         CacheFilter_2__2__0, CacheFilter_2__3__7, CacheFilter_2__3__6, 
         CacheFilter_2__3__5, CacheFilter_2__3__4, CacheFilter_2__3__3, 
         CacheFilter_2__3__2, CacheFilter_2__3__1, CacheFilter_2__3__0, 
         CacheFilter_2__4__7, CacheFilter_2__4__6, CacheFilter_2__4__5, 
         CacheFilter_2__4__4, CacheFilter_2__4__3, CacheFilter_2__4__2, 
         CacheFilter_2__4__1, CacheFilter_2__4__0, CacheFilter_3__0__7, 
         CacheFilter_3__0__6, CacheFilter_3__0__5, CacheFilter_3__0__4, 
         CacheFilter_3__0__3, CacheFilter_3__0__2, CacheFilter_3__0__1, 
         CacheFilter_3__0__0, CacheFilter_3__1__7, CacheFilter_3__1__6, 
         CacheFilter_3__1__5, CacheFilter_3__1__4, CacheFilter_3__1__3, 
         CacheFilter_3__1__2, CacheFilter_3__1__1, CacheFilter_3__1__0, 
         CacheFilter_3__2__7, CacheFilter_3__2__6, CacheFilter_3__2__5, 
         CacheFilter_3__2__4, CacheFilter_3__2__3, CacheFilter_3__2__2, 
         CacheFilter_3__2__1, CacheFilter_3__2__0, CacheFilter_3__3__7, 
         CacheFilter_3__3__6, CacheFilter_3__3__5, CacheFilter_3__3__4, 
         CacheFilter_3__3__3, CacheFilter_3__3__2, CacheFilter_3__3__1, 
         CacheFilter_3__3__0, CacheFilter_3__4__7, CacheFilter_3__4__6, 
         CacheFilter_3__4__5, CacheFilter_3__4__4, CacheFilter_3__4__3, 
         CacheFilter_3__4__2, CacheFilter_3__4__1, CacheFilter_3__4__0, 
         CacheFilter_4__0__7, CacheFilter_4__0__6, CacheFilter_4__0__5, 
         CacheFilter_4__0__4, CacheFilter_4__0__3, CacheFilter_4__0__2, 
         CacheFilter_4__0__1, CacheFilter_4__0__0, CacheFilter_4__1__7, 
         CacheFilter_4__1__6, CacheFilter_4__1__5, CacheFilter_4__1__4, 
         CacheFilter_4__1__3, CacheFilter_4__1__2, CacheFilter_4__1__1, 
         CacheFilter_4__1__0, CacheFilter_4__2__7, CacheFilter_4__2__6, 
         CacheFilter_4__2__5, CacheFilter_4__2__4, CacheFilter_4__2__3, 
         CacheFilter_4__2__2, CacheFilter_4__2__1, CacheFilter_4__2__0, 
         CacheFilter_4__3__7, CacheFilter_4__3__6, CacheFilter_4__3__5, 
         CacheFilter_4__3__4, CacheFilter_4__3__3, CacheFilter_4__3__2, 
         CacheFilter_4__3__1, CacheFilter_4__3__0, CacheFilter_4__4__7, 
         CacheFilter_4__4__6, CacheFilter_4__4__5, CacheFilter_4__4__4, 
         CacheFilter_4__4__3, CacheFilter_4__4__2, CacheFilter_4__4__1, 
         CacheFilter_4__4__0, CacheWindow_0__0__7, CacheWindow_0__0__6, 
         CacheWindow_0__0__5, CacheWindow_0__0__4, CacheWindow_0__0__3, 
         CacheWindow_0__0__2, CacheWindow_0__0__1, CacheWindow_0__0__0, 
         CacheWindow_0__1__7, CacheWindow_0__1__6, CacheWindow_0__1__5, 
         CacheWindow_0__1__4, CacheWindow_0__1__3, CacheWindow_0__1__2, 
         CacheWindow_0__1__1, CacheWindow_0__1__0, CacheWindow_0__2__7, 
         CacheWindow_0__2__6, CacheWindow_0__2__5, CacheWindow_0__2__4, 
         CacheWindow_0__2__3, CacheWindow_0__2__2, CacheWindow_0__2__1, 
         CacheWindow_0__2__0, CacheWindow_0__3__7, CacheWindow_0__3__6, 
         CacheWindow_0__3__5, CacheWindow_0__3__4, CacheWindow_0__3__3, 
         CacheWindow_0__3__2, CacheWindow_0__3__1, CacheWindow_0__3__0, 
         CacheWindow_0__4__7, CacheWindow_0__4__6, CacheWindow_0__4__5, 
         CacheWindow_0__4__4, CacheWindow_0__4__3, CacheWindow_0__4__2, 
         CacheWindow_0__4__1, CacheWindow_0__4__0, CacheWindow_1__0__7, 
         CacheWindow_1__0__6, CacheWindow_1__0__5, CacheWindow_1__0__4, 
         CacheWindow_1__0__3, CacheWindow_1__0__2, CacheWindow_1__0__1, 
         CacheWindow_1__0__0, CacheWindow_1__1__7, CacheWindow_1__1__6, 
         CacheWindow_1__1__5, CacheWindow_1__1__4, CacheWindow_1__1__3, 
         CacheWindow_1__1__2, CacheWindow_1__1__1, CacheWindow_1__1__0, 
         CacheWindow_1__2__7, CacheWindow_1__2__6, CacheWindow_1__2__5, 
         CacheWindow_1__2__4, CacheWindow_1__2__3, CacheWindow_1__2__2, 
         CacheWindow_1__2__1, CacheWindow_1__2__0, CacheWindow_1__3__7, 
         CacheWindow_1__3__6, CacheWindow_1__3__5, CacheWindow_1__3__4, 
         CacheWindow_1__3__3, CacheWindow_1__3__2, CacheWindow_1__3__1, 
         CacheWindow_1__3__0, CacheWindow_1__4__7, CacheWindow_1__4__6, 
         CacheWindow_1__4__5, CacheWindow_1__4__4, CacheWindow_1__4__3, 
         CacheWindow_1__4__2, CacheWindow_1__4__1, CacheWindow_1__4__0, 
         CacheWindow_2__0__7, CacheWindow_2__0__6, CacheWindow_2__0__5, 
         CacheWindow_2__0__4, CacheWindow_2__0__3, CacheWindow_2__0__2, 
         CacheWindow_2__0__1, CacheWindow_2__0__0, CacheWindow_2__1__7, 
         CacheWindow_2__1__6, CacheWindow_2__1__5, CacheWindow_2__1__4, 
         CacheWindow_2__1__3, CacheWindow_2__1__2, CacheWindow_2__1__1, 
         CacheWindow_2__1__0, CacheWindow_2__2__7, CacheWindow_2__2__6, 
         CacheWindow_2__2__5, CacheWindow_2__2__4, CacheWindow_2__2__3, 
         CacheWindow_2__2__2, CacheWindow_2__2__1, CacheWindow_2__2__0, 
         CacheWindow_2__3__7, CacheWindow_2__3__6, CacheWindow_2__3__5, 
         CacheWindow_2__3__4, CacheWindow_2__3__3, CacheWindow_2__3__2, 
         CacheWindow_2__3__1, CacheWindow_2__3__0, CacheWindow_2__4__7, 
         CacheWindow_2__4__6, CacheWindow_2__4__5, CacheWindow_2__4__4, 
         CacheWindow_2__4__3, CacheWindow_2__4__2, CacheWindow_2__4__1, 
         CacheWindow_2__4__0, CacheWindow_3__0__7, CacheWindow_3__0__6, 
         CacheWindow_3__0__5, CacheWindow_3__0__4, CacheWindow_3__0__3, 
         CacheWindow_3__0__2, CacheWindow_3__0__1, CacheWindow_3__0__0, 
         CacheWindow_3__1__7, CacheWindow_3__1__6, CacheWindow_3__1__5, 
         CacheWindow_3__1__4, CacheWindow_3__1__3, CacheWindow_3__1__2, 
         CacheWindow_3__1__1, CacheWindow_3__1__0, CacheWindow_3__2__7, 
         CacheWindow_3__2__6, CacheWindow_3__2__5, CacheWindow_3__2__4, 
         CacheWindow_3__2__3, CacheWindow_3__2__2, CacheWindow_3__2__1, 
         CacheWindow_3__2__0, CacheWindow_3__3__7, CacheWindow_3__3__6, 
         CacheWindow_3__3__5, CacheWindow_3__3__4, CacheWindow_3__3__3, 
         CacheWindow_3__3__2, CacheWindow_3__3__1, CacheWindow_3__3__0, 
         CacheWindow_3__4__7, CacheWindow_3__4__6, CacheWindow_3__4__5, 
         CacheWindow_3__4__4, CacheWindow_3__4__3, CacheWindow_3__4__2, 
         CacheWindow_3__4__1, CacheWindow_3__4__0, CacheWindow_4__0__7, 
         CacheWindow_4__0__6, CacheWindow_4__0__5, CacheWindow_4__0__4, 
         CacheWindow_4__0__3, CacheWindow_4__0__2, CacheWindow_4__0__1, 
         CacheWindow_4__0__0, CacheWindow_4__1__7, CacheWindow_4__1__6, 
         CacheWindow_4__1__5, CacheWindow_4__1__4, CacheWindow_4__1__3, 
         CacheWindow_4__1__2, CacheWindow_4__1__1, CacheWindow_4__1__0, 
         CacheWindow_4__2__7, CacheWindow_4__2__6, CacheWindow_4__2__5, 
         CacheWindow_4__2__4, CacheWindow_4__2__3, CacheWindow_4__2__2, 
         CacheWindow_4__2__1, CacheWindow_4__2__0, CacheWindow_4__3__7, 
         CacheWindow_4__3__6, CacheWindow_4__3__5, CacheWindow_4__3__4, 
         CacheWindow_4__3__3, CacheWindow_4__3__2, CacheWindow_4__3__1, 
         CacheWindow_4__3__0, CacheWindow_4__4__7, CacheWindow_4__4__6, 
         CacheWindow_4__4__5, CacheWindow_4__4__4, CacheWindow_4__4__3, 
         CacheWindow_4__4__2, CacheWindow_4__4__1, CacheWindow_4__4__0, 
         Calculating, CalcStarted, CalcStartRST, AccStartCalc, AccFinishCalc, 
         PWR, CONTROLLER_NxtState_3, CONTROLLER_NxtState_2, 
         CONTROLLER_NxtState_1, CONTROLLER_NxtState_0, CONTROLLER_Restart, 
         CONTROLLER_CntRST, CONTROLLER_CntEN, CONTROLLER_NxtRow_7, 
         CONTROLLER_NxtRow_6, CONTROLLER_NxtRow_5, CONTROLLER_NxtRow_4, 
         CONTROLLER_NxtRow_3, CONTROLLER_NxtRow_2, CONTROLLER_NxtRow_1, 
         CONTROLLER_NxtRow_0, CONTROLLER_NxtCol_7, CONTROLLER_NxtCol_6, 
         CONTROLLER_NxtCol_5, CONTROLLER_NxtCol_4, CONTROLLER_NxtCol_3, 
         CONTROLLER_NxtCol_2, CONTROLLER_NxtCol_1, CONTROLLER_NxtCol_0, 
         CONTROLLER_CurRow_7, CONTROLLER_CurRow_6, CONTROLLER_CurRow_5, 
         CONTROLLER_CurRow_4, CONTROLLER_CurRow_3, CONTROLLER_CurRow_2, 
         CONTROLLER_CurRow_1, CONTROLLER_CurRow_0, CONTROLLER_CurCol_7, 
         CONTROLLER_CurCol_6, CONTROLLER_CurCol_5, CONTROLLER_CurCol_4, 
         CONTROLLER_CurCol_3, CONTROLLER_CurCol_2, CONTROLLER_CurCol_1, 
         CONTROLLER_CurCol_0, CONTROLLER_NxtState_4, CONTROLLER_FilterAddr_17, 
         CONTROLLER_nx8, CONTROLLER_nx12, CONTROLLER_nx14, CONTROLLER_nx58, 
         CONTROLLER_nx70, CONTROLLER_nx74, CONTROLLER_nx78, CONTROLLER_nx124, 
         CONTROLLER_nx138, CONTROLLER_nx142, CONTROLLER_nx150, CONTROLLER_nx168, 
         CONTROLLER_nx210, CONTROLLER_nx216, CONTROLLER_nx254, CONTROLLER_nx260, 
         CONTROLLER_nx306, CONTROLLER_nx310, CONTROLLER_nx320, CONTROLLER_nx322, 
         CONTROLLER_nx346, CONTROLLER_nx374, CONTROLLER_nx390, CONTROLLER_nx426, 
         CONTROLLER_nx444, CONTROLLER_nx468, CONTROLLER_nx482, CONTROLLER_nx492, 
         CONTROLLER_nx502, CONTROLLER_nx561, CONTROLLER_nx563, CONTROLLER_nx565, 
         CONTROLLER_nx567, CONTROLLER_nx571, CONTROLLER_nx575, CONTROLLER_nx577, 
         CONTROLLER_nx581, CONTROLLER_nx583, CONTROLLER_nx585, CONTROLLER_nx593, 
         CONTROLLER_nx599, CONTROLLER_nx602, CONTROLLER_nx606, CONTROLLER_nx609, 
         CONTROLLER_nx613, CONTROLLER_nx616, CONTROLLER_nx622, CONTROLLER_nx625, 
         CONTROLLER_nx632, CONTROLLER_nx634, CONTROLLER_nx638, CONTROLLER_nx640, 
         CONTROLLER_nx645, CONTROLLER_nx647, CONTROLLER_nx650, CONTROLLER_nx654, 
         CONTROLLER_nx656, CONTROLLER_nx662, CONTROLLER_nx665, CONTROLLER_nx667, 
         CONTROLLER_nx671, CONTROLLER_nx673, CONTROLLER_nx675, CONTROLLER_nx677, 
         CONTROLLER_nx679, CONTROLLER_nx685, CONTROLLER_nx691, CONTROLLER_nx693, 
         CONTROLLER_nx696, CONTROLLER_nx699, CONTROLLER_nx701, CONTROLLER_nx704, 
         CONTROLLER_nx709, CONTROLLER_nx711, CONTROLLER_nx716, CONTROLLER_nx718, 
         CONTROLLER_nx723, CONTROLLER_nx727, CONTROLLER_nx729, CONTROLLER_nx732, 
         CONTROLLER_nx735, CONTROLLER_nx738, CONTROLLER_nx740, CONTROLLER_nx744, 
         CONTROLLER_nx749, CONTROLLER_nx751, CONTROLLER_nx753, CONTROLLER_nx756, 
         CONTROLLER_nx758, CONTROLLER_nx763, CONTROLLER_nx765, CONTROLLER_nx767, 
         CONTROLLER_nx770, CONTROLLER_nx773, CONTROLLER_nx776, CONTROLLER_nx778, 
         CONTROLLER_nx781, CONTROLLER_nx791, CONTROLLER_nx793, CONTROLLER_nx795, 
         CONTROLLER_nx797, CONTROLLER_nx799, CONTROLLER_nx801, CONTROLLER_nx803, 
         CONTROLLER_nx805, CONTROLLER_nx807, CONTROLLER_nx809, CONTROLLER_nx811, 
         CONTROLLER_nx813, CONTROLLER_nx815, CONTROLLER_nx817, CONTROLLER_nx823, 
         CONTROLLER_nx829, CONTROLLER_STATE_NOT_CLK, CONTROLLER_STATE_nx152, 
         CONTROLLER_STATE_nx162, CONTROLLER_STATE_nx172, CONTROLLER_STATE_nx182, 
         CONTROLLER_STATE_nx192, CONTROLLER_STATE_nx206, CONTROLLER_ROW_NOT_CLK, 
         CONTROLLER_ROW_nx212, CONTROLLER_ROW_nx222, CONTROLLER_ROW_nx232, 
         CONTROLLER_ROW_nx242, CONTROLLER_ROW_nx252, CONTROLLER_ROW_nx262, 
         CONTROLLER_ROW_nx272, CONTROLLER_ROW_nx282, CONTROLLER_ROW_nx296, 
         CONTROLLER_ROW_nx327, CONTROLLER_ROW_nx335, CONTROLLER_ROW_nx337, 
         CONTROLLER_COL_NOT_CLK, CONTROLLER_COL_nx212, CONTROLLER_COL_nx222, 
         CONTROLLER_COL_nx232, CONTROLLER_COL_nx242, CONTROLLER_COL_nx252, 
         CONTROLLER_COL_nx262, CONTROLLER_COL_nx272, CONTROLLER_COL_nx282, 
         CONTROLLER_COL_nx296, CONTROLLER_COL_nx327, CONTROLLER_COL_nx335, 
         CONTROLLER_COL_nx337, CALC_FLIP_FLOP_2_NOT_CLK, CALCULATOR_CounterEN, 
         CALCULATOR_CounterRST, CALCULATOR_CalculatingBooth, 
         CALCULATOR_CounterOut_3, CALCULATOR_CounterOut_2, 
         CALCULATOR_CounterOut_1, CALCULATOR_CounterOut_0, 
         CALCULATOR_L1FirstOperands_0__7, CALCULATOR_L1FirstOperands_0__6, 
         CALCULATOR_L1FirstOperands_0__5, CALCULATOR_L1FirstOperands_0__4, 
         CALCULATOR_L1FirstOperands_0__3, CALCULATOR_L1FirstOperands_0__2, 
         CALCULATOR_L1FirstOperands_0__1, CALCULATOR_L1FirstOperands_0__0, 
         CALCULATOR_L1FirstOperands_1__7, CALCULATOR_L1FirstOperands_1__6, 
         CALCULATOR_L1FirstOperands_1__5, CALCULATOR_L1FirstOperands_1__4, 
         CALCULATOR_L1FirstOperands_1__3, CALCULATOR_L1FirstOperands_1__2, 
         CALCULATOR_L1FirstOperands_1__1, CALCULATOR_L1FirstOperands_1__0, 
         CALCULATOR_L1FirstOperands_2__7, CALCULATOR_L1FirstOperands_2__6, 
         CALCULATOR_L1FirstOperands_2__5, CALCULATOR_L1FirstOperands_2__4, 
         CALCULATOR_L1FirstOperands_2__3, CALCULATOR_L1FirstOperands_2__2, 
         CALCULATOR_L1FirstOperands_2__1, CALCULATOR_L1FirstOperands_2__0, 
         CALCULATOR_L1FirstOperands_3__7, CALCULATOR_L1FirstOperands_3__6, 
         CALCULATOR_L1FirstOperands_3__5, CALCULATOR_L1FirstOperands_3__4, 
         CALCULATOR_L1FirstOperands_3__3, CALCULATOR_L1FirstOperands_3__2, 
         CALCULATOR_L1FirstOperands_3__1, CALCULATOR_L1FirstOperands_3__0, 
         CALCULATOR_L1FirstOperands_4__7, CALCULATOR_L1FirstOperands_4__6, 
         CALCULATOR_L1FirstOperands_4__5, CALCULATOR_L1FirstOperands_4__4, 
         CALCULATOR_L1FirstOperands_4__3, CALCULATOR_L1FirstOperands_4__2, 
         CALCULATOR_L1FirstOperands_4__1, CALCULATOR_L1FirstOperands_4__0, 
         CALCULATOR_L1FirstOperands_5__7, CALCULATOR_L1FirstOperands_5__6, 
         CALCULATOR_L1FirstOperands_5__5, CALCULATOR_L1FirstOperands_5__4, 
         CALCULATOR_L1FirstOperands_5__3, CALCULATOR_L1FirstOperands_5__2, 
         CALCULATOR_L1FirstOperands_5__1, CALCULATOR_L1FirstOperands_5__0, 
         CALCULATOR_L1FirstOperands_6__7, CALCULATOR_L1FirstOperands_6__6, 
         CALCULATOR_L1FirstOperands_6__5, CALCULATOR_L1FirstOperands_6__4, 
         CALCULATOR_L1FirstOperands_6__3, CALCULATOR_L1FirstOperands_6__2, 
         CALCULATOR_L1FirstOperands_6__1, CALCULATOR_L1FirstOperands_6__0, 
         CALCULATOR_L1FirstOperands_7__7, CALCULATOR_L1FirstOperands_7__6, 
         CALCULATOR_L1FirstOperands_7__5, CALCULATOR_L1FirstOperands_7__4, 
         CALCULATOR_L1FirstOperands_7__3, CALCULATOR_L1FirstOperands_7__2, 
         CALCULATOR_L1FirstOperands_7__1, CALCULATOR_L1FirstOperands_7__0, 
         CALCULATOR_L1FirstOperands_8__7, CALCULATOR_L1FirstOperands_8__6, 
         CALCULATOR_L1FirstOperands_8__5, CALCULATOR_L1FirstOperands_8__4, 
         CALCULATOR_L1FirstOperands_8__3, CALCULATOR_L1FirstOperands_8__2, 
         CALCULATOR_L1FirstOperands_8__1, CALCULATOR_L1FirstOperands_8__0, 
         CALCULATOR_L1FirstOperands_9__7, CALCULATOR_L1FirstOperands_9__6, 
         CALCULATOR_L1FirstOperands_9__5, CALCULATOR_L1FirstOperands_9__4, 
         CALCULATOR_L1FirstOperands_9__3, CALCULATOR_L1FirstOperands_9__2, 
         CALCULATOR_L1FirstOperands_9__1, CALCULATOR_L1FirstOperands_9__0, 
         CALCULATOR_L1FirstOperands_10__7, CALCULATOR_L1FirstOperands_10__6, 
         CALCULATOR_L1FirstOperands_10__5, CALCULATOR_L1FirstOperands_10__4, 
         CALCULATOR_L1FirstOperands_10__3, CALCULATOR_L1FirstOperands_10__2, 
         CALCULATOR_L1FirstOperands_10__1, CALCULATOR_L1FirstOperands_10__0, 
         CALCULATOR_L1FirstOperands_11__7, CALCULATOR_L1FirstOperands_11__6, 
         CALCULATOR_L1FirstOperands_11__5, CALCULATOR_L1FirstOperands_11__4, 
         CALCULATOR_L1FirstOperands_11__3, CALCULATOR_L1FirstOperands_11__2, 
         CALCULATOR_L1FirstOperands_11__1, CALCULATOR_L1FirstOperands_11__0, 
         CALCULATOR_L1SecondOperands_0__7, CALCULATOR_L1SecondOperands_0__6, 
         CALCULATOR_L1SecondOperands_0__5, CALCULATOR_L1SecondOperands_0__4, 
         CALCULATOR_L1SecondOperands_0__3, CALCULATOR_L1SecondOperands_0__2, 
         CALCULATOR_L1SecondOperands_0__1, CALCULATOR_L1SecondOperands_0__0, 
         CALCULATOR_L1SecondOperands_1__7, CALCULATOR_L1SecondOperands_1__6, 
         CALCULATOR_L1SecondOperands_1__5, CALCULATOR_L1SecondOperands_1__4, 
         CALCULATOR_L1SecondOperands_1__3, CALCULATOR_L1SecondOperands_1__2, 
         CALCULATOR_L1SecondOperands_1__1, CALCULATOR_L1SecondOperands_1__0, 
         CALCULATOR_L1SecondOperands_2__7, CALCULATOR_L1SecondOperands_2__6, 
         CALCULATOR_L1SecondOperands_2__5, CALCULATOR_L1SecondOperands_2__4, 
         CALCULATOR_L1SecondOperands_2__3, CALCULATOR_L1SecondOperands_2__2, 
         CALCULATOR_L1SecondOperands_2__1, CALCULATOR_L1SecondOperands_2__0, 
         CALCULATOR_L1SecondOperands_3__7, CALCULATOR_L1SecondOperands_3__6, 
         CALCULATOR_L1SecondOperands_3__5, CALCULATOR_L1SecondOperands_3__4, 
         CALCULATOR_L1SecondOperands_3__3, CALCULATOR_L1SecondOperands_3__2, 
         CALCULATOR_L1SecondOperands_3__1, CALCULATOR_L1SecondOperands_3__0, 
         CALCULATOR_L1SecondOperands_4__7, CALCULATOR_L1SecondOperands_4__6, 
         CALCULATOR_L1SecondOperands_4__5, CALCULATOR_L1SecondOperands_4__4, 
         CALCULATOR_L1SecondOperands_4__3, CALCULATOR_L1SecondOperands_4__2, 
         CALCULATOR_L1SecondOperands_4__1, CALCULATOR_L1SecondOperands_4__0, 
         CALCULATOR_L1SecondOperands_5__7, CALCULATOR_L1SecondOperands_5__6, 
         CALCULATOR_L1SecondOperands_5__5, CALCULATOR_L1SecondOperands_5__4, 
         CALCULATOR_L1SecondOperands_5__3, CALCULATOR_L1SecondOperands_5__2, 
         CALCULATOR_L1SecondOperands_5__1, CALCULATOR_L1SecondOperands_5__0, 
         CALCULATOR_L1SecondOperands_6__7, CALCULATOR_L1SecondOperands_6__6, 
         CALCULATOR_L1SecondOperands_6__5, CALCULATOR_L1SecondOperands_6__4, 
         CALCULATOR_L1SecondOperands_6__3, CALCULATOR_L1SecondOperands_6__2, 
         CALCULATOR_L1SecondOperands_6__1, CALCULATOR_L1SecondOperands_6__0, 
         CALCULATOR_L1SecondOperands_7__7, CALCULATOR_L1SecondOperands_7__6, 
         CALCULATOR_L1SecondOperands_7__5, CALCULATOR_L1SecondOperands_7__4, 
         CALCULATOR_L1SecondOperands_7__3, CALCULATOR_L1SecondOperands_7__2, 
         CALCULATOR_L1SecondOperands_7__1, CALCULATOR_L1SecondOperands_7__0, 
         CALCULATOR_L1SecondOperands_8__7, CALCULATOR_L1SecondOperands_8__6, 
         CALCULATOR_L1SecondOperands_8__5, CALCULATOR_L1SecondOperands_8__4, 
         CALCULATOR_L1SecondOperands_8__3, CALCULATOR_L1SecondOperands_8__2, 
         CALCULATOR_L1SecondOperands_8__1, CALCULATOR_L1SecondOperands_8__0, 
         CALCULATOR_L1SecondOperands_9__7, CALCULATOR_L1SecondOperands_9__6, 
         CALCULATOR_L1SecondOperands_9__5, CALCULATOR_L1SecondOperands_9__4, 
         CALCULATOR_L1SecondOperands_9__3, CALCULATOR_L1SecondOperands_9__2, 
         CALCULATOR_L1SecondOperands_9__1, CALCULATOR_L1SecondOperands_9__0, 
         CALCULATOR_L1SecondOperands_10__7, CALCULATOR_L1SecondOperands_10__6, 
         CALCULATOR_L1SecondOperands_10__5, CALCULATOR_L1SecondOperands_10__4, 
         CALCULATOR_L1SecondOperands_10__3, CALCULATOR_L1SecondOperands_10__2, 
         CALCULATOR_L1SecondOperands_10__1, CALCULATOR_L1SecondOperands_10__0, 
         CALCULATOR_L1SecondOperands_11__7, CALCULATOR_L1SecondOperands_11__6, 
         CALCULATOR_L1SecondOperands_11__5, CALCULATOR_L1SecondOperands_11__4, 
         CALCULATOR_L1SecondOperands_11__3, CALCULATOR_L1SecondOperands_11__2, 
         CALCULATOR_L1SecondOperands_11__1, CALCULATOR_L1SecondOperands_11__0, 
         CALCULATOR_L1Results_0__7, CALCULATOR_L1Results_0__6, 
         CALCULATOR_L1Results_0__5, CALCULATOR_L1Results_0__4, 
         CALCULATOR_L1Results_0__3, CALCULATOR_L1Results_0__2, 
         CALCULATOR_L1Results_0__1, CALCULATOR_L1Results_0__0, 
         CALCULATOR_L1Results_1__7, CALCULATOR_L1Results_1__6, 
         CALCULATOR_L1Results_1__5, CALCULATOR_L1Results_1__4, 
         CALCULATOR_L1Results_1__3, CALCULATOR_L1Results_1__2, 
         CALCULATOR_L1Results_1__1, CALCULATOR_L1Results_1__0, 
         CALCULATOR_L1Results_2__7, CALCULATOR_L1Results_2__6, 
         CALCULATOR_L1Results_2__5, CALCULATOR_L1Results_2__4, 
         CALCULATOR_L1Results_2__3, CALCULATOR_L1Results_2__2, 
         CALCULATOR_L1Results_2__1, CALCULATOR_L1Results_2__0, 
         CALCULATOR_L1Results_3__7, CALCULATOR_L1Results_3__6, 
         CALCULATOR_L1Results_3__5, CALCULATOR_L1Results_3__4, 
         CALCULATOR_L1Results_3__3, CALCULATOR_L1Results_3__2, 
         CALCULATOR_L1Results_3__1, CALCULATOR_L1Results_3__0, 
         CALCULATOR_L1Results_4__7, CALCULATOR_L1Results_4__6, 
         CALCULATOR_L1Results_4__5, CALCULATOR_L1Results_4__4, 
         CALCULATOR_L1Results_4__3, CALCULATOR_L1Results_4__2, 
         CALCULATOR_L1Results_4__1, CALCULATOR_L1Results_4__0, 
         CALCULATOR_L1Results_5__7, CALCULATOR_L1Results_5__6, 
         CALCULATOR_L1Results_5__5, CALCULATOR_L1Results_5__4, 
         CALCULATOR_L1Results_5__3, CALCULATOR_L1Results_5__2, 
         CALCULATOR_L1Results_5__1, CALCULATOR_L1Results_5__0, 
         CALCULATOR_L1Results_6__7, CALCULATOR_L1Results_6__6, 
         CALCULATOR_L1Results_6__5, CALCULATOR_L1Results_6__4, 
         CALCULATOR_L1Results_6__3, CALCULATOR_L1Results_6__2, 
         CALCULATOR_L1Results_6__1, CALCULATOR_L1Results_6__0, 
         CALCULATOR_L1Results_7__7, CALCULATOR_L1Results_7__6, 
         CALCULATOR_L1Results_7__5, CALCULATOR_L1Results_7__4, 
         CALCULATOR_L1Results_7__3, CALCULATOR_L1Results_7__2, 
         CALCULATOR_L1Results_7__1, CALCULATOR_L1Results_7__0, 
         CALCULATOR_L1Results_8__7, CALCULATOR_L1Results_8__6, 
         CALCULATOR_L1Results_8__5, CALCULATOR_L1Results_8__4, 
         CALCULATOR_L1Results_8__3, CALCULATOR_L1Results_8__2, 
         CALCULATOR_L1Results_8__1, CALCULATOR_L1Results_8__0, 
         CALCULATOR_L1Results_9__7, CALCULATOR_L1Results_9__6, 
         CALCULATOR_L1Results_9__5, CALCULATOR_L1Results_9__4, 
         CALCULATOR_L1Results_9__3, CALCULATOR_L1Results_9__2, 
         CALCULATOR_L1Results_9__1, CALCULATOR_L1Results_9__0, 
         CALCULATOR_L1Results_10__7, CALCULATOR_L1Results_10__6, 
         CALCULATOR_L1Results_10__5, CALCULATOR_L1Results_10__4, 
         CALCULATOR_L1Results_10__3, CALCULATOR_L1Results_10__2, 
         CALCULATOR_L1Results_10__1, CALCULATOR_L1Results_10__0, 
         CALCULATOR_L1Results_11__7, CALCULATOR_L1Results_11__6, 
         CALCULATOR_L1Results_11__5, CALCULATOR_L1Results_11__4, 
         CALCULATOR_L1Results_11__3, CALCULATOR_L1Results_11__2, 
         CALCULATOR_L1Results_11__1, CALCULATOR_L1Results_11__0, 
         CALCULATOR_L2Results_0__7, CALCULATOR_L2Results_0__6, 
         CALCULATOR_L2Results_0__5, CALCULATOR_L2Results_0__4, 
         CALCULATOR_L2Results_0__3, CALCULATOR_L2Results_0__2, 
         CALCULATOR_L2Results_0__1, CALCULATOR_L2Results_0__0, 
         CALCULATOR_L2Results_1__7, CALCULATOR_L2Results_1__6, 
         CALCULATOR_L2Results_1__5, CALCULATOR_L2Results_1__4, 
         CALCULATOR_L2Results_1__3, CALCULATOR_L2Results_1__2, 
         CALCULATOR_L2Results_1__1, CALCULATOR_L2Results_1__0, 
         CALCULATOR_L2Results_2__7, CALCULATOR_L2Results_2__6, 
         CALCULATOR_L2Results_2__5, CALCULATOR_L2Results_2__4, 
         CALCULATOR_L2Results_2__3, CALCULATOR_L2Results_2__2, 
         CALCULATOR_L2Results_2__1, CALCULATOR_L2Results_2__0, 
         CALCULATOR_L2Results_3__7, CALCULATOR_L2Results_3__6, 
         CALCULATOR_L2Results_3__5, CALCULATOR_L2Results_3__4, 
         CALCULATOR_L2Results_3__3, CALCULATOR_L2Results_3__2, 
         CALCULATOR_L2Results_3__1, CALCULATOR_L2Results_3__0, 
         CALCULATOR_L2Results_4__7, CALCULATOR_L2Results_4__6, 
         CALCULATOR_L2Results_4__5, CALCULATOR_L2Results_4__4, 
         CALCULATOR_L2Results_4__3, CALCULATOR_L2Results_4__2, 
         CALCULATOR_L2Results_4__1, CALCULATOR_L2Results_4__0, 
         CALCULATOR_L2Results_5__7, CALCULATOR_L2Results_5__6, 
         CALCULATOR_L2Results_5__5, CALCULATOR_L2Results_5__4, 
         CALCULATOR_L2Results_5__3, CALCULATOR_L2Results_5__2, 
         CALCULATOR_L2Results_5__1, CALCULATOR_L2Results_5__0, 
         CALCULATOR_L3Results_0__7, CALCULATOR_L3Results_0__6, 
         CALCULATOR_L3Results_0__5, CALCULATOR_L3Results_0__4, 
         CALCULATOR_L3Results_0__3, CALCULATOR_L3Results_0__2, 
         CALCULATOR_L3Results_0__1, CALCULATOR_L3Results_0__0, 
         CALCULATOR_L3Results_1__7, CALCULATOR_L3Results_1__6, 
         CALCULATOR_L3Results_1__5, CALCULATOR_L3Results_1__4, 
         CALCULATOR_L3Results_1__3, CALCULATOR_L3Results_1__2, 
         CALCULATOR_L3Results_1__1, CALCULATOR_L3Results_1__0, 
         CALCULATOR_L3Results_2__7, CALCULATOR_L3Results_2__6, 
         CALCULATOR_L3Results_2__5, CALCULATOR_L3Results_2__4, 
         CALCULATOR_L3Results_2__3, CALCULATOR_L3Results_2__2, 
         CALCULATOR_L3Results_2__1, CALCULATOR_L3Results_2__0, 
         CALCULATOR_L4Results_0__7, CALCULATOR_L4Results_0__6, 
         CALCULATOR_L4Results_0__5, CALCULATOR_L4Results_0__4, 
         CALCULATOR_L4Results_0__3, CALCULATOR_L4Results_0__2, 
         CALCULATOR_L4Results_0__1, CALCULATOR_L4Results_0__0, 
         CALCULATOR_L5FirstOperands_1__7, CALCULATOR_L5FirstOperands_1__6, 
         CALCULATOR_L5FirstOperands_1__5, CALCULATOR_L5FirstOperands_1__4, 
         CALCULATOR_L5FirstOperands_1__3, CALCULATOR_L5FirstOperands_1__2, 
         CALCULATOR_L5FirstOperands_1__1, CALCULATOR_L5FirstOperands_1__0, 
         CALCULATOR_L5SecondOperands_1__7, CALCULATOR_L5SecondOperands_1__6, 
         CALCULATOR_L5SecondOperands_1__5, CALCULATOR_L5SecondOperands_1__4, 
         CALCULATOR_L5SecondOperands_1__3, CALCULATOR_L5SecondOperands_1__2, 
         CALCULATOR_L5SecondOperands_1__1, CALCULATOR_L5SecondOperands_1__0, 
         CALCULATOR_L5Results_1__7, CALCULATOR_L5Results_1__6, 
         CALCULATOR_L5Results_1__5, CALCULATOR_L5Results_1__4, 
         CALCULATOR_L5Results_1__3, CALCULATOR_L5Results_1__2, 
         CALCULATOR_L5Results_1__1, CALCULATOR_L5Results_1__0, CALCULATOR_nx22, 
         CALCULATOR_nx78, CALCULATOR_nx990, CALCULATOR_nx993, CALCULATOR_nx995, 
         CALCULATOR_nx1001, CALCULATOR_nx1003, CALCULATOR_nx1007, 
         CALCULATOR_nx1009, CALCULATOR_nx1012, CALCULATOR_nx1014, 
         CALCULATOR_nx1043, CALCULATOR_CalculatingBooth_dup_1146, 
         CALCULATOR_CalculatingBooth_dup_1181, 
         CALCULATOR_CalculatingBooth_dup_1224, 
         CALCULATOR_CalculatingBooth_dup_1315, CALCULATOR_Start_dup_1144, 
         CALCULATOR_Start_dup_1149, CALCULATOR_Start_dup_1154, 
         CALCULATOR_Start_dup_1159, CALCULATOR_Start_dup_1164, 
         CALCULATOR_Start_dup_1169, CALCULATOR_Start_dup_1174, 
         CALCULATOR_Start_dup_1179, CALCULATOR_Start_dup_1184, 
         CALCULATOR_Start_dup_1189, CALCULATOR_Start_dup_1194, 
         CALCULATOR_Start_dup_1199, CALCULATOR_Start_dup_1204, 
         CALCULATOR_Start_dup_1209, CALCULATOR_Start_dup_1222, 
         CALCULATOR_Start_dup_1235, CALCULATOR_Start_dup_1248, 
         CALCULATOR_Start_dup_1261, CALCULATOR_Start_dup_1274, 
         CALCULATOR_Start_dup_1287, CALCULATOR_Start_dup_1300, 
         CALCULATOR_Start_dup_1313, CALCULATOR_Start_dup_1326, 
         CALCULATOR_Start_dup_1339, CALCULATOR_Start_dup_1352, CALCULATOR_nx1111, 
         CALCULATOR_ACCELERATOR_COUNTER_nx6, CALCULATOR_ACCELERATOR_COUNTER_nx12, 
         CALCULATOR_ACCELERATOR_COUNTER_nx18, 
         CALCULATOR_ACCELERATOR_COUNTER_nx81, 
         CALCULATOR_ACCELERATOR_COUNTER_nx91, 
         CALCULATOR_ACCELERATOR_COUNTER_nx101, 
         CALCULATOR_ACCELERATOR_COUNTER_nx111, 
         CALCULATOR_ACCELERATOR_COUNTER_nx133, 
         CALCULATOR_ACCELERATOR_COUNTER_nx139, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_AddPToBoothOperand, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothOperand_16, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothOperand_15, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothOperand_14, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothOperand_13, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothOperand_12, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothOperand_11, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothOperand_10, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothOperand_9, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothOperand_8, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothOperand_7, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothOperand_6, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothOperand_5, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothOperand_4, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothOperand_3, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothOperand_2, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothOperand_1, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothOperand_0, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_16, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_15, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_14, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_13, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_12, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_11, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_10, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_9, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_8, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_7, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_6, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_5, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_4, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_3, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_2, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_1, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_16, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_15, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_14, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_13, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_12, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_11, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_10, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_9, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_8, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_7, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_6, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_5, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_4, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_3, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_2, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_1, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_0, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx0, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx6, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx12, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx18, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx24, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx30, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx40, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx44, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx48, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx52, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx56, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx62, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx154, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx316, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx336, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx356, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx376, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx396, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx416, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx436, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx454, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx456, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx379, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx381, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx383, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx387, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx389, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx391, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx395, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx399, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx401, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx403, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx405, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx409, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx411, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx413, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx415, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx419, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx421, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx423, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx425, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx429, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx431, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx433, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx435, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx439, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx441, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx443, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx445, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx449, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx451, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx453, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx455, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx461, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx463, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx467, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx469, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx471, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx475, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx477, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx479, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx483, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx485, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx487, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx491, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx493, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx495, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx499, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx501, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx503, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx507, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx509, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx511, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx515, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx517, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx529, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx531, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx534, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx537, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx540, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx544, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx547, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx551, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx554, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx558, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx561, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx565, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx568, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_WindowCellShiftedLeft_16, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_16, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_15, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_14, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_13, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_12, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_11, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_10, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_16, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_15, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_14, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_13, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_12, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_11, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_10, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_9, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_8, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_7, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_6, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_5, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_4, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_3, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_2, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_1, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_0, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_16, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_15, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_14, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_13, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_12, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_11, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_10, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_9, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_8, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_7, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_6, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_5, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_4, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_3, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_2, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_1, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_0, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_16, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_15, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_14, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_13, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_12, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_11, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_10, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_9, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_8, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_7, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_6, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_5, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_4, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_3, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_2, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_1, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_0, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx4, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx8, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx12, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx16, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx20, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx24, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx80, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx328, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx384, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx564, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642, 
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_AddPToBoothOperand, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothOperand_16, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothOperand_15, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothOperand_14, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothOperand_13, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothOperand_12, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothOperand_11, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothOperand_10, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothOperand_9, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothOperand_8, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothOperand_7, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothOperand_6, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothOperand_5, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothOperand_4, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothOperand_3, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothOperand_2, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothOperand_1, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothOperand_0, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_16, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_15, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_14, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_13, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_12, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_11, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_10, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_9, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_8, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_7, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_6, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_5, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_4, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_3, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_2, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_1, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_16, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_15, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_14, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_13, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_12, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_11, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_10, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_9, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_8, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_7, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_6, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_5, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_4, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_3, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_2, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_1, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_0, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx0, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx6, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx12, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx18, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx24, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx30, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx40, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx44, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx48, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx52, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx56, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx62, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx154, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx316, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx336, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx356, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx376, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx396, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx416, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx436, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx454, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx456, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx379, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx381, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx383, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx387, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx389, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx391, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx395, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx399, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx401, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx403, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx405, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx409, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx411, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx413, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx415, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx419, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx421, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx423, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx425, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx429, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx431, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx433, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx435, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx439, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx441, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx443, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx445, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx449, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx451, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx453, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx455, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx461, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx463, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx467, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx469, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx471, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx475, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx477, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx479, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx483, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx485, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx487, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx491, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx493, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx495, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx499, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx501, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx503, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx507, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx509, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx511, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx515, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx517, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx529, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx531, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx534, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx537, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx540, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx544, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx547, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx551, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx554, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx558, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx561, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx565, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx568, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_WindowCellShiftedLeft_16, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_16, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_15, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_14, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_13, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_12, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_11, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_10, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_16, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_15, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_14, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_13, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_12, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_11, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_10, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_9, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_8, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_7, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_6, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_5, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_4, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_3, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_2, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_1, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_0, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_16, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_15, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_14, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_13, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_12, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_11, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_10, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_9, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_8, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_7, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_6, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_5, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_4, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_3, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_2, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_1, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_0, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_16, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_15, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_14, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_13, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_12, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_11, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_10, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_9, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_8, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_7, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_6, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_5, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_4, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_3, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_2, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_1, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_0, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx4, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx8, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx12, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx16, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx20, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx24, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx80, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx328, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx384, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642, 
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_AddPToBoothOperand, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothOperand_16, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothOperand_15, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothOperand_14, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothOperand_13, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothOperand_12, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothOperand_11, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothOperand_10, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothOperand_9, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothOperand_8, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothOperand_7, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothOperand_6, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothOperand_5, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothOperand_4, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothOperand_3, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothOperand_2, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothOperand_1, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothOperand_0, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_16, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_15, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_14, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_13, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_12, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_11, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_10, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_9, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_8, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_7, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_6, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_5, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_4, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_3, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_2, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_1, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_16, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_15, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_14, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_13, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_12, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_11, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_10, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_9, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_8, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_7, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_6, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_5, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_4, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_3, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_2, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_1, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_0, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx0, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx6, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx12, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx18, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx24, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx30, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx40, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx44, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx48, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx52, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx56, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx62, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx154, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx316, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx336, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx356, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx376, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx396, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx416, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx436, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx454, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx456, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx379, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx381, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx383, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx387, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx389, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx391, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx395, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx399, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx401, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx403, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx405, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx409, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx411, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx413, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx415, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx419, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx421, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx423, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx425, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx429, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx431, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx433, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx435, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx439, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx441, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx443, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx445, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx449, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx451, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx453, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx455, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx461, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx463, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx467, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx469, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx471, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx475, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx477, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx479, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx483, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx485, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx487, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx491, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx493, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx495, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx499, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx501, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx503, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx507, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx509, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx511, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx515, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx517, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx529, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx531, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx534, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx537, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx540, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx544, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx547, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx551, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx554, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx558, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx561, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx565, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx568, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_WindowCellShiftedLeft_16, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_16, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_15, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_14, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_13, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_12, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_11, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_10, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_16, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_15, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_14, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_13, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_12, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_11, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_10, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_9, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_8, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_7, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_6, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_5, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_4, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_3, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_2, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_1, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_0, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_16, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_15, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_14, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_13, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_12, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_11, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_10, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_9, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_8, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_7, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_6, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_5, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_4, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_3, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_2, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_1, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_0, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_16, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_15, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_14, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_13, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_12, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_11, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_10, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_9, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_8, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_7, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_6, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_5, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_4, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_3, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_2, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_1, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_0, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx4, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx8, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx12, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx16, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx20, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx24, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx80, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx328, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx384, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642, 
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_AddPToBoothOperand, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothOperand_16, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothOperand_15, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothOperand_14, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothOperand_13, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothOperand_12, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothOperand_11, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothOperand_10, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothOperand_9, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothOperand_8, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothOperand_7, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothOperand_6, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothOperand_5, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothOperand_4, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothOperand_3, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothOperand_2, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothOperand_1, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothOperand_0, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_16, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_15, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_14, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_13, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_12, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_11, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_10, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_9, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_8, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_7, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_6, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_5, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_4, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_3, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_2, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_1, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_16, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_15, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_14, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_13, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_12, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_11, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_10, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_9, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_8, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_7, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_6, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_5, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_4, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_3, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_2, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_1, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_0, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx0, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx6, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx12, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx18, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx24, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx30, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx40, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx44, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx48, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx52, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx56, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx62, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx154, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx316, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx336, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx356, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx376, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx396, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx416, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx436, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx454, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx456, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx379, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx381, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx383, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx387, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx389, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx391, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx395, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx399, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx401, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx403, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx405, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx409, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx411, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx413, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx415, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx419, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx421, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx423, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx425, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx429, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx431, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx433, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx435, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx439, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx441, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx443, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx445, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx449, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx451, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx453, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx455, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx461, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx463, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx467, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx469, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx471, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx475, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx477, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx479, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx483, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx485, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx487, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx491, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx493, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx495, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx499, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx501, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx503, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx507, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx509, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx511, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx515, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx517, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx529, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx531, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx534, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx537, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx540, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx544, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx547, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx551, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx554, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx558, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx561, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx565, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx568, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_WindowCellShiftedLeft_16, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_16, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_15, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_14, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_13, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_12, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_11, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_10, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_16, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_15, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_14, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_13, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_12, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_11, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_10, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_9, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_8, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_7, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_6, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_5, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_4, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_3, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_2, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_1, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_0, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_16, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_15, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_14, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_13, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_12, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_11, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_10, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_9, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_8, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_7, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_6, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_5, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_4, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_3, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_2, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_1, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_0, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_16, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_15, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_14, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_13, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_12, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_11, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_10, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_9, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_8, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_7, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_6, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_5, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_4, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_3, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_2, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_1, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_0, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx4, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx8, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx12, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx16, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx20, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx24, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx80, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx328, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx384, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642, 
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_AddPToBoothOperand, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothOperand_16, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothOperand_15, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothOperand_14, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothOperand_13, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothOperand_12, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothOperand_11, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothOperand_10, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothOperand_9, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothOperand_8, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothOperand_7, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothOperand_6, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothOperand_5, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothOperand_4, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothOperand_3, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothOperand_2, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothOperand_1, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothOperand_0, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_16, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_15, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_14, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_13, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_12, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_11, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_10, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_9, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_8, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_7, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_6, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_5, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_4, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_3, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_2, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_1, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_16, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_15, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_14, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_13, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_12, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_11, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_10, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_9, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_8, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_7, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_6, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_5, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_4, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_3, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_2, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_1, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_0, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx0, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx6, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx12, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx18, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx24, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx30, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx40, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx44, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx48, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx52, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx56, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx62, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx154, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx316, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx336, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx356, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx376, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx396, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx416, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx436, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx454, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx456, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx379, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx381, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx383, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx387, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx389, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx391, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx395, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx399, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx401, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx403, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx405, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx409, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx411, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx413, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx415, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx419, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx421, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx423, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx425, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx429, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx431, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx433, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx435, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx439, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx441, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx443, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx445, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx449, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx451, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx453, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx455, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx461, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx463, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx467, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx469, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx471, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx475, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx477, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx479, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx483, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx485, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx487, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx491, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx493, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx495, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx499, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx501, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx503, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx507, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx509, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx511, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx515, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx517, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx529, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx531, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx534, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx537, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx540, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx544, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx547, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx551, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx554, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx558, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx561, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx565, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx568, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_WindowCellShiftedLeft_16, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_16, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_15, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_14, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_13, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_12, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_11, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_10, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_16, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_15, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_14, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_13, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_12, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_11, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_10, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_9, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_8, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_7, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_6, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_5, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_4, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_3, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_2, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_1, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_0, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_16, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_15, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_14, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_13, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_12, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_11, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_10, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_9, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_8, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_7, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_6, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_5, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_4, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_3, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_2, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_1, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_0, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_16, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_15, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_14, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_13, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_12, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_11, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_10, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_9, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_8, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_7, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_6, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_5, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_4, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_3, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_2, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_1, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_0, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx4, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx8, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx12, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx16, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx20, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx24, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx80, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx328, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx384, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642, 
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_AddPToBoothOperand, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothOperand_16, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothOperand_15, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothOperand_14, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothOperand_13, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothOperand_12, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothOperand_11, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothOperand_10, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothOperand_9, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothOperand_8, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothOperand_7, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothOperand_6, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothOperand_5, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothOperand_4, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothOperand_3, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothOperand_2, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothOperand_1, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothOperand_0, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_16, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_15, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_14, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_13, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_12, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_11, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_10, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_9, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_8, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_7, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_6, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_5, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_4, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_3, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_2, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_1, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_16, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_15, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_14, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_13, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_12, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_11, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_10, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_9, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_8, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_7, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_6, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_5, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_4, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_3, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_2, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_1, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_0, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx0, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx6, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx12, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx18, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx24, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx30, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx40, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx44, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx48, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx52, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx56, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx62, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx154, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx316, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx336, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx356, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx376, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx396, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx416, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx436, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx454, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx456, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx379, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx381, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx383, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx387, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx389, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx391, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx395, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx399, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx401, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx403, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx405, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx409, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx411, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx413, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx415, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx419, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx421, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx423, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx425, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx429, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx431, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx433, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx435, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx439, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx441, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx443, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx445, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx449, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx451, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx453, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx455, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx461, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx463, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx467, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx469, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx471, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx475, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx477, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx479, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx483, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx485, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx487, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx491, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx493, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx495, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx499, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx501, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx503, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx507, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx509, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx511, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx515, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx517, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx529, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx531, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx534, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx537, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx540, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx544, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx547, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx551, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx554, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx558, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx561, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx565, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx568, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_WindowCellShiftedLeft_16, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_16, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_15, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_14, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_13, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_12, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_11, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_10, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_16, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_15, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_14, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_13, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_12, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_11, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_10, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_9, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_8, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_7, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_6, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_5, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_4, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_3, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_2, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_1, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_0, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_16, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_15, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_14, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_13, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_12, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_11, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_10, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_9, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_8, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_7, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_6, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_5, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_4, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_3, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_2, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_1, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_0, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_16, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_15, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_14, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_13, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_12, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_11, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_10, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_9, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_8, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_7, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_6, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_5, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_4, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_3, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_2, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_1, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_0, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx4, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx8, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx12, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx16, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx20, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx24, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx80, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx328, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx384, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642, 
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_AddPToBoothOperand, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothOperand_16, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothOperand_15, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothOperand_14, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothOperand_13, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothOperand_12, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothOperand_11, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothOperand_10, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothOperand_9, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothOperand_8, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothOperand_7, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothOperand_6, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothOperand_5, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothOperand_4, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothOperand_3, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothOperand_2, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothOperand_1, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothOperand_0, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_16, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_15, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_14, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_13, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_12, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_11, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_10, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_9, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_8, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_7, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_6, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_5, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_4, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_3, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_2, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_1, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_16, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_15, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_14, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_13, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_12, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_11, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_10, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_9, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_8, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_7, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_6, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_5, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_4, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_3, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_2, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_1, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_0, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx0, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx6, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx12, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx18, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx24, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx30, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx40, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx44, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx48, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx52, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx56, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx62, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx154, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx316, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx336, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx356, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx376, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx396, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx416, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx436, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx454, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx456, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx379, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx381, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx383, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx387, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx389, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx391, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx395, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx399, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx401, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx403, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx405, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx409, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx411, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx413, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx415, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx419, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx421, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx423, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx425, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx429, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx431, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx433, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx435, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx439, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx441, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx443, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx445, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx449, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx451, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx453, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx455, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx461, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx463, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx467, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx469, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx471, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx475, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx477, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx479, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx483, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx485, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx487, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx491, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx493, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx495, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx499, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx501, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx503, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx507, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx509, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx511, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx515, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx517, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx529, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx531, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx534, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx537, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx540, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx544, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx547, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx551, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx554, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx558, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx561, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx565, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx568, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_WindowCellShiftedLeft_16, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_16, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_15, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_14, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_13, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_12, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_11, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_10, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_16, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_15, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_14, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_13, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_12, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_11, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_10, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_9, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_8, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_7, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_6, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_5, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_4, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_3, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_2, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_1, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_0, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_16, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_15, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_14, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_13, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_12, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_11, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_10, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_9, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_8, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_7, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_6, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_5, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_4, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_3, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_2, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_1, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_0, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_16, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_15, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_14, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_13, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_12, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_11, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_10, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_9, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_8, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_7, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_6, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_5, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_4, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_3, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_2, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_1, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_0, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx4, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx8, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx12, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx16, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx20, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx24, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx80, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx328, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx384, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642, 
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_AddPToBoothOperand, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothOperand_16, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothOperand_15, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothOperand_14, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothOperand_13, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothOperand_12, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothOperand_11, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothOperand_10, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothOperand_9, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothOperand_8, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothOperand_7, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothOperand_6, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothOperand_5, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothOperand_4, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothOperand_3, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothOperand_2, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothOperand_1, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothOperand_0, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_16, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_15, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_14, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_13, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_12, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_11, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_10, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_9, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_8, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_7, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_6, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_5, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_4, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_3, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_2, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_1, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_16, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_15, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_14, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_13, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_12, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_11, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_10, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_9, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_8, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_7, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_6, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_5, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_4, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_3, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_2, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_1, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_0, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx0, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx6, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx12, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx18, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx24, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx30, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx40, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx44, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx48, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx52, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx56, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx62, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx154, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx316, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx336, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx356, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx376, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx396, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx416, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx436, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx454, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx456, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx379, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx381, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx383, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx387, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx389, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx391, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx395, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx399, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx401, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx403, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx405, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx409, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx411, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx413, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx415, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx419, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx421, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx423, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx425, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx429, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx431, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx433, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx435, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx439, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx441, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx443, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx445, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx449, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx451, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx453, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx455, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx461, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx463, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx467, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx469, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx471, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx475, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx477, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx479, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx483, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx485, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx487, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx491, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx493, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx495, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx499, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx501, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx503, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx507, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx509, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx511, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx515, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx517, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx529, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx531, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx534, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx537, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx540, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx544, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx547, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx551, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx554, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx558, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx561, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx565, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx568, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_WindowCellShiftedLeft_16, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_16, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_15, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_14, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_13, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_12, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_11, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_10, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_16, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_15, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_14, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_13, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_12, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_11, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_10, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_9, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_8, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_7, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_6, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_5, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_4, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_3, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_2, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_1, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_0, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_16, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_15, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_14, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_13, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_12, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_11, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_10, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_9, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_8, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_7, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_6, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_5, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_4, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_3, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_2, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_1, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_0, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_16, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_15, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_14, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_13, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_12, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_11, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_10, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_9, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_8, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_7, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_6, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_5, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_4, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_3, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_2, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_1, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_0, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx4, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx8, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx12, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx16, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx20, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx24, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx80, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx328, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx384, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642, 
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_AddPToBoothOperand, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothOperand_16, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothOperand_15, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothOperand_14, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothOperand_13, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothOperand_12, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothOperand_11, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothOperand_10, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothOperand_9, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothOperand_8, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothOperand_7, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothOperand_6, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothOperand_5, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothOperand_4, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothOperand_3, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothOperand_2, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothOperand_1, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothOperand_0, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_16, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_15, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_14, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_13, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_12, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_11, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_10, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_9, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_8, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_7, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_6, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_5, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_4, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_3, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_2, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_1, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_16, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_15, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_14, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_13, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_12, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_11, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_10, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_9, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_8, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_7, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_6, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_5, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_4, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_3, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_2, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_1, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_0, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx0, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx6, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx12, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx18, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx24, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx30, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx40, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx44, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx48, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx52, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx56, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx62, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx154, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx316, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx336, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx356, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx376, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx396, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx416, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx436, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx454, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx456, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx379, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx381, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx383, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx387, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx389, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx391, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx395, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx399, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx401, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx403, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx405, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx409, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx411, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx413, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx415, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx419, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx421, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx423, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx425, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx429, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx431, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx433, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx435, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx439, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx441, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx443, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx445, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx449, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx451, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx453, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx455, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx461, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx463, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx467, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx469, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx471, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx475, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx477, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx479, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx483, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx485, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx487, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx491, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx493, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx495, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx499, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx501, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx503, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx507, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx509, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx511, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx515, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx517, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx529, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx531, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx534, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx537, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx540, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx544, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx547, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx551, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx554, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx558, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx561, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx565, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx568, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_WindowCellShiftedLeft_16, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_16, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_15, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_14, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_13, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_12, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_11, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_10, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_16, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_15, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_14, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_13, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_12, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_11, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_10, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_9, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_8, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_7, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_6, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_5, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_4, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_3, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_2, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_1, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_0, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_16, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_15, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_14, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_13, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_12, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_11, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_10, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_9, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_8, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_7, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_6, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_5, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_4, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_3, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_2, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_1, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_0, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_16, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_15, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_14, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_13, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_12, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_11, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_10, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_9, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_8, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_7, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_6, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_5, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_4, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_3, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_2, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_1, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_0, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx4, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx8, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx12, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx16, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx20, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx24, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx80, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx328, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx384, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642, 
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_AddPToBoothOperand, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothOperand_16, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothOperand_15, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothOperand_14, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothOperand_13, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothOperand_12, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothOperand_11, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothOperand_10, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothOperand_9, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothOperand_8, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothOperand_7, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothOperand_6, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothOperand_5, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothOperand_4, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothOperand_3, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothOperand_2, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothOperand_1, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothOperand_0, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_16, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_15, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_14, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_13, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_12, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_11, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_10, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_9, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_8, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_7, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_6, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_5, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_4, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_3, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_2, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_1, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_16, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_15, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_14, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_13, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_12, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_11, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_10, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_9, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_8, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_7, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_6, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_5, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_4, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_3, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_2, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_1, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_0, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx0, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx6, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx12, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx18, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx24, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx30, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx40, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx44, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx48, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx52, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx56, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx62, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx154, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx316, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx336, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx356, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx376, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx396, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx416, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx436, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx454, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx456, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx379, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx381, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx383, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx387, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx389, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx391, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx395, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx399, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx401, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx403, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx405, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx409, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx411, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx413, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx415, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx419, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx421, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx423, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx425, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx429, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx431, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx433, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx435, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx439, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx441, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx443, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx445, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx449, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx451, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx453, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx455, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx461, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx463, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx467, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx469, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx471, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx475, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx477, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx479, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx483, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx485, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx487, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx491, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx493, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx495, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx499, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx501, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx503, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx507, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx509, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx511, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx515, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx517, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx529, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx531, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx534, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx537, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx540, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx544, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx547, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx551, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx554, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx558, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx561, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx565, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx568, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_WindowCellShiftedLeft_16, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_16, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_15, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_14, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_13, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_12, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_11, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_10, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_16, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_15, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_14, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_13, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_12, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_11, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_10, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_9, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_8, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_7, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_6, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_5, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_4, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_3, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_2, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_1, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_0, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_16, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_15, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_14, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_13, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_12, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_11, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_10, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_9, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_8, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_7, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_6, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_5, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_4, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_3, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_2, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_1, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_0, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_16, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_15, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_14, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_13, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_12, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_11, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_10, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_9, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_8, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_7, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_6, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_5, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_4, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_3, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_2, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_1, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_0, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx4, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx8, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx12, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx16, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx20, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx24, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx80, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx328, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx384, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642, 
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_AddPToBoothOperand, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothOperand_16, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothOperand_15, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothOperand_14, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothOperand_13, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothOperand_12, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothOperand_11, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothOperand_10, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothOperand_9, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothOperand_8, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothOperand_7, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothOperand_6, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothOperand_5, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothOperand_4, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothOperand_3, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothOperand_2, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothOperand_1, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothOperand_0, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_16, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_15, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_14, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_13, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_12, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_11, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_10, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_9, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_8, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_7, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_6, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_5, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_4, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_3, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_2, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_1, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_16, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_15, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_14, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_13, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_12, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_11, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_10, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_9, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_8, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_7, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_6, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_5, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_4, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_3, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_2, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_1, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_0, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx0, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx6, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx12, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx18, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx24, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx30, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx40, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx44, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx48, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx52, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx56, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx62, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx154, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx316, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx336, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx356, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx376, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx396, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx416, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx436, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx454, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx456, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx379, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx381, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx383, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx387, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx389, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx391, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx395, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx399, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx401, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx403, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx405, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx409, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx411, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx413, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx415, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx419, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx421, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx423, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx425, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx429, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx431, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx433, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx435, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx439, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx441, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx443, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx445, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx449, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx451, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx453, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx455, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx461, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx463, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx467, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx469, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx471, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx475, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx477, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx479, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx483, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx485, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx487, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx491, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx493, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx495, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx499, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx501, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx503, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx507, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx509, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx511, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx515, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx517, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx529, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx531, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx534, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx537, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx540, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx544, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx547, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx551, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx554, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx558, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx561, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx565, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx568, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_WindowCellShiftedLeft_16, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_16, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_15, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_14, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_13, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_12, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_11, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_10, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_16, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_15, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_14, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_13, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_12, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_11, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_10, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_9, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_8, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_7, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_6, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_5, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_4, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_3, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_2, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_1, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_0, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_16, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_15, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_14, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_13, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_12, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_11, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_10, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_9, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_8, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_7, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_6, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_5, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_4, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_3, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_2, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_1, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_0, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_16, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_15, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_14, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_13, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_12, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_11, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_10, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_9, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_8, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_7, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_6, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_5, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_4, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_3, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_2, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_1, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_0, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx4, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx8, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx12, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx16, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx20, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx24, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx80, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx328, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx384, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642, 
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_AddPToBoothOperand, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothOperand_16, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothOperand_15, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothOperand_14, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothOperand_13, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothOperand_12, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothOperand_11, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothOperand_10, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothOperand_9, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothOperand_8, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothOperand_7, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothOperand_6, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothOperand_5, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothOperand_4, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothOperand_3, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothOperand_2, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothOperand_1, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothOperand_0, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_16, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_15, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_14, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_13, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_12, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_11, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_10, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_9, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_8, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_7, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_6, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_5, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_4, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_3, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_2, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_1, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_16, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_15, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_14, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_13, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_12, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_11, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_10, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_9, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_8, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_7, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_6, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_5, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_4, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_3, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_2, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_1, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_0, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx0, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx6, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx12, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx18, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx24, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx30, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx40, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx44, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx48, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx52, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx56, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx62, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx154, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx316, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx336, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx356, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx376, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx396, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx416, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx436, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx454, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx456, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx379, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx381, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx383, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx387, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx389, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx391, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx395, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx399, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx401, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx403, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx405, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx409, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx411, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx413, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx415, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx419, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx421, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx423, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx425, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx429, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx431, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx433, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx435, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx439, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx441, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx443, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx445, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx449, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx451, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx453, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx455, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx461, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx463, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx467, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx469, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx471, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx475, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx477, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx479, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx483, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx485, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx487, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx491, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx493, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx495, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx499, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx501, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx503, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx507, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx509, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx511, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx515, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx517, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx529, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx531, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx534, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx537, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx540, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx544, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx547, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx551, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx554, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx558, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx561, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx565, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx568, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_WindowCellShiftedLeft_16, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_16, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_15, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_14, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_13, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_12, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_11, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_10, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_16, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_15, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_14, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_13, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_12, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_11, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_10, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_9, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_8, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_7, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_6, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_5, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_4, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_3, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_2, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_1, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_0, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_16, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_15, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_14, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_13, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_12, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_11, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_10, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_9, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_8, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_7, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_6, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_5, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_4, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_3, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_2, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_1, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_0, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_16, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_15, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_14, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_13, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_12, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_11, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_10, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_9, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_8, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_7, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_6, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_5, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_4, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_3, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_2, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_1, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_0, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx4, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx8, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx12, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx16, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx20, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx24, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx80, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx328, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx384, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642, 
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_AddPToBoothOperand, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothOperand_16, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothOperand_15, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothOperand_14, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothOperand_13, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothOperand_12, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothOperand_11, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothOperand_10, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothOperand_9, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothOperand_8, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothOperand_7, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothOperand_6, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothOperand_5, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothOperand_4, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothOperand_3, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothOperand_2, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothOperand_1, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothOperand_0, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_16, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_15, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_14, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_13, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_12, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_11, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_10, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_9, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_8, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_7, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_6, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_5, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_4, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_3, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_2, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_1, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_16, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_15, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_14, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_13, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_12, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_11, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_10, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_9, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_8, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_7, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_6, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_5, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_4, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_3, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_2, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_1, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_0, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx154, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx316, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx336, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx356, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx376, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx396, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx416, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx436, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx454, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx456, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx379, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx381, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx383, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx387, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx389, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx391, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx395, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx399, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx401, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx403, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx405, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx409, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx411, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx413, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx415, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx419, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx421, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx423, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx425, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx429, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx431, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx433, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx435, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx439, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx441, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx443, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx445, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx449, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx451, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx453, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx455, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx461, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx463, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx467, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx469, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx471, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx475, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx477, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx479, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx483, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx485, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx487, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx491, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx493, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx495, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx499, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx501, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx503, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx507, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx509, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx511, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx515, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx517, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_WindowCellShiftedLeft_16, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_16, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_15, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_14, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_13, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_12, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_11, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_10, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_16, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_15, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_14, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_13, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_12, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_11, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_10, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_9, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_8, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_7, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_6, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_5, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_4, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_3, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_2, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_1, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_0, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_16, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_15, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_14, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_13, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_12, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_11, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_10, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_9, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_8, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_7, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_6, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_5, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_4, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_3, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_2, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_1, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_0, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_16, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_15, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_14, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_13, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_12, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_11, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_10, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_9, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_8, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_7, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_6, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_5, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_4, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_3, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_2, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_1, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_0, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx4, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx8, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx12, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx16, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx20, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx24, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx80, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx328, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx384, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642, 
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_AddPToBoothOperand, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothOperand_16, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothOperand_15, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothOperand_14, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothOperand_13, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothOperand_12, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothOperand_11, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothOperand_10, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothOperand_9, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothOperand_8, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothOperand_7, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothOperand_6, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothOperand_5, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothOperand_4, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothOperand_3, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothOperand_2, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothOperand_1, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothOperand_0, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_16, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_15, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_14, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_13, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_12, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_11, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_10, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_9, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_8, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_7, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_6, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_5, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_4, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_3, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_2, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_1, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_16, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_15, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_14, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_13, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_12, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_11, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_10, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_9, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_8, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_7, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_6, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_5, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_4, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_3, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_2, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_1, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_0, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx0, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx6, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx12, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx18, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx24, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx30, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx40, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx44, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx48, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx52, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx56, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx62, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx154, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx316, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx336, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx356, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx376, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx396, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx416, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx436, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx454, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx456, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx379, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx381, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx383, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx387, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx389, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx391, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx395, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx399, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx401, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx403, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx405, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx409, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx411, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx413, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx415, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx419, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx421, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx423, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx425, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx429, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx431, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx433, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx435, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx439, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx441, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx443, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx445, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx449, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx451, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx453, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx455, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx461, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx463, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx467, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx469, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx471, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx475, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx477, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx479, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx483, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx485, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx487, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx491, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx493, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx495, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx499, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx501, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx503, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx507, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx509, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx511, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx515, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx517, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx529, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx531, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx534, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx537, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx540, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx544, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx547, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx551, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx554, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx558, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx561, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx565, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx568, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_WindowCellShiftedLeft_16, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_16, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_15, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_14, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_13, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_12, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_11, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_10, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_16, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_15, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_14, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_13, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_12, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_11, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_10, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_9, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_8, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_7, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_6, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_5, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_4, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_3, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_2, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_1, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_0, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_16, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_15, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_14, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_13, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_12, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_11, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_10, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_9, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_8, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_7, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_6, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_5, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_4, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_3, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_2, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_1, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_0, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_16, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_15, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_14, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_13, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_12, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_11, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_10, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_9, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_8, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_7, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_6, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_5, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_4, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_3, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_2, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_1, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_0, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx4, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx8, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx12, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx16, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx20, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx24, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx80, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx328, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx384, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642, 
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_AddPToBoothOperand, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothOperand_16, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothOperand_15, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothOperand_14, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothOperand_13, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothOperand_12, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothOperand_11, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothOperand_10, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothOperand_9, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothOperand_8, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothOperand_7, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothOperand_6, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothOperand_5, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothOperand_4, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothOperand_3, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothOperand_2, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothOperand_1, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothOperand_0, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_16, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_15, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_14, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_13, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_12, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_11, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_10, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_9, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_8, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_7, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_6, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_5, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_4, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_3, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_2, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_1, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_16, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_15, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_14, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_13, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_12, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_11, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_10, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_9, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_8, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_7, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_6, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_5, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_4, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_3, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_2, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_1, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_0, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx0, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx6, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx12, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx18, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx24, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx30, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx40, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx44, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx48, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx52, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx56, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx62, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx154, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx316, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx336, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx356, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx376, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx396, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx416, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx436, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx454, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx456, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx379, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx381, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx383, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx387, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx389, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx391, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx395, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx399, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx401, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx403, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx405, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx409, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx411, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx413, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx415, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx419, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx421, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx423, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx425, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx429, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx431, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx433, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx435, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx439, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx441, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx443, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx445, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx449, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx451, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx453, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx455, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx461, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx463, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx467, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx469, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx471, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx475, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx477, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx479, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx483, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx485, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx487, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx491, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx493, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx495, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx499, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx501, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx503, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx507, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx509, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx511, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx515, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx517, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx529, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx531, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx534, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx537, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx540, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx544, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx547, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx551, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx554, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx558, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx561, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx565, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx568, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_WindowCellShiftedLeft_16, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_16, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_15, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_14, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_13, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_12, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_11, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_10, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_16, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_15, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_14, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_13, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_12, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_11, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_10, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_9, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_8, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_7, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_6, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_5, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_4, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_3, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_2, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_1, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_0, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_16, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_15, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_14, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_13, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_12, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_11, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_10, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_9, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_8, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_7, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_6, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_5, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_4, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_3, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_2, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_1, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_0, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_16, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_15, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_14, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_13, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_12, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_11, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_10, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_9, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_8, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_7, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_6, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_5, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_4, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_3, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_2, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_1, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_0, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_nx4, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_nx8, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_nx12, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_nx16, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_nx20, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_nx24, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_nx80, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_nx328, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_nx384, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642, 
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_AddPToBoothOperand, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothOperand_16, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothOperand_15, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothOperand_14, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothOperand_13, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothOperand_12, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothOperand_11, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothOperand_10, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothOperand_9, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothOperand_8, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothOperand_7, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothOperand_6, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothOperand_5, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothOperand_4, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothOperand_3, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothOperand_2, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothOperand_1, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothOperand_0, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_16, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_15, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_14, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_13, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_12, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_11, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_10, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_9, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_8, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_7, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_6, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_5, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_4, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_3, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_2, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_1, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_16, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_15, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_14, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_13, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_12, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_11, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_10, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_9, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_8, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_7, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_6, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_5, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_4, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_3, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_2, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_1, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_0, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx0, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx6, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx12, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx18, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx24, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx30, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx40, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx44, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx48, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx52, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx56, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx62, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx154, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx316, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx336, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx356, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx376, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx396, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx416, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx436, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx454, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx456, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx379, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx381, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx383, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx387, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx389, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx391, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx395, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx399, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx401, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx403, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx405, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx409, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx411, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx413, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx415, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx419, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx421, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx423, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx425, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx429, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx431, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx433, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx435, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx439, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx441, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx443, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx445, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx449, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx451, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx453, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx455, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx461, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx463, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx467, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx469, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx471, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx475, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx477, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx479, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx483, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx485, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx487, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx491, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx493, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx495, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx499, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx501, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx503, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx507, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx509, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx511, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx515, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx517, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx529, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx531, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx534, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx537, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx540, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx544, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx547, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx551, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx554, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx558, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx561, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx565, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx568, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_WindowCellShiftedLeft_16, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_16, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_15, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_14, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_13, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_12, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_11, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_10, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_16, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_15, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_14, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_13, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_12, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_11, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_10, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_9, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_8, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_7, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_6, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_5, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_4, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_3, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_2, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_1, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_0, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_16, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_15, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_14, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_13, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_12, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_11, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_10, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_9, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_8, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_7, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_6, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_5, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_4, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_3, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_2, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_1, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_0, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_16, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_15, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_14, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_13, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_12, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_11, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_10, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_9, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_8, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_7, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_6, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_5, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_4, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_3, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_2, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_1, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_0, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_nx4, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_nx8, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_nx12, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_nx16, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_nx20, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_nx24, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_nx80, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_nx328, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_nx384, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642, 
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_AddPToBoothOperand, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothOperand_16, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothOperand_15, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothOperand_14, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothOperand_13, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothOperand_12, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothOperand_11, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothOperand_10, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothOperand_9, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothOperand_8, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothOperand_7, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothOperand_6, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothOperand_5, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothOperand_4, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothOperand_3, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothOperand_2, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothOperand_1, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothOperand_0, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_16, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_15, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_14, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_13, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_12, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_11, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_10, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_9, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_8, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_7, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_6, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_5, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_4, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_3, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_2, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_1, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_16, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_15, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_14, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_13, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_12, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_11, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_10, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_9, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_8, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_7, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_6, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_5, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_4, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_3, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_2, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_1, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_0, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx0, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx6, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx12, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx18, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx24, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx30, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx40, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx44, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx48, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx52, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx56, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx62, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx154, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx316, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx336, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx356, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx376, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx396, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx416, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx436, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx454, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx456, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx379, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx381, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx383, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx387, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx389, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx391, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx395, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx399, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx401, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx403, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx405, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx409, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx411, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx413, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx415, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx419, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx421, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx423, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx425, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx429, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx431, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx433, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx435, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx439, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx441, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx443, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx445, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx449, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx451, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx453, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx455, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx461, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx463, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx467, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx469, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx471, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx475, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx477, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx479, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx483, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx485, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx487, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx491, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx493, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx495, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx499, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx501, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx503, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx507, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx509, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx511, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx515, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx517, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx529, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx531, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx534, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx537, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx540, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx544, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx547, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx551, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx554, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx558, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx561, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx565, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx568, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_WindowCellShiftedLeft_16, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_16, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_15, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_14, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_13, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_12, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_11, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_10, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_16, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_15, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_14, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_13, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_12, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_11, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_10, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_9, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_8, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_7, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_6, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_5, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_4, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_3, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_2, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_1, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_0, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_16, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_15, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_14, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_13, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_12, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_11, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_10, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_9, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_8, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_7, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_6, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_5, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_4, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_3, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_2, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_1, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_0, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_16, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_15, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_14, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_13, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_12, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_11, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_10, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_9, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_8, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_7, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_6, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_5, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_4, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_3, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_2, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_1, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_0, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_nx4, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_nx8, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_nx12, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_nx16, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_nx20, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_nx24, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_nx80, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_nx328, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_nx384, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642, 
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_AddPToBoothOperand, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothOperand_16, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothOperand_15, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothOperand_14, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothOperand_13, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothOperand_12, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothOperand_11, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothOperand_10, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothOperand_9, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothOperand_8, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothOperand_7, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothOperand_6, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothOperand_5, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothOperand_4, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothOperand_3, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothOperand_2, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothOperand_1, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothOperand_0, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_16, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_15, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_14, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_13, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_12, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_11, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_10, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_9, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_8, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_7, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_6, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_5, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_4, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_3, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_2, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_1, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_16, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_15, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_14, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_13, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_12, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_11, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_10, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_9, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_8, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_7, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_6, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_5, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_4, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_3, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_2, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_1, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_0, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx0, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx6, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx12, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx18, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx24, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx30, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx40, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx44, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx48, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx52, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx56, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx62, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx154, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx316, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx336, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx356, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx376, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx396, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx416, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx436, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx454, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx456, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx379, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx381, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx383, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx387, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx389, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx391, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx395, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx399, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx401, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx403, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx405, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx409, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx411, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx413, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx415, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx419, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx421, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx423, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx425, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx429, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx431, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx433, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx435, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx439, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx441, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx443, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx445, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx449, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx451, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx453, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx455, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx461, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx463, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx467, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx469, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx471, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx475, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx477, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx479, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx483, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx485, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx487, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx491, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx493, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx495, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx499, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx501, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx503, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx507, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx509, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx511, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx515, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx517, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx529, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx531, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx534, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx537, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx540, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx544, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx547, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx551, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx554, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx558, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx561, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx565, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx568, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_WindowCellShiftedLeft_16, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_16, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_15, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_14, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_13, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_12, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_11, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_10, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_16, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_15, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_14, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_13, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_12, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_11, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_10, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_9, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_8, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_7, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_6, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_5, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_4, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_3, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_2, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_1, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_0, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_16, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_15, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_14, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_13, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_12, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_11, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_10, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_9, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_8, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_7, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_6, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_5, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_4, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_3, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_2, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_1, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_0, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_16, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_15, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_14, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_13, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_12, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_11, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_10, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_9, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_8, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_7, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_6, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_5, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_4, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_3, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_2, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_1, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_0, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_nx4, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_nx8, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_nx12, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_nx16, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_nx20, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_nx24, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_nx80, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_nx328, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_nx384, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642, 
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_AddPToBoothOperand, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothOperand_16, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothOperand_15, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothOperand_14, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothOperand_13, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothOperand_12, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothOperand_11, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothOperand_10, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothOperand_9, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothOperand_8, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothOperand_7, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothOperand_6, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothOperand_5, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothOperand_4, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothOperand_3, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothOperand_2, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothOperand_1, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothOperand_0, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_16, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_15, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_14, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_13, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_12, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_11, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_10, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_9, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_8, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_7, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_6, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_5, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_4, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_3, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_2, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_1, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_16, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_15, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_14, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_13, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_12, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_11, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_10, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_9, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_8, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_7, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_6, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_5, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_4, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_3, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_2, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_1, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_0, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx0, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx6, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx12, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx18, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx24, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx30, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx40, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx44, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx48, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx52, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx56, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx62, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx154, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx316, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx336, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx356, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx376, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx396, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx416, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx436, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx454, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx456, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx379, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx381, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx383, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx387, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx389, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx391, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx395, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx399, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx401, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx403, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx405, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx409, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx411, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx413, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx415, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx419, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx421, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx423, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx425, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx429, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx431, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx433, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx435, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx439, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx441, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx443, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx445, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx449, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx451, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx453, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx455, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx461, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx463, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx467, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx469, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx471, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx475, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx477, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx479, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx483, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx485, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx487, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx491, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx493, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx495, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx499, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx501, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx503, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx507, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx509, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx511, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx515, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx517, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx529, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx531, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx534, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx537, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx540, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx544, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx547, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx551, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx554, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx558, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx561, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx565, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx568, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_WindowCellShiftedLeft_16, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_16, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_15, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_14, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_13, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_12, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_11, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_10, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_16, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_15, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_14, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_13, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_12, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_11, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_10, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_9, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_8, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_7, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_6, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_5, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_4, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_3, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_2, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_1, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_0, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_16, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_15, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_14, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_13, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_12, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_11, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_10, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_9, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_8, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_7, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_6, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_5, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_4, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_3, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_2, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_1, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_0, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_16, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_15, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_14, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_13, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_12, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_11, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_10, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_9, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_8, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_7, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_6, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_5, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_4, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_3, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_2, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_1, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_0, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx4, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx8, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx12, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx16, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx20, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx24, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx80, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx328, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx384, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642, 
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_AddPToBoothOperand, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothOperand_16, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothOperand_15, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothOperand_14, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothOperand_13, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothOperand_12, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothOperand_11, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothOperand_10, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothOperand_9, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothOperand_8, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothOperand_7, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothOperand_6, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothOperand_5, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothOperand_4, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothOperand_3, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothOperand_2, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothOperand_1, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothOperand_0, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_16, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_15, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_14, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_13, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_12, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_11, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_10, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_9, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_8, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_7, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_6, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_5, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_4, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_3, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_2, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_1, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_16, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_15, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_14, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_13, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_12, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_11, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_10, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_9, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_8, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_7, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_6, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_5, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_4, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_3, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_2, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_1, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_0, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx0, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx6, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx12, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx18, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx24, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx30, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx40, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx44, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx48, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx52, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx56, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx62, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx154, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx316, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx336, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx356, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx376, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx396, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx416, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx436, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx454, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx456, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx379, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx381, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx383, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx387, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx389, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx391, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx395, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx399, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx401, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx403, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx405, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx409, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx411, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx413, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx415, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx419, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx421, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx423, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx425, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx429, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx431, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx433, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx435, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx439, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx441, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx443, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx445, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx449, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx451, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx453, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx455, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx461, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx463, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx467, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx469, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx471, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx475, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx477, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx479, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx483, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx485, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx487, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx491, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx493, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx495, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx499, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx501, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx503, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx507, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx509, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx511, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx515, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx517, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx529, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx531, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx534, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx537, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx540, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx544, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx547, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx551, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx554, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx558, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx561, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx565, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx568, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_WindowCellShiftedLeft_16, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_16, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_15, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_14, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_13, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_12, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_11, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_10, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_16, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_15, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_14, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_13, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_12, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_11, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_10, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_9, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_8, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_7, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_6, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_5, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_4, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_3, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_2, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_1, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_0, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_16, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_15, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_14, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_13, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_12, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_11, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_10, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_9, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_8, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_7, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_6, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_5, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_4, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_3, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_2, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_1, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_0, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_16, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_15, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_14, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_13, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_12, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_11, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_10, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_9, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_8, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_7, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_6, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_5, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_4, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_3, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_2, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_1, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_0, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_nx4, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_nx8, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_nx12, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_nx16, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_nx20, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_nx24, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_nx80, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_nx328, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_nx384, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642, 
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_AddPToBoothOperand, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothOperand_16, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothOperand_15, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothOperand_14, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothOperand_13, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothOperand_12, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothOperand_11, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothOperand_10, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothOperand_9, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothOperand_8, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothOperand_7, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothOperand_6, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothOperand_5, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothOperand_4, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothOperand_3, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothOperand_2, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothOperand_1, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothOperand_0, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_16, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_15, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_14, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_13, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_12, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_11, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_10, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_9, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_8, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_7, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_6, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_5, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_4, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_3, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_2, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_1, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_16, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_15, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_14, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_13, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_12, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_11, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_10, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_9, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_8, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_7, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_6, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_5, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_4, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_3, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_2, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_1, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_0, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx0, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx6, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx12, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx18, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx24, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx30, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx40, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx44, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx48, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx52, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx56, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx62, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx154, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx316, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx336, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx356, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx376, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx396, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx416, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx436, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx454, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx456, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx379, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx381, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx383, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx387, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx389, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx391, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx395, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx399, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx401, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx403, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx405, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx409, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx411, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx413, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx415, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx419, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx421, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx423, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx425, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx429, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx431, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx433, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx435, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx439, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx441, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx443, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx445, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx449, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx451, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx453, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx455, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx461, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx463, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx467, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx469, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx471, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx475, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx477, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx479, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx483, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx485, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx487, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx491, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx493, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx495, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx499, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx501, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx503, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx507, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx509, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx511, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx515, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx517, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx529, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx531, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx534, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx537, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx540, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx544, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx547, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx551, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx554, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx558, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx561, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx565, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx568, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_WindowCellShiftedLeft_16, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_16, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_15, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_14, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_13, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_12, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_11, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_10, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_16, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_15, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_14, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_13, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_12, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_11, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_10, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_9, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_8, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_7, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_6, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_5, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_4, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_3, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_2, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_1, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_0, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_16, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_15, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_14, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_13, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_12, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_11, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_10, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_9, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_8, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_7, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_6, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_5, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_4, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_3, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_2, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_1, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_0, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_16, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_15, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_14, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_13, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_12, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_11, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_10, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_9, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_8, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_7, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_6, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_5, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_4, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_3, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_2, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_1, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_0, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_nx4, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_nx8, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_nx12, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_nx16, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_nx20, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_nx24, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_nx80, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_nx328, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_nx384, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642, 
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_AddPToBoothOperand, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothOperand_16, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothOperand_15, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothOperand_14, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothOperand_13, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothOperand_12, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothOperand_11, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothOperand_10, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothOperand_9, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothOperand_8, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothOperand_7, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothOperand_6, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothOperand_5, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothOperand_4, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothOperand_3, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothOperand_2, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothOperand_1, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothOperand_0, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_16, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_15, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_14, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_13, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_12, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_11, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_10, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_9, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_8, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_7, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_6, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_5, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_4, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_3, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_2, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_1, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_16, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_15, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_14, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_13, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_12, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_11, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_10, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_9, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_8, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_7, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_6, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_5, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_4, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_3, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_2, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_1, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_0, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx0, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx6, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx12, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx18, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx24, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx30, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx40, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx44, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx48, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx52, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx56, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx62, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx154, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx316, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx336, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx356, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx376, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx396, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx416, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx436, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx454, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx456, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx379, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx381, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx383, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx387, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx389, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx391, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx395, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx399, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx401, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx403, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx405, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx409, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx411, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx413, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx415, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx419, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx421, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx423, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx425, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx429, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx431, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx433, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx435, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx439, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx441, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx443, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx445, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx449, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx451, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx453, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx455, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx461, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx463, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx467, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx469, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx471, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx475, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx477, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx479, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx483, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx485, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx487, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx491, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx493, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx495, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx499, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx501, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx503, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx507, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx509, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx511, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx515, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx517, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx529, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx531, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx534, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx537, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx540, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx544, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx547, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx551, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx554, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx558, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx561, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx565, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx568, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_WindowCellShiftedLeft_16, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_16, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_15, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_14, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_13, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_12, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_11, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_10, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_16, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_15, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_14, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_13, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_12, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_11, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_10, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_9, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_8, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_7, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_6, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_5, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_4, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_3, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_2, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_1, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_0, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_16, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_15, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_14, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_13, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_12, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_11, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_10, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_9, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_8, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_7, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_6, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_5, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_4, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_3, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_2, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_1, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_0, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_16, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_15, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_14, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_13, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_12, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_11, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_10, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_9, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_8, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_7, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_6, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_5, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_4, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_3, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_2, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_1, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_0, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_nx4, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_nx8, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_nx12, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_nx16, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_nx20, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_nx24, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_nx80, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_nx328, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_nx384, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642, 
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_AddPToBoothOperand, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothOperand_16, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothOperand_15, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothOperand_14, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothOperand_13, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothOperand_12, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothOperand_11, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothOperand_10, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothOperand_9, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothOperand_8, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothOperand_7, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothOperand_6, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothOperand_5, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothOperand_4, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothOperand_3, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothOperand_2, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothOperand_1, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothOperand_0, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_16, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_15, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_14, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_13, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_12, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_11, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_10, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_9, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_8, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_7, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_6, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_5, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_4, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_3, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_2, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_1, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_16, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_15, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_14, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_13, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_12, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_11, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_10, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_9, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_8, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_7, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_6, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_5, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_4, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_3, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_2, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_1, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_0, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx0, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx6, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx12, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx18, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx24, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx30, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx40, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx44, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx48, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx52, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx56, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx62, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx154, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx316, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx336, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx356, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx376, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx396, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx416, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx436, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx454, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx456, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx379, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx381, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx383, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx387, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx389, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx391, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx395, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx399, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx401, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx403, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx405, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx409, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx411, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx413, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx415, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx419, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx421, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx423, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx425, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx429, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx431, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx433, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx435, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx439, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx441, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx443, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx445, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx449, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx451, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx453, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx455, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx461, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx463, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx467, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx469, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx471, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx475, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx477, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx479, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx483, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx485, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx487, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx491, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx493, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx495, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx499, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx501, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx503, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx507, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx509, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx511, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx515, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx517, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx529, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx531, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx534, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx537, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx540, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx544, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx547, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx551, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx554, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx558, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx561, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx565, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx568, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_WindowCellShiftedLeft_16, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDin_16, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDin_15, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDin_14, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDin_13, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDin_12, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDin_11, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDin_10, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_16, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_15, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_14, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_13, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_12, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_11, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_10, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_9, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_8, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_7, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_6, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_5, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_4, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_3, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_2, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_1, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_0, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_16, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_15, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_14, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_13, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_12, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_11, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_10, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_9, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_8, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_7, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_6, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_5, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_4, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_3, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_2, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_1, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_0, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_16, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_15, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_14, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_13, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_12, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_11, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_10, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_9, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_8, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_7, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_6, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_5, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_4, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_3, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_2, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_1, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_0, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_nx4, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_nx8, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_nx12, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_nx16, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_nx20, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_nx24, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_nx80, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_nx328, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_nx384, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642, 
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_AddPToBoothOperand, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothOperand_16, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothOperand_15, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothOperand_14, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothOperand_13, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothOperand_12, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothOperand_11, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothOperand_10, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothOperand_9, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothOperand_8, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothOperand_7, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothOperand_6, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothOperand_5, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothOperand_4, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothOperand_3, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothOperand_2, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothOperand_1, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothOperand_0, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_16, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_15, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_14, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_13, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_12, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_11, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_10, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_9, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_8, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_7, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_6, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_5, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_4, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_3, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_2, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_1, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_16, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_15, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_14, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_13, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_12, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_11, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_10, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_9, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_8, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_7, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_6, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_5, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_4, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_3, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_2, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_1, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_0, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx0, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx6, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx12, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx18, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx24, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx30, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx40, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx44, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx48, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx52, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx56, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx62, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx154, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx316, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx336, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx356, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx376, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx396, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx416, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx436, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx454, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx456, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx379, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx381, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx383, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx387, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx389, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx391, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx395, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx399, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx401, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx403, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx405, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx409, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx411, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx413, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx415, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx419, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx421, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx423, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx425, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx429, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx431, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx433, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx435, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx439, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx441, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx443, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx445, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx449, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx451, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx453, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx455, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx461, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx463, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx467, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx469, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx471, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx475, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx477, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx479, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx483, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx485, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx487, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx491, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx493, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx495, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx499, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx501, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx503, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx507, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx509, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx511, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx515, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx517, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx529, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx531, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx534, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx537, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx540, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx544, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx547, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx551, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx554, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx558, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx561, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx565, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx568, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_WindowCellShiftedLeft_16, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_16, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_15, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_14, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_13, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_12, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_11, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_10, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_16, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_15, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_14, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_13, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_12, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_11, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_10, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_9, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_8, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_7, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_6, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_5, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_4, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_3, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_2, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_1, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_0, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_16, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_15, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_14, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_13, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_12, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_11, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_10, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_9, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_8, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_7, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_6, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_5, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_4, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_3, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_2, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_1, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_0, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_16, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_15, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_14, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_13, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_12, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_11, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_10, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_9, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_8, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_7, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_6, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_5, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_4, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_3, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_2, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_1, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_0, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_nx4, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_nx8, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_nx12, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_nx16, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_nx20, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_nx24, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_nx80, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_nx328, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_nx384, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642, 
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_AddPToBoothOperand, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothOperand_16, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothOperand_15, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothOperand_14, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothOperand_13, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothOperand_12, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothOperand_11, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothOperand_10, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothOperand_9, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothOperand_8, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothOperand_7, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothOperand_6, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothOperand_5, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothOperand_4, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothOperand_3, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothOperand_2, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothOperand_1, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothOperand_0, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_16, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_15, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_14, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_13, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_12, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_11, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_10, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_9, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_8, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_7, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_6, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_5, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_4, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_3, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_2, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_1, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_16, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_15, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_14, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_13, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_12, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_11, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_10, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_9, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_8, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_7, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_6, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_5, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_4, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_3, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_2, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_1, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_0, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx0, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx6, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx12, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx18, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx24, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx30, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx40, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx44, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx48, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx52, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx56, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx62, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx154, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx316, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx336, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx356, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx376, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx396, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx416, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx436, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx454, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx456, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx379, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx381, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx383, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx387, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx389, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx391, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx395, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx399, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx401, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx403, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx405, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx409, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx411, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx413, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx415, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx419, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx421, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx423, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx425, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx429, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx431, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx433, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx435, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx439, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx441, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx443, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx445, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx449, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx451, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx453, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx455, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx461, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx463, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx467, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx469, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx471, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx475, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx477, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx479, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx483, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx485, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx487, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx491, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx493, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx495, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx499, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx501, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx503, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx507, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx509, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx511, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx515, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx517, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx529, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx531, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx534, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx537, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx540, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx544, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx547, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx551, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx554, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx558, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx561, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx565, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx568, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_WindowCellShiftedLeft_16, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_16, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_15, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_14, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_13, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_12, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_11, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_10, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_16, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_15, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_14, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_13, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_12, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_11, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_10, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_9, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_8, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_7, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_6, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_5, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_4, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_3, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_2, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_1, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_0, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_16, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_15, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_14, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_13, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_12, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_11, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_10, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_9, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_8, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_7, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_6, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_5, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_4, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_3, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_2, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_1, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_0, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_16, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_15, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_14, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_13, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_12, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_11, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_10, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_9, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_8, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_7, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_6, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_5, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_4, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_3, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_2, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_1, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_0, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_nx4, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_nx8, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_nx12, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_nx16, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_nx20, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_nx24, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_nx80, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_nx328, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_nx384, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642, 
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644, 
         CACHE_nx941, CACHE_EN_dup_1491, CACHE_EN_dup_1359, CACHE_EN_dup_1227, 
         CACHE_EN_dup_1161, CACHE_EN_dup_1095, CACHE_EN, CACHE_nx955, 
         CACHE_EN_dup_1502, CACHE_EN_dup_1370, CACHE_EN_dup_1238, 
         CACHE_EN_dup_1172, CACHE_EN_dup_1106, CACHE_EN_dup_1084, 
         CACHE_RST_dup_1073, CACHE_RST_dup_1094, CACHE_RST_dup_1116, 
         CACHE_RST_dup_1138, CACHE_RST_dup_1160, CACHE_RST_dup_1182, 
         CACHE_RST_dup_1204, CACHE_RST_dup_1226, CACHE_RST_dup_1248, 
         CACHE_RST_dup_1270, CACHE_RST_dup_1292, CACHE_RST_dup_1314, 
         CACHE_RST_dup_1336, CACHE_RST_dup_1358, CACHE_RST_dup_1380, 
         CACHE_RST_dup_1402, CACHE_RST_dup_1424, CACHE_RST_dup_1446, 
         CACHE_RST_dup_1468, CACHE_RST_dup_1490, CACHE_RST_dup_1512, 
         CACHE_RST_dup_1534, CACHE_RST_dup_1556, CACHE_RST_dup_1578, 
         CACHE_RST_dup_1600, CACHE_nx1025, CACHE_EN_dup_1293, CACHE_EN_dup_1403, 
         CACHE_EN_dup_1513, CACHE_nx1033, CACHE_EN_dup_1304, CACHE_EN_dup_1414, 
         CACHE_EN_dup_1524, CACHE_nx1041, CACHE_nx1043, CACHE_nx1045, 
         CACHE_nx1047, CACHE_L0_0_L1_0_Fij_nx212, CACHE_L0_0_L1_0_Fij_nx222, 
         CACHE_L0_0_L1_0_Fij_nx232, CACHE_L0_0_L1_0_Fij_nx242, 
         CACHE_L0_0_L1_0_Fij_nx252, CACHE_L0_0_L1_0_Fij_nx262, 
         CACHE_L0_0_L1_0_Fij_nx272, CACHE_L0_0_L1_0_Fij_nx282, 
         CACHE_L0_0_L1_0_Fij_nx296, CACHE_L0_0_L1_0_Fij_nx331, 
         CACHE_L0_0_L1_0_Fij_nx333, CACHE_L0_0_L1_0_Wij_nx212, 
         CACHE_L0_0_L1_0_Wij_nx222, CACHE_L0_0_L1_0_Wij_nx232, 
         CACHE_L0_0_L1_0_Wij_nx242, CACHE_L0_0_L1_0_Wij_nx252, 
         CACHE_L0_0_L1_0_Wij_nx262, CACHE_L0_0_L1_0_Wij_nx272, 
         CACHE_L0_0_L1_0_Wij_nx282, CACHE_L0_0_L1_0_Wij_nx296, 
         CACHE_L0_0_L1_0_Wij_nx331, CACHE_L0_0_L1_0_Wij_nx333, 
         CACHE_L0_0_L1_1_Fij_nx212, CACHE_L0_0_L1_1_Fij_nx222, 
         CACHE_L0_0_L1_1_Fij_nx232, CACHE_L0_0_L1_1_Fij_nx242, 
         CACHE_L0_0_L1_1_Fij_nx252, CACHE_L0_0_L1_1_Fij_nx262, 
         CACHE_L0_0_L1_1_Fij_nx272, CACHE_L0_0_L1_1_Fij_nx282, 
         CACHE_L0_0_L1_1_Fij_nx296, CACHE_L0_0_L1_1_Fij_nx331, 
         CACHE_L0_0_L1_1_Fij_nx333, CACHE_L0_0_L1_1_Wij_nx212, 
         CACHE_L0_0_L1_1_Wij_nx222, CACHE_L0_0_L1_1_Wij_nx232, 
         CACHE_L0_0_L1_1_Wij_nx242, CACHE_L0_0_L1_1_Wij_nx252, 
         CACHE_L0_0_L1_1_Wij_nx262, CACHE_L0_0_L1_1_Wij_nx272, 
         CACHE_L0_0_L1_1_Wij_nx282, CACHE_L0_0_L1_1_Wij_nx296, 
         CACHE_L0_0_L1_1_Wij_nx331, CACHE_L0_0_L1_1_Wij_nx333, 
         CACHE_L0_0_L1_2_Fij_nx212, CACHE_L0_0_L1_2_Fij_nx222, 
         CACHE_L0_0_L1_2_Fij_nx232, CACHE_L0_0_L1_2_Fij_nx242, 
         CACHE_L0_0_L1_2_Fij_nx252, CACHE_L0_0_L1_2_Fij_nx262, 
         CACHE_L0_0_L1_2_Fij_nx272, CACHE_L0_0_L1_2_Fij_nx282, 
         CACHE_L0_0_L1_2_Fij_nx296, CACHE_L0_0_L1_2_Fij_nx331, 
         CACHE_L0_0_L1_2_Fij_nx333, CACHE_L0_0_L1_2_Wij_nx212, 
         CACHE_L0_0_L1_2_Wij_nx222, CACHE_L0_0_L1_2_Wij_nx232, 
         CACHE_L0_0_L1_2_Wij_nx242, CACHE_L0_0_L1_2_Wij_nx252, 
         CACHE_L0_0_L1_2_Wij_nx262, CACHE_L0_0_L1_2_Wij_nx272, 
         CACHE_L0_0_L1_2_Wij_nx282, CACHE_L0_0_L1_2_Wij_nx296, 
         CACHE_L0_0_L1_2_Wij_nx331, CACHE_L0_0_L1_2_Wij_nx333, 
         CACHE_L0_0_L1_3_Fij_nx212, CACHE_L0_0_L1_3_Fij_nx222, 
         CACHE_L0_0_L1_3_Fij_nx232, CACHE_L0_0_L1_3_Fij_nx242, 
         CACHE_L0_0_L1_3_Fij_nx252, CACHE_L0_0_L1_3_Fij_nx262, 
         CACHE_L0_0_L1_3_Fij_nx272, CACHE_L0_0_L1_3_Fij_nx282, 
         CACHE_L0_0_L1_3_Fij_nx296, CACHE_L0_0_L1_3_Fij_nx331, 
         CACHE_L0_0_L1_3_Fij_nx333, CACHE_L0_0_L1_3_Wij_nx212, 
         CACHE_L0_0_L1_3_Wij_nx222, CACHE_L0_0_L1_3_Wij_nx232, 
         CACHE_L0_0_L1_3_Wij_nx242, CACHE_L0_0_L1_3_Wij_nx252, 
         CACHE_L0_0_L1_3_Wij_nx262, CACHE_L0_0_L1_3_Wij_nx272, 
         CACHE_L0_0_L1_3_Wij_nx282, CACHE_L0_0_L1_3_Wij_nx296, 
         CACHE_L0_0_L1_3_Wij_nx331, CACHE_L0_0_L1_3_Wij_nx333, 
         CACHE_L0_0_L1_4_Fij_nx212, CACHE_L0_0_L1_4_Fij_nx222, 
         CACHE_L0_0_L1_4_Fij_nx232, CACHE_L0_0_L1_4_Fij_nx242, 
         CACHE_L0_0_L1_4_Fij_nx252, CACHE_L0_0_L1_4_Fij_nx262, 
         CACHE_L0_0_L1_4_Fij_nx272, CACHE_L0_0_L1_4_Fij_nx282, 
         CACHE_L0_0_L1_4_Fij_nx296, CACHE_L0_0_L1_4_Fij_nx331, 
         CACHE_L0_0_L1_4_Fij_nx333, CACHE_L0_0_L1_4_Wij_nx212, 
         CACHE_L0_0_L1_4_Wij_nx222, CACHE_L0_0_L1_4_Wij_nx232, 
         CACHE_L0_0_L1_4_Wij_nx242, CACHE_L0_0_L1_4_Wij_nx252, 
         CACHE_L0_0_L1_4_Wij_nx262, CACHE_L0_0_L1_4_Wij_nx272, 
         CACHE_L0_0_L1_4_Wij_nx282, CACHE_L0_0_L1_4_Wij_nx296, 
         CACHE_L0_0_L1_4_Wij_nx331, CACHE_L0_0_L1_4_Wij_nx333, 
         CACHE_L0_1_L1_0_Fij_nx212, CACHE_L0_1_L1_0_Fij_nx222, 
         CACHE_L0_1_L1_0_Fij_nx232, CACHE_L0_1_L1_0_Fij_nx242, 
         CACHE_L0_1_L1_0_Fij_nx252, CACHE_L0_1_L1_0_Fij_nx262, 
         CACHE_L0_1_L1_0_Fij_nx272, CACHE_L0_1_L1_0_Fij_nx282, 
         CACHE_L0_1_L1_0_Fij_nx296, CACHE_L0_1_L1_0_Fij_nx331, 
         CACHE_L0_1_L1_0_Fij_nx333, CACHE_L0_1_L1_0_Wij_nx212, 
         CACHE_L0_1_L1_0_Wij_nx222, CACHE_L0_1_L1_0_Wij_nx232, 
         CACHE_L0_1_L1_0_Wij_nx242, CACHE_L0_1_L1_0_Wij_nx252, 
         CACHE_L0_1_L1_0_Wij_nx262, CACHE_L0_1_L1_0_Wij_nx272, 
         CACHE_L0_1_L1_0_Wij_nx282, CACHE_L0_1_L1_0_Wij_nx296, 
         CACHE_L0_1_L1_0_Wij_nx331, CACHE_L0_1_L1_0_Wij_nx333, 
         CACHE_L0_1_L1_1_Fij_nx212, CACHE_L0_1_L1_1_Fij_nx222, 
         CACHE_L0_1_L1_1_Fij_nx232, CACHE_L0_1_L1_1_Fij_nx242, 
         CACHE_L0_1_L1_1_Fij_nx252, CACHE_L0_1_L1_1_Fij_nx262, 
         CACHE_L0_1_L1_1_Fij_nx272, CACHE_L0_1_L1_1_Fij_nx282, 
         CACHE_L0_1_L1_1_Fij_nx296, CACHE_L0_1_L1_1_Fij_nx331, 
         CACHE_L0_1_L1_1_Fij_nx333, CACHE_L0_1_L1_1_Wij_nx212, 
         CACHE_L0_1_L1_1_Wij_nx222, CACHE_L0_1_L1_1_Wij_nx232, 
         CACHE_L0_1_L1_1_Wij_nx242, CACHE_L0_1_L1_1_Wij_nx252, 
         CACHE_L0_1_L1_1_Wij_nx262, CACHE_L0_1_L1_1_Wij_nx272, 
         CACHE_L0_1_L1_1_Wij_nx282, CACHE_L0_1_L1_1_Wij_nx296, 
         CACHE_L0_1_L1_1_Wij_nx331, CACHE_L0_1_L1_1_Wij_nx333, 
         CACHE_L0_1_L1_2_Fij_nx212, CACHE_L0_1_L1_2_Fij_nx222, 
         CACHE_L0_1_L1_2_Fij_nx232, CACHE_L0_1_L1_2_Fij_nx242, 
         CACHE_L0_1_L1_2_Fij_nx252, CACHE_L0_1_L1_2_Fij_nx262, 
         CACHE_L0_1_L1_2_Fij_nx272, CACHE_L0_1_L1_2_Fij_nx282, 
         CACHE_L0_1_L1_2_Fij_nx296, CACHE_L0_1_L1_2_Fij_nx331, 
         CACHE_L0_1_L1_2_Fij_nx333, CACHE_L0_1_L1_2_Wij_nx212, 
         CACHE_L0_1_L1_2_Wij_nx222, CACHE_L0_1_L1_2_Wij_nx232, 
         CACHE_L0_1_L1_2_Wij_nx242, CACHE_L0_1_L1_2_Wij_nx252, 
         CACHE_L0_1_L1_2_Wij_nx262, CACHE_L0_1_L1_2_Wij_nx272, 
         CACHE_L0_1_L1_2_Wij_nx282, CACHE_L0_1_L1_2_Wij_nx296, 
         CACHE_L0_1_L1_2_Wij_nx331, CACHE_L0_1_L1_2_Wij_nx333, 
         CACHE_L0_1_L1_3_Fij_nx212, CACHE_L0_1_L1_3_Fij_nx222, 
         CACHE_L0_1_L1_3_Fij_nx232, CACHE_L0_1_L1_3_Fij_nx242, 
         CACHE_L0_1_L1_3_Fij_nx252, CACHE_L0_1_L1_3_Fij_nx262, 
         CACHE_L0_1_L1_3_Fij_nx272, CACHE_L0_1_L1_3_Fij_nx282, 
         CACHE_L0_1_L1_3_Fij_nx296, CACHE_L0_1_L1_3_Fij_nx331, 
         CACHE_L0_1_L1_3_Fij_nx333, CACHE_L0_1_L1_3_Wij_nx212, 
         CACHE_L0_1_L1_3_Wij_nx222, CACHE_L0_1_L1_3_Wij_nx232, 
         CACHE_L0_1_L1_3_Wij_nx242, CACHE_L0_1_L1_3_Wij_nx252, 
         CACHE_L0_1_L1_3_Wij_nx262, CACHE_L0_1_L1_3_Wij_nx272, 
         CACHE_L0_1_L1_3_Wij_nx282, CACHE_L0_1_L1_3_Wij_nx296, 
         CACHE_L0_1_L1_3_Wij_nx331, CACHE_L0_1_L1_3_Wij_nx333, 
         CACHE_L0_1_L1_4_Fij_nx212, CACHE_L0_1_L1_4_Fij_nx222, 
         CACHE_L0_1_L1_4_Fij_nx232, CACHE_L0_1_L1_4_Fij_nx242, 
         CACHE_L0_1_L1_4_Fij_nx252, CACHE_L0_1_L1_4_Fij_nx262, 
         CACHE_L0_1_L1_4_Fij_nx272, CACHE_L0_1_L1_4_Fij_nx282, 
         CACHE_L0_1_L1_4_Fij_nx296, CACHE_L0_1_L1_4_Fij_nx331, 
         CACHE_L0_1_L1_4_Fij_nx333, CACHE_L0_1_L1_4_Wij_nx212, 
         CACHE_L0_1_L1_4_Wij_nx222, CACHE_L0_1_L1_4_Wij_nx232, 
         CACHE_L0_1_L1_4_Wij_nx242, CACHE_L0_1_L1_4_Wij_nx252, 
         CACHE_L0_1_L1_4_Wij_nx262, CACHE_L0_1_L1_4_Wij_nx272, 
         CACHE_L0_1_L1_4_Wij_nx282, CACHE_L0_1_L1_4_Wij_nx296, 
         CACHE_L0_1_L1_4_Wij_nx331, CACHE_L0_1_L1_4_Wij_nx333, 
         CACHE_L0_2_L1_0_Fij_nx212, CACHE_L0_2_L1_0_Fij_nx222, 
         CACHE_L0_2_L1_0_Fij_nx232, CACHE_L0_2_L1_0_Fij_nx242, 
         CACHE_L0_2_L1_0_Fij_nx252, CACHE_L0_2_L1_0_Fij_nx262, 
         CACHE_L0_2_L1_0_Fij_nx272, CACHE_L0_2_L1_0_Fij_nx282, 
         CACHE_L0_2_L1_0_Fij_nx296, CACHE_L0_2_L1_0_Fij_nx331, 
         CACHE_L0_2_L1_0_Fij_nx333, CACHE_L0_2_L1_0_Wij_nx212, 
         CACHE_L0_2_L1_0_Wij_nx222, CACHE_L0_2_L1_0_Wij_nx232, 
         CACHE_L0_2_L1_0_Wij_nx242, CACHE_L0_2_L1_0_Wij_nx252, 
         CACHE_L0_2_L1_0_Wij_nx262, CACHE_L0_2_L1_0_Wij_nx272, 
         CACHE_L0_2_L1_0_Wij_nx282, CACHE_L0_2_L1_0_Wij_nx296, 
         CACHE_L0_2_L1_0_Wij_nx331, CACHE_L0_2_L1_0_Wij_nx333, 
         CACHE_L0_2_L1_1_Fij_nx212, CACHE_L0_2_L1_1_Fij_nx222, 
         CACHE_L0_2_L1_1_Fij_nx232, CACHE_L0_2_L1_1_Fij_nx242, 
         CACHE_L0_2_L1_1_Fij_nx252, CACHE_L0_2_L1_1_Fij_nx262, 
         CACHE_L0_2_L1_1_Fij_nx272, CACHE_L0_2_L1_1_Fij_nx282, 
         CACHE_L0_2_L1_1_Fij_nx296, CACHE_L0_2_L1_1_Fij_nx331, 
         CACHE_L0_2_L1_1_Fij_nx333, CACHE_L0_2_L1_1_Wij_nx212, 
         CACHE_L0_2_L1_1_Wij_nx222, CACHE_L0_2_L1_1_Wij_nx232, 
         CACHE_L0_2_L1_1_Wij_nx242, CACHE_L0_2_L1_1_Wij_nx252, 
         CACHE_L0_2_L1_1_Wij_nx262, CACHE_L0_2_L1_1_Wij_nx272, 
         CACHE_L0_2_L1_1_Wij_nx282, CACHE_L0_2_L1_1_Wij_nx296, 
         CACHE_L0_2_L1_1_Wij_nx331, CACHE_L0_2_L1_1_Wij_nx333, 
         CACHE_L0_2_L1_2_Fij_nx212, CACHE_L0_2_L1_2_Fij_nx222, 
         CACHE_L0_2_L1_2_Fij_nx232, CACHE_L0_2_L1_2_Fij_nx242, 
         CACHE_L0_2_L1_2_Fij_nx252, CACHE_L0_2_L1_2_Fij_nx262, 
         CACHE_L0_2_L1_2_Fij_nx272, CACHE_L0_2_L1_2_Fij_nx282, 
         CACHE_L0_2_L1_2_Fij_nx296, CACHE_L0_2_L1_2_Fij_nx331, 
         CACHE_L0_2_L1_2_Fij_nx333, CACHE_L0_2_L1_2_Wij_nx212, 
         CACHE_L0_2_L1_2_Wij_nx222, CACHE_L0_2_L1_2_Wij_nx232, 
         CACHE_L0_2_L1_2_Wij_nx242, CACHE_L0_2_L1_2_Wij_nx252, 
         CACHE_L0_2_L1_2_Wij_nx262, CACHE_L0_2_L1_2_Wij_nx272, 
         CACHE_L0_2_L1_2_Wij_nx282, CACHE_L0_2_L1_2_Wij_nx296, 
         CACHE_L0_2_L1_2_Wij_nx331, CACHE_L0_2_L1_2_Wij_nx333, 
         CACHE_L0_2_L1_3_Fij_nx212, CACHE_L0_2_L1_3_Fij_nx222, 
         CACHE_L0_2_L1_3_Fij_nx232, CACHE_L0_2_L1_3_Fij_nx242, 
         CACHE_L0_2_L1_3_Fij_nx252, CACHE_L0_2_L1_3_Fij_nx262, 
         CACHE_L0_2_L1_3_Fij_nx272, CACHE_L0_2_L1_3_Fij_nx282, 
         CACHE_L0_2_L1_3_Fij_nx296, CACHE_L0_2_L1_3_Fij_nx331, 
         CACHE_L0_2_L1_3_Fij_nx333, CACHE_L0_2_L1_3_Wij_nx212, 
         CACHE_L0_2_L1_3_Wij_nx222, CACHE_L0_2_L1_3_Wij_nx232, 
         CACHE_L0_2_L1_3_Wij_nx242, CACHE_L0_2_L1_3_Wij_nx252, 
         CACHE_L0_2_L1_3_Wij_nx262, CACHE_L0_2_L1_3_Wij_nx272, 
         CACHE_L0_2_L1_3_Wij_nx282, CACHE_L0_2_L1_3_Wij_nx296, 
         CACHE_L0_2_L1_3_Wij_nx331, CACHE_L0_2_L1_3_Wij_nx333, 
         CACHE_L0_2_L1_4_Fij_nx212, CACHE_L0_2_L1_4_Fij_nx222, 
         CACHE_L0_2_L1_4_Fij_nx232, CACHE_L0_2_L1_4_Fij_nx242, 
         CACHE_L0_2_L1_4_Fij_nx252, CACHE_L0_2_L1_4_Fij_nx262, 
         CACHE_L0_2_L1_4_Fij_nx272, CACHE_L0_2_L1_4_Fij_nx282, 
         CACHE_L0_2_L1_4_Fij_nx296, CACHE_L0_2_L1_4_Fij_nx331, 
         CACHE_L0_2_L1_4_Fij_nx333, CACHE_L0_2_L1_4_Wij_nx212, 
         CACHE_L0_2_L1_4_Wij_nx222, CACHE_L0_2_L1_4_Wij_nx232, 
         CACHE_L0_2_L1_4_Wij_nx242, CACHE_L0_2_L1_4_Wij_nx252, 
         CACHE_L0_2_L1_4_Wij_nx262, CACHE_L0_2_L1_4_Wij_nx272, 
         CACHE_L0_2_L1_4_Wij_nx282, CACHE_L0_2_L1_4_Wij_nx296, 
         CACHE_L0_2_L1_4_Wij_nx331, CACHE_L0_2_L1_4_Wij_nx333, 
         CACHE_L0_3_L1_0_Fij_nx212, CACHE_L0_3_L1_0_Fij_nx222, 
         CACHE_L0_3_L1_0_Fij_nx232, CACHE_L0_3_L1_0_Fij_nx242, 
         CACHE_L0_3_L1_0_Fij_nx252, CACHE_L0_3_L1_0_Fij_nx262, 
         CACHE_L0_3_L1_0_Fij_nx272, CACHE_L0_3_L1_0_Fij_nx282, 
         CACHE_L0_3_L1_0_Fij_nx296, CACHE_L0_3_L1_0_Fij_nx331, 
         CACHE_L0_3_L1_0_Fij_nx333, CACHE_L0_3_L1_0_Wij_nx212, 
         CACHE_L0_3_L1_0_Wij_nx222, CACHE_L0_3_L1_0_Wij_nx232, 
         CACHE_L0_3_L1_0_Wij_nx242, CACHE_L0_3_L1_0_Wij_nx252, 
         CACHE_L0_3_L1_0_Wij_nx262, CACHE_L0_3_L1_0_Wij_nx272, 
         CACHE_L0_3_L1_0_Wij_nx282, CACHE_L0_3_L1_0_Wij_nx296, 
         CACHE_L0_3_L1_0_Wij_nx331, CACHE_L0_3_L1_0_Wij_nx333, 
         CACHE_L0_3_L1_1_Fij_nx212, CACHE_L0_3_L1_1_Fij_nx222, 
         CACHE_L0_3_L1_1_Fij_nx232, CACHE_L0_3_L1_1_Fij_nx242, 
         CACHE_L0_3_L1_1_Fij_nx252, CACHE_L0_3_L1_1_Fij_nx262, 
         CACHE_L0_3_L1_1_Fij_nx272, CACHE_L0_3_L1_1_Fij_nx282, 
         CACHE_L0_3_L1_1_Fij_nx296, CACHE_L0_3_L1_1_Fij_nx331, 
         CACHE_L0_3_L1_1_Fij_nx333, CACHE_L0_3_L1_1_Wij_nx212, 
         CACHE_L0_3_L1_1_Wij_nx222, CACHE_L0_3_L1_1_Wij_nx232, 
         CACHE_L0_3_L1_1_Wij_nx242, CACHE_L0_3_L1_1_Wij_nx252, 
         CACHE_L0_3_L1_1_Wij_nx262, CACHE_L0_3_L1_1_Wij_nx272, 
         CACHE_L0_3_L1_1_Wij_nx282, CACHE_L0_3_L1_1_Wij_nx296, 
         CACHE_L0_3_L1_1_Wij_nx331, CACHE_L0_3_L1_1_Wij_nx333, 
         CACHE_L0_3_L1_2_Fij_nx212, CACHE_L0_3_L1_2_Fij_nx222, 
         CACHE_L0_3_L1_2_Fij_nx232, CACHE_L0_3_L1_2_Fij_nx242, 
         CACHE_L0_3_L1_2_Fij_nx252, CACHE_L0_3_L1_2_Fij_nx262, 
         CACHE_L0_3_L1_2_Fij_nx272, CACHE_L0_3_L1_2_Fij_nx282, 
         CACHE_L0_3_L1_2_Fij_nx296, CACHE_L0_3_L1_2_Fij_nx331, 
         CACHE_L0_3_L1_2_Fij_nx333, CACHE_L0_3_L1_2_Wij_nx212, 
         CACHE_L0_3_L1_2_Wij_nx222, CACHE_L0_3_L1_2_Wij_nx232, 
         CACHE_L0_3_L1_2_Wij_nx242, CACHE_L0_3_L1_2_Wij_nx252, 
         CACHE_L0_3_L1_2_Wij_nx262, CACHE_L0_3_L1_2_Wij_nx272, 
         CACHE_L0_3_L1_2_Wij_nx282, CACHE_L0_3_L1_2_Wij_nx296, 
         CACHE_L0_3_L1_2_Wij_nx331, CACHE_L0_3_L1_2_Wij_nx333, 
         CACHE_L0_3_L1_3_Fij_nx212, CACHE_L0_3_L1_3_Fij_nx222, 
         CACHE_L0_3_L1_3_Fij_nx232, CACHE_L0_3_L1_3_Fij_nx242, 
         CACHE_L0_3_L1_3_Fij_nx252, CACHE_L0_3_L1_3_Fij_nx262, 
         CACHE_L0_3_L1_3_Fij_nx272, CACHE_L0_3_L1_3_Fij_nx282, 
         CACHE_L0_3_L1_3_Fij_nx296, CACHE_L0_3_L1_3_Fij_nx331, 
         CACHE_L0_3_L1_3_Fij_nx333, CACHE_L0_3_L1_3_Wij_nx212, 
         CACHE_L0_3_L1_3_Wij_nx222, CACHE_L0_3_L1_3_Wij_nx232, 
         CACHE_L0_3_L1_3_Wij_nx242, CACHE_L0_3_L1_3_Wij_nx252, 
         CACHE_L0_3_L1_3_Wij_nx262, CACHE_L0_3_L1_3_Wij_nx272, 
         CACHE_L0_3_L1_3_Wij_nx282, CACHE_L0_3_L1_3_Wij_nx296, 
         CACHE_L0_3_L1_3_Wij_nx331, CACHE_L0_3_L1_3_Wij_nx333, 
         CACHE_L0_3_L1_4_Fij_nx212, CACHE_L0_3_L1_4_Fij_nx222, 
         CACHE_L0_3_L1_4_Fij_nx232, CACHE_L0_3_L1_4_Fij_nx242, 
         CACHE_L0_3_L1_4_Fij_nx252, CACHE_L0_3_L1_4_Fij_nx262, 
         CACHE_L0_3_L1_4_Fij_nx272, CACHE_L0_3_L1_4_Fij_nx282, 
         CACHE_L0_3_L1_4_Fij_nx296, CACHE_L0_3_L1_4_Fij_nx331, 
         CACHE_L0_3_L1_4_Fij_nx333, CACHE_L0_3_L1_4_Wij_nx212, 
         CACHE_L0_3_L1_4_Wij_nx222, CACHE_L0_3_L1_4_Wij_nx232, 
         CACHE_L0_3_L1_4_Wij_nx242, CACHE_L0_3_L1_4_Wij_nx252, 
         CACHE_L0_3_L1_4_Wij_nx262, CACHE_L0_3_L1_4_Wij_nx272, 
         CACHE_L0_3_L1_4_Wij_nx282, CACHE_L0_3_L1_4_Wij_nx296, 
         CACHE_L0_3_L1_4_Wij_nx331, CACHE_L0_3_L1_4_Wij_nx333, 
         CACHE_L0_4_L1_0_Fij_nx212, CACHE_L0_4_L1_0_Fij_nx222, 
         CACHE_L0_4_L1_0_Fij_nx232, CACHE_L0_4_L1_0_Fij_nx242, 
         CACHE_L0_4_L1_0_Fij_nx252, CACHE_L0_4_L1_0_Fij_nx262, 
         CACHE_L0_4_L1_0_Fij_nx272, CACHE_L0_4_L1_0_Fij_nx282, 
         CACHE_L0_4_L1_0_Fij_nx296, CACHE_L0_4_L1_0_Fij_nx331, 
         CACHE_L0_4_L1_0_Fij_nx333, CACHE_L0_4_L1_0_Wij_nx212, 
         CACHE_L0_4_L1_0_Wij_nx222, CACHE_L0_4_L1_0_Wij_nx232, 
         CACHE_L0_4_L1_0_Wij_nx242, CACHE_L0_4_L1_0_Wij_nx252, 
         CACHE_L0_4_L1_0_Wij_nx262, CACHE_L0_4_L1_0_Wij_nx272, 
         CACHE_L0_4_L1_0_Wij_nx282, CACHE_L0_4_L1_0_Wij_nx296, 
         CACHE_L0_4_L1_0_Wij_nx331, CACHE_L0_4_L1_0_Wij_nx333, 
         CACHE_L0_4_L1_1_Fij_nx212, CACHE_L0_4_L1_1_Fij_nx222, 
         CACHE_L0_4_L1_1_Fij_nx232, CACHE_L0_4_L1_1_Fij_nx242, 
         CACHE_L0_4_L1_1_Fij_nx252, CACHE_L0_4_L1_1_Fij_nx262, 
         CACHE_L0_4_L1_1_Fij_nx272, CACHE_L0_4_L1_1_Fij_nx282, 
         CACHE_L0_4_L1_1_Fij_nx296, CACHE_L0_4_L1_1_Fij_nx331, 
         CACHE_L0_4_L1_1_Fij_nx333, CACHE_L0_4_L1_1_Wij_nx212, 
         CACHE_L0_4_L1_1_Wij_nx222, CACHE_L0_4_L1_1_Wij_nx232, 
         CACHE_L0_4_L1_1_Wij_nx242, CACHE_L0_4_L1_1_Wij_nx252, 
         CACHE_L0_4_L1_1_Wij_nx262, CACHE_L0_4_L1_1_Wij_nx272, 
         CACHE_L0_4_L1_1_Wij_nx282, CACHE_L0_4_L1_1_Wij_nx296, 
         CACHE_L0_4_L1_1_Wij_nx331, CACHE_L0_4_L1_1_Wij_nx333, 
         CACHE_L0_4_L1_2_Fij_nx212, CACHE_L0_4_L1_2_Fij_nx222, 
         CACHE_L0_4_L1_2_Fij_nx232, CACHE_L0_4_L1_2_Fij_nx242, 
         CACHE_L0_4_L1_2_Fij_nx252, CACHE_L0_4_L1_2_Fij_nx262, 
         CACHE_L0_4_L1_2_Fij_nx272, CACHE_L0_4_L1_2_Fij_nx282, 
         CACHE_L0_4_L1_2_Fij_nx296, CACHE_L0_4_L1_2_Fij_nx331, 
         CACHE_L0_4_L1_2_Fij_nx333, CACHE_L0_4_L1_2_Wij_nx212, 
         CACHE_L0_4_L1_2_Wij_nx222, CACHE_L0_4_L1_2_Wij_nx232, 
         CACHE_L0_4_L1_2_Wij_nx242, CACHE_L0_4_L1_2_Wij_nx252, 
         CACHE_L0_4_L1_2_Wij_nx262, CACHE_L0_4_L1_2_Wij_nx272, 
         CACHE_L0_4_L1_2_Wij_nx282, CACHE_L0_4_L1_2_Wij_nx296, 
         CACHE_L0_4_L1_2_Wij_nx331, CACHE_L0_4_L1_2_Wij_nx333, 
         CACHE_L0_4_L1_3_Fij_nx212, CACHE_L0_4_L1_3_Fij_nx222, 
         CACHE_L0_4_L1_3_Fij_nx232, CACHE_L0_4_L1_3_Fij_nx242, 
         CACHE_L0_4_L1_3_Fij_nx252, CACHE_L0_4_L1_3_Fij_nx262, 
         CACHE_L0_4_L1_3_Fij_nx272, CACHE_L0_4_L1_3_Fij_nx282, 
         CACHE_L0_4_L1_3_Fij_nx296, CACHE_L0_4_L1_3_Fij_nx331, 
         CACHE_L0_4_L1_3_Fij_nx333, CACHE_L0_4_L1_3_Wij_nx212, 
         CACHE_L0_4_L1_3_Wij_nx222, CACHE_L0_4_L1_3_Wij_nx232, 
         CACHE_L0_4_L1_3_Wij_nx242, CACHE_L0_4_L1_3_Wij_nx252, 
         CACHE_L0_4_L1_3_Wij_nx262, CACHE_L0_4_L1_3_Wij_nx272, 
         CACHE_L0_4_L1_3_Wij_nx282, CACHE_L0_4_L1_3_Wij_nx296, 
         CACHE_L0_4_L1_3_Wij_nx331, CACHE_L0_4_L1_3_Wij_nx333, 
         CACHE_L0_4_L1_4_Fij_nx212, CACHE_L0_4_L1_4_Fij_nx222, 
         CACHE_L0_4_L1_4_Fij_nx232, CACHE_L0_4_L1_4_Fij_nx242, 
         CACHE_L0_4_L1_4_Fij_nx252, CACHE_L0_4_L1_4_Fij_nx262, 
         CACHE_L0_4_L1_4_Fij_nx272, CACHE_L0_4_L1_4_Fij_nx282, 
         CACHE_L0_4_L1_4_Fij_nx296, CACHE_L0_4_L1_4_Fij_nx331, 
         CACHE_L0_4_L1_4_Fij_nx333, CACHE_L0_4_L1_4_Wij_nx212, 
         CACHE_L0_4_L1_4_Wij_nx222, CACHE_L0_4_L1_4_Wij_nx232, 
         CACHE_L0_4_L1_4_Wij_nx242, CACHE_L0_4_L1_4_Wij_nx252, 
         CACHE_L0_4_L1_4_Wij_nx262, CACHE_L0_4_L1_4_Wij_nx272, 
         CACHE_L0_4_L1_4_Wij_nx282, CACHE_L0_4_L1_4_Wij_nx296, 
         CACHE_L0_4_L1_4_Wij_nx331, CACHE_L0_4_L1_4_Wij_nx333, nx619, nx621, 
         nx623, nx625, nx627, nx629, nx631, nx633, nx635, nx637, nx639, nx641, 
         nx643, nx647, nx649, nx651, nx653, nx655, nx657, nx659, nx661, nx663, 
         nx665, nx669, nx671, nx673, nx675, nx677, nx679, nx681, nx683, nx685, 
         nx687, nx689, nx691, nx693, nx695, nx697, nx699, nx701, nx703, nx705, 
         nx707, nx709, nx711, nx713, nx715, nx717, nx719, nx721, nx723, nx725, 
         nx727, nx729, nx731, nx733, nx735, nx737, nx739, nx741, nx743, nx745, 
         nx747, nx749, nx751, nx753, nx755, nx757, nx759, nx761, nx763, nx765, 
         nx767, nx769, nx771, nx773, nx775, nx777, nx779, nx781, nx783, nx785, 
         nx787, nx789, nx791, nx793, nx795, nx797, nx799, nx801, nx803, nx805, 
         nx807, nx809, nx811, nx813, nx815, nx817, nx819, nx821, nx823, nx825, 
         nx827, nx829, nx831, nx833, nx835, nx837, nx839, nx841, nx843, nx845, 
         nx847, nx849, nx851, nx853, nx855, nx857, nx859, nx861, nx863, nx865, 
         nx867, nx871, nx873, nx875, nx877, nx879, nx881, nx883, nx885, nx887, 
         nx889, nx891, nx893, nx895, nx897, nx899, nx901, nx903, nx905, nx907, 
         nx909, nx911, nx913, nx915, nx917, nx919, nx921, nx923, nx925, nx927, 
         nx929, nx931, nx933, nx935, nx937, nx939, nx941, nx943, nx945, nx947, 
         nx949, nx951, nx953, nx955, nx957, nx959, nx961, nx963, nx965, nx967, 
         nx969, nx971, nx973, nx975, nx977, nx979, nx981, nx983, nx985, nx987, 
         nx989, nx991, nx993, nx995, nx997, nx999, nx1001, nx1003, nx1005, 
         nx1007, nx1009, nx1011, nx1013, nx1015, nx1017, nx1019, nx1021, nx1023, 
         nx1025, nx1027, nx1029, nx1031, nx1033, nx1035, nx1037, nx1039, nx1041, 
         nx1043, nx1045, nx1047, nx1049, nx1051, nx1053, nx1055, nx1057, nx1059, 
         nx1061, nx1063, nx1065, nx1067, nx1069, nx1071, nx1073, nx1075, nx1077, 
         nx1079, nx1081, nx1083, nx1085, nx1087, nx1089, nx1091, nx1093, nx1095, 
         nx1097, nx1099, nx1101, nx1103, nx1105, nx1107, nx1109, nx1111, nx1113, 
         nx1115, nx1119, nx1121, nx1123, nx1125, nx1127, nx1129, nx1131, nx1133, 
         nx1135, nx1137, nx1139, nx1141, nx1143, nx1145, nx1147, nx1149, nx1151, 
         nx1153, nx1155, nx1157, nx1159, nx1161, nx1163, nx1165, nx1167, nx1169, 
         nx1171, nx1173, nx1175, nx1177, nx1179, nx1181, nx1183, nx1185, nx1187, 
         nx1189, nx1191, nx1193, nx1195, nx1197, nx1199, nx1201, nx1203, nx1205, 
         nx1207, nx1209, nx1211, nx1213, nx1215, nx1217, nx1219, nx1221, nx1223, 
         nx1225, nx1227, nx1229, nx1231, nx1233, nx1235, nx1237, nx1239, nx1241, 
         nx1243, nx1245, nx1247, nx1249, nx1251, nx1253, nx1255, nx1257, nx1259, 
         nx1261, nx1263, nx1265, nx1267, nx1269, nx1271, nx1273, nx1275, nx1277, 
         nx1279, nx1281, nx1283, nx1285, nx1287, nx1289, nx1291, nx1293, nx1295, 
         nx1297, nx1299, nx1301, nx1303, nx1305, nx1307, nx1309, nx1311, nx1313, 
         nx1315, nx1317, nx1319, nx1321, nx1323, nx1325, nx1327, nx1329, nx1331, 
         nx1333, nx1335, nx1337, nx1339, nx1341, nx1343, nx1345, nx1347, nx1349, 
         nx1351, nx1353, nx1355, nx1357, nx1359, nx1361, nx1363, nx1367, nx1369, 
         nx1371, nx1373, nx1375, nx1377, nx1379, nx1381, nx1383, nx1385, nx1387, 
         nx1389, nx1391, nx1393, nx1395, nx1397, nx1399, nx1401, nx1403, nx1405, 
         nx1407, nx1409, nx1411, nx1413, nx1415, nx1417, nx1419, nx1421, nx1423, 
         nx1425, nx1427, nx1429, nx1431, nx1433, nx1435, nx1437, nx1439, nx1441, 
         nx1443, nx1445, nx1447, nx1449, nx1451, nx1453, nx1455, nx1457, nx1459, 
         nx1461, nx1463, nx1465, nx1467, nx1469, nx1471, nx1473, nx1475, nx1477, 
         nx1479, nx1481, nx1483, nx1485, nx1487, nx1489, nx1491, nx1493, nx1495, 
         nx1497, nx1499, nx1501, nx1503, nx1505, nx1507, nx1509, nx1511, nx1513, 
         nx1515, nx1517, nx1519, nx1521, nx1523, nx1525, nx1527, nx1529, nx1531, 
         nx1533, nx1535, nx1537, nx1539, nx1541, nx1543, nx1545, nx1547, nx1549, 
         nx1551, nx1553, nx1555, nx1557, nx1559, nx1561, nx1563, nx1565, nx1567, 
         nx1569, nx1571, nx1573, nx1575, nx1577, nx1579, nx1581, nx1583, nx1585, 
         nx1587, nx1589, nx1591, nx1593, nx1595, nx1597, nx1599, nx1601, nx1603, 
         nx1605, nx1607, nx1609, nx1611, nx1615, nx1617, nx1619, nx1621, nx1623, 
         nx1625, nx1627, nx1629, nx1631, nx1633, nx1635, nx1637, nx1639, nx1641, 
         nx1643, nx1645, nx1647, nx1649, nx1651, nx1653, nx1655, nx1657, nx1659, 
         nx1661, nx1663, nx1665, nx1667, nx1669, nx1671, nx1673, nx1675, nx1677, 
         nx1679, nx1681, nx1683, nx1685, nx1687, nx1689, nx1691, nx1693, nx1695, 
         nx1697, nx1699, nx1701, nx1703, nx1705, nx1707, nx1709, nx1711, nx1713, 
         nx1715, nx1717, nx1719, nx1721, nx1723, nx1725, nx1727, nx1729, nx1731, 
         nx1733, nx1735, nx1737, nx1739, nx1741, nx1743, nx1745, nx1747, nx1749, 
         nx1751, nx1753, nx1755, nx1757, nx1759, nx1761, nx1763, nx1765, nx1767, 
         nx1769, nx1771, nx1773, nx1775, nx1777, nx1779, nx1781, nx1783, nx1785, 
         nx1787, nx1789, nx1791, nx1793, nx1795, nx1797, nx1799, nx1801, nx1803, 
         nx1805, nx1807, nx1809, nx1811, nx1813, nx1815, nx1817, nx1819, nx1821, 
         nx1823, nx1825, nx1827, nx1829, nx1831, nx1833, nx1835, nx1837, nx1839, 
         nx1841, nx1843, nx1845, nx1847, nx1849, nx1851, nx1853, nx1855, nx1857, 
         nx1859, nx1863, nx1865, nx1867, nx1869, nx1871, nx1873, nx1875, nx1877, 
         nx1879, nx1881, nx1883, nx1885, nx1887, nx1889, nx1891, nx1893, nx1895, 
         nx1897, nx1899, nx1901, nx1903, nx1905, nx1907, nx1909, nx1911, nx1913, 
         nx1915, nx1917, nx1919, nx1921, nx1923, nx1925, nx1927, nx1929, nx1931, 
         nx1933, nx1935, nx1937, nx1939, nx1941, nx1943, nx1945, nx1947, nx1949, 
         nx1951, nx1953, nx1955, nx1957, nx1959, nx1961, nx1963, nx1965, nx1967, 
         nx1969, nx1971, nx1973, nx1975, nx1977, nx1979, nx1981, nx1983, nx1985, 
         nx1987, nx1989, nx1991, nx1993, nx1995, nx1997, nx1999, nx2001, nx2003, 
         nx2005, nx2007, nx2009, nx2011, nx2013, nx2015, nx2017, nx2019, nx2021, 
         nx2023, nx2025, nx2027, nx2029, nx2031, nx2033, nx2035, nx2037, nx2039, 
         nx2041, nx2043, nx2045, nx2047, nx2049, nx2051, nx2053, nx2055, nx2057, 
         nx2059, nx2061, nx2063, nx2065, nx2067, nx2069, nx2071, nx2073, nx2075, 
         nx2077, nx2079, nx2081, nx2083, nx2085, nx2087, nx2089, nx2091, nx2093, 
         nx2095, nx2097, nx2099, nx2101, nx2103, nx2105, nx2107, nx2111, nx2113, 
         nx2115, nx2117, nx2119, nx2121, nx2123, nx2125, nx2127, nx2129, nx2131, 
         nx2133, nx2135, nx2137, nx2139, nx2141, nx2143, nx2145, nx2147, nx2149, 
         nx2151, nx2153, nx2155, nx2157, nx2159, nx2161, nx2163, nx2165, nx2167, 
         nx2169, nx2171, nx2173, nx2175, nx2177, nx2179, nx2181, nx2183, nx2185, 
         nx2187, nx2189, nx2191, nx2193, nx2195, nx2197, nx2199, nx2201, nx2203, 
         nx2205, nx2207, nx2209, nx2211, nx2213, nx2215, nx2217, nx2219, nx2221, 
         nx2223, nx2225, nx2227, nx2229, nx2231, nx2233, nx2235, nx2237, nx2239, 
         nx2241, nx2243, nx2245, nx2247, nx2249, nx2251, nx2253, nx2255, nx2257, 
         nx2259, nx2261, nx2263, nx2265, nx2267, nx2269, nx2271, nx2273, nx2275, 
         nx2277, nx2279, nx2281, nx2283, nx2285, nx2287, nx2289, nx2291, nx2293, 
         nx2295, nx2297, nx2299, nx2301, nx2303, nx2305, nx2307, nx2309, nx2311, 
         nx2313, nx2315, nx2317, nx2319, nx2321, nx2323, nx2325, nx2327, nx2329, 
         nx2331, nx2333, nx2335, nx2337, nx2339, nx2341, nx2343, nx2345, nx2347, 
         nx2349, nx2351, nx2353, nx2355, nx2359, nx2361, nx2363, nx2365, nx2367, 
         nx2369, nx2371, nx2373, nx2375, nx2377, nx2379, nx2381, nx2383, nx2385, 
         nx2387, nx2389, nx2391, nx2393, nx2395, nx2397, nx2399, nx2401, nx2403, 
         nx2405, nx2407, nx2409, nx2411, nx2413, nx2415, nx2417, nx2419, nx2421, 
         nx2423, nx2425, nx2427, nx2429, nx2431, nx2433, nx2435, nx2437, nx2439, 
         nx2441, nx2443, nx2445, nx2447, nx2449, nx2451, nx2453, nx2455, nx2457, 
         nx2459, nx2461, nx2463, nx2465, nx2467, nx2469, nx2471, nx2473, nx2475, 
         nx2477, nx2479, nx2481, nx2483, nx2485, nx2487, nx2489, nx2491, nx2493, 
         nx2495, nx2497, nx2499, nx2501, nx2503, nx2505, nx2507, nx2509, nx2511, 
         nx2513, nx2515, nx2517, nx2519, nx2521, nx2523, nx2525, nx2527, nx2529, 
         nx2531, nx2533, nx2535, nx2537, nx2539, nx2541, nx2543, nx2545, nx2547, 
         nx2549, nx2551, nx2553, nx2555, nx2557, nx2559, nx2561, nx2563, nx2565, 
         nx2567, nx2569, nx2571, nx2573, nx2575, nx2577, nx2579, nx2581, nx2583, 
         nx2585, nx2587, nx2589, nx2591, nx2593, nx2595, nx2597, nx2599, nx2601, 
         nx2603, nx2607, nx2609, nx2611, nx2613, nx2615, nx2617, nx2619, nx2621, 
         nx2623, nx2625, nx2627, nx2629, nx2631, nx2633, nx2635, nx2637, nx2639, 
         nx2641, nx2643, nx2645, nx2647, nx2649, nx2651, nx2653, nx2655, nx2657, 
         nx2659, nx2661, nx2663, nx2665, nx2667, nx2669, nx2671, nx2673, nx2675, 
         nx2677, nx2679, nx2681, nx2683, nx2685, nx2687, nx2689, nx2691, nx2693, 
         nx2695, nx2697, nx2699, nx2701, nx2703, nx2705, nx2707, nx2709, nx2711, 
         nx2713, nx2715, nx2717, nx2719, nx2721, nx2723, nx2725, nx2727, nx2729, 
         nx2731, nx2733, nx2735, nx2737, nx2739, nx2741, nx2743, nx2745, nx2747, 
         nx2749, nx2751, nx2753, nx2755, nx2757, nx2759, nx2761, nx2763, nx2765, 
         nx2767, nx2769, nx2771, nx2773, nx2775, nx2777, nx2779, nx2781, nx2783, 
         nx2785, nx2787, nx2789, nx2791, nx2793, nx2795, nx2797, nx2799, nx2801, 
         nx2803, nx2805, nx2807, nx2809, nx2811, nx2813, nx2815, nx2817, nx2819, 
         nx2821, nx2823, nx2825, nx2827, nx2829, nx2831, nx2833, nx2835, nx2837, 
         nx2839, nx2841, nx2843, nx2845, nx2847, nx2849, nx2851, nx2855, nx2857, 
         nx2859, nx2861, nx2863, nx2865, nx2867, nx2869, nx2871, nx2873, nx2875, 
         nx2877, nx2879, nx2881, nx2883, nx2885, nx2887, nx2889, nx2891, nx2893, 
         nx2895, nx2897, nx2899, nx2901, nx2903, nx2905, nx2907, nx2909, nx2911, 
         nx2913, nx2915, nx2917, nx2919, nx2921, nx2923, nx2925, nx2927, nx2929, 
         nx2931, nx2933, nx2935, nx2937, nx2939, nx2941, nx2943, nx2945, nx2947, 
         nx2949, nx2951, nx2953, nx2955, nx2957, nx2959, nx2961, nx2963, nx2965, 
         nx2967, nx2969, nx2971, nx2973, nx2975, nx2977, nx2979, nx2981, nx2983, 
         nx2985, nx2987, nx2989, nx2991, nx2993, nx2995, nx2997, nx2999, nx3001, 
         nx3003, nx3005, nx3007, nx3009, nx3011, nx3013, nx3015, nx3017, nx3019, 
         nx3021, nx3023, nx3025, nx3027, nx3029, nx3031, nx3033, nx3035, nx3037, 
         nx3039, nx3041, nx3043, nx3045, nx3047, nx3049, nx3051, nx3053, nx3055, 
         nx3057, nx3059, nx3061, nx3063, nx3065, nx3067, nx3069, nx3071, nx3073, 
         nx3075, nx3077, nx3079, nx3081, nx3083, nx3085, nx3087, nx3089, nx3091, 
         nx3093, nx3095, nx3097, nx3099, nx3103, nx3105, nx3107, nx3109, nx3111, 
         nx3113, nx3115, nx3117, nx3119, nx3121, nx3123, nx3125, nx3127, nx3129, 
         nx3131, nx3133, nx3135, nx3137, nx3139, nx3141, nx3143, nx3145, nx3147, 
         nx3149, nx3151, nx3153, nx3155, nx3157, nx3159, nx3161, nx3163, nx3165, 
         nx3167, nx3169, nx3171, nx3173, nx3175, nx3177, nx3179, nx3181, nx3183, 
         nx3185, nx3187, nx3189, nx3191, nx3193, nx3195, nx3197, nx3199, nx3201, 
         nx3203, nx3205, nx3207, nx3209, nx3211, nx3213, nx3215, nx3217, nx3219, 
         nx3221, nx3223, nx3225, nx3227, nx3229, nx3231, nx3233, nx3235, nx3237, 
         nx3239, nx3241, nx3243, nx3245, nx3247, nx3249, nx3251, nx3253, nx3255, 
         nx3257, nx3259, nx3261, nx3263, nx3265, nx3267, nx3269, nx3271, nx3273, 
         nx3275, nx3277, nx3279, nx3281, nx3283, nx3285, nx3287, nx3289, nx3291, 
         nx3293, nx3295, nx3297, nx3299, nx3301, nx3303, nx3305, nx3307, nx3309, 
         nx3311, nx3313, nx3315, nx3317, nx3319, nx3321, nx3323, nx3325, nx3327, 
         nx3329, nx3331, nx3333, nx3335, nx3337, nx3339, nx3341, nx3343, nx3345, 
         nx3347, nx3351, nx3353, nx3355, nx3357, nx3359, nx3361, nx3363, nx3365, 
         nx3367, nx3369, nx3371, nx3373, nx3375, nx3377, nx3379, nx3381, nx3383, 
         nx3385, nx3387, nx3389, nx3391, nx3393, nx3395, nx3397, nx3399, nx3401, 
         nx3403, nx3405, nx3407, nx3409, nx3411, nx3413, nx3415, nx3417, nx3419, 
         nx3421, nx3423, nx3425, nx3427, nx3429, nx3431, nx3433, nx3435, nx3437, 
         nx3439, nx3441, nx3443, nx3445, nx3447, nx3449, nx3451, nx3453, nx3455, 
         nx3457, nx3459, nx3461, nx3463, nx3465, nx3467, nx3469, nx3471, nx3473, 
         nx3475, nx3477, nx3479, nx3481, nx3483, nx3485, nx3487, nx3489, nx3491, 
         nx3493, nx3495, nx3497, nx3499, nx3501, nx3503, nx3505, nx3507, nx3509, 
         nx3511, nx3513, nx3515, nx3517, nx3519, nx3521, nx3523, nx3525, nx3527, 
         nx3529, nx3531, nx3533, nx3535, nx3537, nx3539, nx3541, nx3543, nx3545, 
         nx3547, nx3549, nx3551, nx3553, nx3555, nx3557, nx3559, nx3561, nx3563, 
         nx3565, nx3567, nx3569, nx3571, nx3573, nx3575, nx3577, nx3579, nx3581, 
         nx3583, nx3585, nx3587, nx3589, nx3591, nx3593, nx3595, nx3599, nx3601, 
         nx3603, nx3605, nx3607, nx3609, nx3611, nx3613, nx3615, nx3617, nx3619, 
         nx3621, nx3623, nx3625, nx3627, nx3629, nx3631, nx3633, nx3635, nx3637, 
         nx3639, nx3641, nx3643, nx3645, nx3647, nx3649, nx3651, nx3653, nx3655, 
         nx3657, nx3659, nx3661, nx3663, nx3665, nx3667, nx3669, nx3671, nx3673, 
         nx3675, nx3677, nx3679, nx3681, nx3683, nx3685, nx3687, nx3689, nx3691, 
         nx3693, nx3695, nx3697, nx3699, nx3701, nx3703, nx3705, nx3707, nx3709, 
         nx3711, nx3713, nx3715, nx3717, nx3719, nx3721, nx3723, nx3725, nx3727, 
         nx3729, nx3731, nx3733, nx3735, nx3737, nx3739, nx3741, nx3743, nx3745, 
         nx3747, nx3749, nx3751, nx3753, nx3755, nx3757, nx3759, nx3761, nx3763, 
         nx3765, nx3767, nx3769, nx3771, nx3773, nx3775, nx3777, nx3779, nx3781, 
         nx3783, nx3785, nx3787, nx3789, nx3791, nx3793, nx3795, nx3797, nx3799, 
         nx3801, nx3803, nx3805, nx3807, nx3809, nx3811, nx3813, nx3815, nx3817, 
         nx3819, nx3821, nx3823, nx3825, nx3827, nx3829, nx3831, nx3833, nx3835, 
         nx3837, nx3839, nx3841, nx3843, nx3847, nx3849, nx3851, nx3853, nx3855, 
         nx3857, nx3859, nx3861, nx3863, nx3865, nx3867, nx3869, nx3871, nx3873, 
         nx3875, nx3877, nx3879, nx3881, nx3883, nx3885, nx3887, nx3889, nx3891, 
         nx3893, nx3895, nx3897, nx3899, nx3901, nx3903, nx3905, nx3907, nx3909, 
         nx3911, nx3913, nx3915, nx3917, nx3919, nx3921, nx3923, nx3925, nx3927, 
         nx3929, nx3931, nx3933, nx3935, nx3937, nx3939, nx3941, nx3943, nx3945, 
         nx3947, nx3949, nx3951, nx3953, nx3955, nx3957, nx3959, nx3961, nx3963, 
         nx3965, nx3967, nx3969, nx3971, nx3973, nx3975, nx3977, nx3979, nx3981, 
         nx3983, nx3985, nx3987, nx3989, nx3991, nx3993, nx3995, nx3997, nx3999, 
         nx4001, nx4003, nx4005, nx4007, nx4009, nx4011, nx4013, nx4015, nx4017, 
         nx4019, nx4021, nx4023, nx4025, nx4027, nx4029, nx4031, nx4033, nx4035, 
         nx4037, nx4039, nx4041, nx4043, nx4045, nx4047, nx4049, nx4051, nx4053, 
         nx4055, nx4057, nx4059, nx4061, nx4063, nx4065, nx4067, nx4069, nx4071, 
         nx4073, nx4075, nx4077, nx4079, nx4081, nx4083, nx4085, nx4087, nx4089, 
         nx4091, nx4095, nx4097, nx4099, nx4101, nx4103, nx4105, nx4107, nx4109, 
         nx4111, nx4113, nx4115, nx4117, nx4119, nx4121, nx4123, nx4125, nx4127, 
         nx4129, nx4131, nx4133, nx4135, nx4137, nx4139, nx4141, nx4143, nx4145, 
         nx4147, nx4149, nx4151, nx4153, nx4155, nx4157, nx4159, nx4161, nx4163, 
         nx4165, nx4167, nx4169, nx4171, nx4173, nx4175, nx4177, nx4179, nx4181, 
         nx4183, nx4185, nx4187, nx4189, nx4191, nx4193, nx4195, nx4197, nx4199, 
         nx4201, nx4203, nx4205, nx4207, nx4209, nx4211, nx4213, nx4215, nx4217, 
         nx4219, nx4221, nx4223, nx4225, nx4227, nx4229, nx4231, nx4233, nx4235, 
         nx4237, nx4239, nx4241, nx4243, nx4245, nx4247, nx4249, nx4251, nx4253, 
         nx4255, nx4257, nx4259, nx4261, nx4263, nx4265, nx4267, nx4269, nx4271, 
         nx4273, nx4275, nx4277, nx4279, nx4281, nx4283, nx4285, nx4287, nx4289, 
         nx4291, nx4293, nx4295, nx4297, nx4299, nx4301, nx4303, nx4305, nx4307, 
         nx4309, nx4311, nx4313, nx4315, nx4317, nx4319, nx4321, nx4323, nx4325, 
         nx4327, nx4329, nx4331, nx4333, nx4335, nx4337, nx4339, nx4343, nx4345, 
         nx4347, nx4349, nx4351, nx4353, nx4355, nx4357, nx4359, nx4361, nx4363, 
         nx4365, nx4367, nx4369, nx4371, nx4373, nx4375, nx4377, nx4379, nx4381, 
         nx4383, nx4385, nx4387, nx4389, nx4391, nx4393, nx4395, nx4397, nx4399, 
         nx4401, nx4403, nx4405, nx4407, nx4409, nx4411, nx4413, nx4415, nx4417, 
         nx4419, nx4421, nx4423, nx4425, nx4427, nx4429, nx4431, nx4433, nx4435, 
         nx4437, nx4439, nx4441, nx4443, nx4445, nx4447, nx4449, nx4451, nx4453, 
         nx4455, nx4457, nx4459, nx4461, nx4463, nx4465, nx4467, nx4469, nx4471, 
         nx4473, nx4475, nx4477, nx4479, nx4481, nx4483, nx4485, nx4487, nx4489, 
         nx4491, nx4493, nx4495, nx4497, nx4499, nx4501, nx4503, nx4505, nx4507, 
         nx4509, nx4511, nx4513, nx4515, nx4517, nx4519, nx4521, nx4523, nx4525, 
         nx4527, nx4529, nx4531, nx4533, nx4535, nx4537, nx4539, nx4541, nx4543, 
         nx4545, nx4547, nx4549, nx4551, nx4553, nx4555, nx4557, nx4559, nx4561, 
         nx4563, nx4565, nx4567, nx4569, nx4571, nx4573, nx4575, nx4577, nx4579, 
         nx4581, nx4583, nx4585, nx4587, nx4591, nx4593, nx4595, nx4597, nx4599, 
         nx4601, nx4603, nx4605, nx4607, nx4609, nx4611, nx4613, nx4615, nx4617, 
         nx4619, nx4621, nx4623, nx4625, nx4627, nx4629, nx4631, nx4633, nx4635, 
         nx4637, nx4639, nx4641, nx4643, nx4645, nx4647, nx4649, nx4651, nx4653, 
         nx4655, nx4657, nx4659, nx4661, nx4663, nx4665, nx4667, nx4669, nx4671, 
         nx4673, nx4675, nx4677, nx4679, nx4681, nx4683, nx4685, nx4687, nx4689, 
         nx4691, nx4693, nx4695, nx4697, nx4699, nx4701, nx4703, nx4705, nx4707, 
         nx4709, nx4711, nx4713, nx4715, nx4717, nx4719, nx4721, nx4723, nx4725, 
         nx4727, nx4729, nx4731, nx4733, nx4735, nx4737, nx4739, nx4741, nx4743, 
         nx4745, nx4747, nx4749, nx4751, nx4753, nx4755, nx4757, nx4759, nx4761, 
         nx4763, nx4765, nx4767, nx4769, nx4771, nx4773, nx4775, nx4777, nx4779, 
         nx4781, nx4783, nx4785, nx4787, nx4789, nx4791, nx4793, nx4795, nx4797, 
         nx4799, nx4801, nx4803, nx4805, nx4807, nx4809, nx4811, nx4813, nx4815, 
         nx4817, nx4819, nx4821, nx4823, nx4825, nx4827, nx4829, nx4831, nx4833, 
         nx4835, nx4839, nx4841, nx4843, nx4845, nx4847, nx4849, nx4851, nx4853, 
         nx4855, nx4857, nx4859, nx4861, nx4863, nx4865, nx4867, nx4869, nx4871, 
         nx4873, nx4875, nx4877, nx4879, nx4881, nx4883, nx4885, nx4887, nx4889, 
         nx4891, nx4893, nx4895, nx4897, nx4899, nx4901, nx4903, nx4905, nx4907, 
         nx4909, nx4911, nx4913, nx4915, nx4917, nx4919, nx4921, nx4923, nx4925, 
         nx4927, nx4929, nx4931, nx4933, nx4935, nx4937, nx4939, nx4941, nx4943, 
         nx4945, nx4947, nx4949, nx4951, nx4953, nx4955, nx4957, nx4959, nx4961, 
         nx4963, nx4965, nx4967, nx4969, nx4971, nx4973, nx4975, nx4977, nx4979, 
         nx4981, nx4983, nx4985, nx4987, nx4989, nx4991, nx4993, nx4995, nx4997, 
         nx4999, nx5001, nx5003, nx5005, nx5007, nx5009, nx5011, nx5013, nx5015, 
         nx5017, nx5019, nx5021, nx5023, nx5025, nx5027, nx5029, nx5031, nx5033, 
         nx5035, nx5037, nx5039, nx5041, nx5043, nx5045, nx5047, nx5049, nx5051, 
         nx5053, nx5055, nx5057, nx5059, nx5061, nx5063, nx5065, nx5067, nx5069, 
         nx5071, nx5073, nx5075, nx5077, nx5079, nx5081, nx5083, nx5087, nx5089, 
         nx5091, nx5093, nx5095, nx5097, nx5099, nx5101, nx5103, nx5105, nx5107, 
         nx5109, nx5111, nx5113, nx5115, nx5117, nx5119, nx5121, nx5123, nx5125, 
         nx5127, nx5129, nx5131, nx5133, nx5135, nx5137, nx5139, nx5141, nx5143, 
         nx5145, nx5147, nx5149, nx5151, nx5153, nx5155, nx5157, nx5159, nx5161, 
         nx5163, nx5165, nx5167, nx5169, nx5171, nx5173, nx5175, nx5177, nx5179, 
         nx5181, nx5183, nx5185, nx5187, nx5189, nx5191, nx5193, nx5195, nx5197, 
         nx5199, nx5201, nx5203, nx5205, nx5207, nx5209, nx5211, nx5213, nx5215, 
         nx5217, nx5219, nx5221, nx5223, nx5225, nx5227, nx5229, nx5231, nx5233, 
         nx5235, nx5237, nx5239, nx5241, nx5243, nx5245, nx5247, nx5249, nx5251, 
         nx5253, nx5255, nx5257, nx5259, nx5261, nx5263, nx5265, nx5267, nx5269, 
         nx5271, nx5273, nx5275, nx5277, nx5279, nx5281, nx5283, nx5285, nx5287, 
         nx5289, nx5291, nx5293, nx5295, nx5297, nx5299, nx5301, nx5303, nx5305, 
         nx5307, nx5309, nx5311, nx5313, nx5315, nx5317, nx5319, nx5321, nx5323, 
         nx5325, nx5327, nx5329, nx5331, nx5335, nx5337, nx5339, nx5341, nx5343, 
         nx5345, nx5347, nx5349, nx5351, nx5353, nx5355, nx5357, nx5359, nx5361, 
         nx5363, nx5365, nx5367, nx5369, nx5371, nx5373, nx5375, nx5377, nx5379, 
         nx5381, nx5383, nx5385, nx5387, nx5389, nx5391, nx5393, nx5395, nx5397, 
         nx5399, nx5401, nx5403, nx5405, nx5407, nx5409, nx5411, nx5413, nx5415, 
         nx5417, nx5419, nx5421, nx5423, nx5425, nx5427, nx5429, nx5431, nx5433, 
         nx5435, nx5437, nx5439, nx5441, nx5443, nx5445, nx5447, nx5449, nx5451, 
         nx5453, nx5455, nx5457, nx5459, nx5461, nx5463, nx5465, nx5467, nx5469, 
         nx5471, nx5473, nx5475, nx5477, nx5479, nx5481, nx5483, nx5485, nx5487, 
         nx5489, nx5491, nx5493, nx5495, nx5497, nx5499, nx5501, nx5503, nx5505, 
         nx5507, nx5509, nx5511, nx5513, nx5515, nx5517, nx5519, nx5521, nx5523, 
         nx5525, nx5527, nx5529, nx5531, nx5533, nx5535, nx5537, nx5539, nx5541, 
         nx5543, nx5545, nx5547, nx5549, nx5551, nx5553, nx5555, nx5557, nx5559, 
         nx5561, nx5563, nx5565, nx5567, nx5569, nx5571, nx5573, nx5575, nx5577, 
         nx5579, nx5583, nx5585, nx5587, nx5589, nx5591, nx5593, nx5595, nx5597, 
         nx5599, nx5601, nx5603, nx5605, nx5607, nx5609, nx5611, nx5613, nx5615, 
         nx5617, nx5619, nx5621, nx5623, nx5625, nx5627, nx5629, nx5631, nx5633, 
         nx5635, nx5637, nx5639, nx5641, nx5643, nx5645, nx5647, nx5649, nx5651, 
         nx5653, nx5655, nx5657, nx5659, nx5661, nx5663, nx5665, nx5667, nx5669, 
         nx5671, nx5673, nx5675, nx5677, nx5679, nx5681, nx5683, nx5685, nx5687, 
         nx5689, nx5691, nx5693, nx5695, nx5697, nx5699, nx5701, nx5703, nx5705, 
         nx5707, nx5709, nx5711, nx5713, nx5715, nx5717, nx5719, nx5721, nx5723, 
         nx5725, nx5727, nx5729, nx5731, nx5733, nx5735, nx5737, nx5739, nx5741, 
         nx5743, nx5745, nx5747, nx5749, nx5751, nx5753, nx5755, nx5757, nx5759, 
         nx5761, nx5763, nx5765, nx5767, nx5769, nx5771, nx5773, nx5775, nx5777, 
         nx5779, nx5781, nx5783, nx5785, nx5787, nx5789, nx5791, nx5793, nx5795, 
         nx5797, nx5799, nx5801, nx5803, nx5805, nx5807, nx5809, nx5811, nx5813, 
         nx5815, nx5817, nx5819, nx5821, nx5823, nx5825, nx5827, nx5831, nx5833, 
         nx5835, nx5837, nx5839, nx5841, nx5843, nx5845, nx5847, nx5849, nx5851, 
         nx5853, nx5855, nx5857, nx5859, nx5861, nx5863, nx5865, nx5867, nx5869, 
         nx5871, nx5873, nx5875, nx5877, nx5879, nx5881, nx5883, nx5885, nx5887, 
         nx5889, nx5891, nx5893, nx5895, nx5897, nx5899, nx5901, nx5903, nx5905, 
         nx5907, nx5909, nx5911, nx5913, nx5915, nx5917, nx5919, nx5921, nx5923, 
         nx5925, nx5927, nx5929, nx5931, nx5933, nx5935, nx5937, nx5939, nx5941, 
         nx5943, nx5945, nx5947, nx5949, nx5951, nx5953, nx5955, nx5957, nx5959, 
         nx5961, nx5963, nx5965, nx5967, nx5969, nx5971, nx5973, nx5975, nx5977, 
         nx5979, nx5981, nx5983, nx5985, nx5987, nx5989, nx5991, nx5993, nx5995, 
         nx5997, nx5999, nx6001, nx6003, nx6005, nx6007, nx6009, nx6011, nx6013, 
         nx6015, nx6017, nx6019, nx6021, nx6023, nx6025, nx6027, nx6029, nx6031, 
         nx6033, nx6035, nx6037, nx6039, nx6041, nx6043, nx6045, nx6047, nx6049, 
         nx6051, nx6053, nx6055, nx6057, nx6059, nx6061, nx6063, nx6065, nx6067, 
         nx6069, nx6071, nx6073, nx6075, nx6079, nx6081, nx6083, nx6085, nx6087, 
         nx6089, nx6091, nx6093, nx6095, nx6097, nx6099, nx6101, nx6103, nx6105, 
         nx6107, nx6109, nx6111, nx6113, nx6115, nx6117, nx6119, nx6121, nx6123, 
         nx6125, nx6127, nx6129, nx6131, nx6133, nx6135, nx6137, nx6139, nx6141, 
         nx6143, nx6145, nx6147, nx6149, nx6151, nx6153, nx6155, nx6157, nx6159, 
         nx6161, nx6163, nx6165, nx6167, nx6169, nx6171, nx6173, nx6175, nx6177, 
         nx6179, nx6181, nx6183, nx6185, nx6187, nx6189, nx6191, nx6193, nx6195, 
         nx6197, nx6199, nx6201, nx6203, nx6205, nx6207, nx6209, nx6211, nx6213, 
         nx6215, nx6217, nx6219, nx6221, nx6223, nx6225, nx6227, nx6229, nx6231, 
         nx6233, nx6235, nx6237, nx6239, nx6241, nx6243, nx6245, nx6247, nx6249, 
         nx6251, nx6253, nx6255, nx6257, nx6259, nx6261, nx6263, nx6265, nx6267, 
         nx6269, nx6271, nx6273, nx6275, nx6277, nx6279, nx6281, nx6283, nx6285, 
         nx6287, nx6289, nx6291, nx6293, nx6295, nx6297, nx6299, nx6301, nx6303, 
         nx6305, nx6307, nx6309, nx6311, nx6313, nx6315, nx6317, nx6319, nx6321, 
         nx6323, nx6327, nx6329, nx6331, nx6333, nx6335, nx6337, nx6339, nx6341, 
         nx6343, nx6345, nx6347, nx6349, nx6351, nx6353, nx6355, nx6357, nx6359, 
         nx6361, nx6363, nx6365, nx6367, nx6369, nx6371, nx6373, nx6375, nx6377, 
         nx6379, nx6381, nx6383, nx6385, nx6387, nx6389, nx6391, nx6393, nx6395, 
         nx6397, nx6399, nx6401, nx6403, nx6405, nx6407, nx6409, nx6411, nx6413, 
         nx6415, nx6417, nx6419, nx6421, nx6423, nx6425, nx6427, nx6429, nx6431, 
         nx6433, nx6435, nx6437, nx6439, nx6441, nx6443, nx6445, nx6447, nx6449, 
         nx6451, nx6453, nx6455, nx6457, nx6459, nx6461, nx6463, nx6465, nx6467, 
         nx6469, nx6471, nx6473, nx6475, nx6477, nx6479, nx6481, nx6483, nx6485, 
         nx6487, nx6489, nx6491, nx6493, nx6495, nx6497, nx6499, nx6501, nx6503, 
         nx6505, nx6507, nx6509, nx6511, nx6513, nx6515, nx6517, nx6519, nx6521, 
         nx6523, nx6525, nx6527, nx6529, nx6531, nx6533, nx6535, nx6537, nx6539, 
         nx6541, nx6543, nx6545, nx6547, nx6549, nx6551, nx6553, nx6555, nx6557, 
         nx6559, nx6561, nx6563, nx6565, nx6567, nx6569, nx6571, nx6575, nx6577, 
         nx6579, nx6581, nx6583, nx6585, nx6587, nx6589, nx6591, nx6593, nx6595, 
         nx6597, nx6599, nx6601, nx6603, nx6605, nx6607, nx6609, nx6611, nx6613, 
         nx6615, nx6617, nx6619, nx6621, nx6623, nx6625, nx6627, nx6629, nx6631, 
         nx6633, nx6635, nx6637, nx6639, nx6641, nx6643, nx6645, nx6647, nx6649, 
         nx6651, nx6653, nx6655, nx6657, nx6659, nx6661, nx6663, nx6665, nx6667, 
         nx6669, nx6671, nx6673, nx6675, nx6677, nx6679, nx6681, nx6683, nx6685, 
         nx6687, nx6689, nx6691, nx6693, nx6695, nx6697, nx6699, nx6701, nx6703, 
         nx6705, nx6707, nx6709, nx6711, nx6713, nx6715, nx6717, nx6719, nx6721, 
         nx6723, nx6725, nx6727, nx6729, nx6731, nx6733, nx6735, nx6737, nx6739, 
         nx6741, nx6743, nx6745, nx6747, nx6749, nx6751, nx6753, nx6755, nx6757, 
         nx6759, nx6761, nx6763, nx6765, nx6767, nx6769, nx6771, nx6773, nx6775, 
         nx6777, nx6779, nx6781, nx6783, nx6785, nx6787, nx6789, nx6791, nx6793, 
         nx6795, nx6797, nx6799, nx6801, nx6803, nx6805, nx6807, nx6809, nx6811, 
         nx6813, nx6815, nx6817, nx6819, nx6823, nx6825, nx6827, nx6829, nx6831, 
         nx6833, nx6835, nx6837, nx6839, nx6841, nx6843, nx6845, nx6847, nx6849, 
         nx6851, nx6853, nx6855, nx6857, nx6859, nx6861, nx6863, nx6865, nx6867, 
         nx6869, nx6871, nx6873, nx6875, nx6877, nx6879, nx6881, nx6883, nx6885, 
         nx6887, nx6889, nx6891, nx6893, nx6895, nx6897, nx6899, nx6901, nx6903, 
         nx6905, nx6909, nx6911, nx6915, nx6917, nx6921, nx6923, nx6927, nx6929, 
         nx6933, nx6935, nx6939, nx6941, nx6945, nx6947, nx6951, nx6953, nx6957, 
         nx6959, nx6963, nx6965, nx6969, nx6971, nx6975, nx6977, nx6981, nx6983, 
         nx6987, nx6989, nx6993, nx6995, nx6999, nx7001, nx7005, nx7007, nx7011, 
         nx7013, nx7017, nx7019, nx7023, nx7025, nx7029, nx7031, nx7035, nx7037, 
         nx7041, nx7043, nx7047, nx7049, nx7053, nx7055, nx7059, nx7061, nx7065, 
         nx7067, nx7071, nx7073, nx7077, nx7079, nx7083, nx7085, nx7089, nx7091, 
         nx7095, nx7097, nx7101, nx7103, nx7107, nx7109, nx7113, nx7115, nx7119, 
         nx7121, nx7125, nx7127, nx7131, nx7133, nx7137, nx7139, nx7143, nx7145, 
         nx7147, nx7151, nx7153, nx7155, nx7157, nx7159, nx7161, nx7163, nx7165, 
         nx7167, nx7171, nx7173, nx7175, nx7179, nx7181, nx7183, nx7185, nx7187, 
         nx7189, nx7191, nx7193, nx7195, nx7199, nx7201, nx7203, nx7207, nx7209, 
         nx7211, nx7213, nx7215, nx7217, nx7219, nx7221, nx7223, nx7227, nx7229, 
         nx7231, nx7235, nx7237, nx7239, nx7241, nx7243, nx7245, nx7247, nx7249, 
         nx7251, nx7255, nx7257, nx7259, nx7263, nx7265, nx7267, nx7269, nx7271, 
         nx7273, nx7275, nx7277, nx7279, nx7283, nx7285, nx7287, nx7289, nx7291, 
         nx7293, nx7295, nx7297, nx7299, nx7301, nx7303, nx7305, nx7307, nx7309, 
         nx7311, nx7313, nx7315, nx7317, nx7319, nx7321, nx7323, nx7325, nx7327, 
         nx7329, nx7331, nx7333, nx7335, nx7337, nx7339, nx7341, nx7343, nx7345, 
         nx7347, nx7349, nx7351, nx7353, nx7355, nx7357, nx7359, nx7361, nx7363, 
         nx7365, nx7367, nx7369, nx7371, nx7373, nx7375, nx7377, nx7379, nx7381, 
         nx7383, nx7385, nx7387, nx7389, nx7391, nx7393, nx7395, nx7397, nx7399, 
         nx7401, nx7403, nx7405, nx7407, nx7409, nx7411, nx7413, nx7415, nx7417, 
         nx7419, nx7421, nx7423, nx7425, nx7427, nx7429, nx7431, nx7433, nx7435, 
         nx7437, nx7439, nx7441, nx7443, nx7445, nx7447, nx7449, nx7451, nx7453, 
         nx7455, nx7457, nx7459, nx7461, nx7463, nx7465, nx7467, nx7469, nx7471, 
         nx7473, nx7475, nx7477, nx7479, nx7481, nx7483, nx7485, nx7487, nx7489, 
         nx7491, nx7493, nx7495, nx7497, nx7499, nx7501, nx7503, nx7505, nx7507, 
         nx7509, nx7511, nx7513, nx7515, nx7517, nx7519, nx7521, nx7523, nx7525, 
         nx7527, nx7529, nx7531, nx7533, nx7535, nx7537, nx7539, nx7541, nx7543, 
         nx7545, nx7547, nx7549, nx7551, nx7553, nx7555, nx7557, nx7559, nx7561, 
         nx7563, nx7565, nx7567, nx7569, nx7571, nx7573, nx7575, nx7577, nx7579, 
         nx7581, nx7583, nx7585, nx7587, nx7589, nx7591, nx7593, nx7595, nx7597, 
         nx7599, nx7601, nx7603, nx7605, nx7607, nx7609, nx7611, nx7613, nx7615, 
         nx7617, nx7619, nx7621, nx7623, nx7625, nx7627, nx7629, nx7631, nx7633, 
         nx7635, nx7637, nx7639, nx7641, nx7643, nx7645, nx7647, nx7649, nx7651, 
         nx7653, nx7655, nx7657, nx7659, nx7661, nx7663, nx7665, nx7667, nx7669, 
         nx7671, nx7673, nx7675, nx7677, nx7679, nx7681, nx7683, nx7685, nx7687, 
         nx7689, nx7691, nx7693, nx7695, nx7697, nx7699, nx7701, nx7703, nx7705, 
         nx7707, nx7709, nx7711, nx7713, nx7715, nx7717, nx7719, nx7721, nx7723, 
         nx7725, nx7727, nx7729, nx7731, nx7733, nx7735, nx7737, nx7739, nx7741, 
         nx7743, nx7745, nx7747, nx7749, nx7751, nx7753, nx7755, nx7757, nx7759, 
         nx7761, nx7763, nx7765, nx7767, nx7769, nx7771, nx7773, nx7775, nx7777, 
         nx7779, nx7781, nx7783, nx7785, nx7787, nx7789, nx7791, nx7793, nx7795, 
         nx7797, nx7799, nx7801, nx7803, nx7805, nx7807, nx7809, nx7811, nx7813, 
         nx7815, nx7817, nx7819, nx7821, nx7823, nx7825, nx7827, nx7829, nx7831, 
         nx7833, nx7835, nx7837, nx7839, nx7841, nx7843, nx7845, nx7847, nx7849, 
         nx7851, nx7853, nx7855, nx7857, nx7859, nx7861, nx7863, nx7865, nx7867, 
         nx7869, nx7871, nx7873, nx7875, nx7877, nx7879, nx7881, nx7883, nx7885, 
         nx7887, nx7889, nx7891, nx7893, nx7895, nx7897, nx7899, nx7901, nx7903, 
         nx7905, nx7907, nx7909, nx7911, nx7913, nx7915, nx7917, nx7919, nx7921, 
         nx7923, nx7925, nx7927, nx7929, nx7931, nx7933, nx7935, nx7937, nx7939, 
         nx7941, nx7943, nx7945, nx7947, nx7949, nx7951, nx7953, nx7955, nx7957, 
         nx7959, nx7961, nx7963, nx7965, nx7967, nx7969, nx7971, nx7973, nx7975, 
         nx7977, nx7979, nx7981, nx7983, nx7985, nx7987, nx7989, nx7991, nx7993, 
         nx7995, nx7997, nx7999, nx8001, nx8003, nx8005, nx8007, nx8009, nx8011, 
         nx8013, nx8015, nx8017, nx8019, nx8021, nx8023, nx8025, nx8027, nx8029, 
         nx8031, nx8033, nx8035, nx8037, nx8039, nx8041, nx8043, nx8045, nx8047, 
         nx8049, nx8051, nx8053, nx8055, nx8057, nx8059, nx8061, nx8063, nx8065, 
         nx8067, nx8069, nx8071, nx8073, nx8075, nx8077, nx8079, nx8081, nx8083, 
         nx8085, nx8087, nx8089, nx8091, nx8093, nx8095, nx8097, nx8099, nx8101, 
         nx8103, nx8105, nx8107, nx8109, nx8111, nx8113, nx8115, nx8117, nx8119, 
         nx8121, nx8123, nx8125, nx8127, nx8129, nx8131, nx8133, nx8135, nx8137, 
         nx8139, nx8141, nx8143, nx8145, nx8147, nx8149, nx8151, nx8153, nx8155, 
         nx8157, nx8159, nx8161, nx8163, nx8165, nx8167, nx8169, nx8171, nx8173, 
         nx8175, nx8177, nx8179, nx8181, nx8183, nx8185, nx8187, nx8189, nx8191, 
         nx8193, nx8195, nx8197, nx8199, nx8201, nx8203, nx8205, nx8207, nx8209, 
         nx8211, nx8213, nx8215, nx8217, nx8219, nx8221, nx8223, nx8225, nx8227, 
         nx8229, nx8231, nx8233, nx8235, nx8237, nx8239, nx8241, nx8243, nx8245, 
         nx8247, nx8249, nx8251, nx8253, nx8255, nx8257, nx8259, nx8261, nx8263, 
         nx8265, nx8267, nx8269, nx8271, nx8273, nx8275, nx8277, nx8279, nx8281, 
         nx8283, nx8285, nx8287, nx8289, nx8291, nx8293, nx8295, nx8297, nx8299, 
         nx8301, nx8303, nx8305, nx8307, nx8309, nx8311, nx8313, nx8315, nx8317, 
         nx8319, nx8321, nx8323, nx8325, nx8327, nx8329, nx8331, nx8333, nx8335, 
         nx8337, nx8339, nx8341, nx8343, nx8345, nx8347, nx8349, nx8351, nx8353, 
         nx8355, nx8357, nx8359, nx8361, nx8363, nx8365, nx8367, nx8369, nx8371, 
         nx8373, nx8375, nx8377, nx8379, nx8381, nx8383, nx8385, nx8387, nx8389, 
         nx8391, nx8393, nx8395, nx8397, nx8399, nx8401, nx8403, nx8405, nx8407, 
         nx8409, nx8411, nx8413, nx8415, nx8417, nx8419, nx8421, nx8423, nx8425, 
         nx8427, nx8429, nx8431, nx8433, nx8435, nx8437, nx8439, nx8441, nx8443, 
         nx8445, nx8447, nx8449, nx8451, nx8453, nx8455, nx8457, nx8459, nx8461, 
         nx8463, nx8465, nx8467, nx8469, nx8471, nx8473, nx8475, nx8477, nx8479, 
         nx8481, nx8483, nx8485, nx8487, nx8489, nx8491, nx8493, nx8495, nx8497, 
         nx8499, nx8501, nx8503, nx8505, nx8507, nx8509, nx8511, nx8513, nx8515, 
         nx8517, nx8519, nx8521, nx8523, nx8525, nx8527, nx8529, nx8531, nx8533, 
         nx8535, nx8537, nx8539, nx8541, nx8543, nx8545, nx8547, nx8549, nx8551, 
         nx8553, nx8555, nx8557, nx8559, nx8561, nx8563, nx8565, nx8567, nx8569, 
         nx8571, nx8573, nx8575, nx8577, nx8579, nx8581, nx8583, nx8585, nx8587, 
         nx8589, nx8591, nx8593, nx8595, nx8597, nx8599, nx8601, nx8603, nx8605, 
         nx8607, nx8609, nx8611, nx8613, nx8615, nx8617, nx8619, nx8621, nx8623, 
         nx8625, nx8627, nx8629, nx8631, nx8633, nx8635, nx8637, nx8639, nx8641, 
         nx8643, nx8645, nx8647, nx8649, nx8651, nx8653, nx8655, nx8657, nx8659, 
         nx8661, nx8663, nx8665, nx8667, nx8669, nx8671, nx8673, nx8675, nx8677, 
         nx8679, nx8681, nx8683, nx8685, nx8687, nx8689, nx8691, nx8693, nx8695, 
         nx8697, nx8699, nx8701, nx8703, nx8705, nx8707, nx8709, nx8711, nx8713, 
         nx8715, nx8717, nx8719, nx8721, nx8723, nx8725, nx8727, nx8729, nx8731, 
         nx8733, nx8735, nx8737, nx8739, nx8741, nx8743, nx8745, nx8747, nx8749, 
         nx8751, nx8753, nx8755, nx8757, nx8759, nx8761, nx8763, nx8765, nx8767, 
         nx8769, nx8771, nx8773, nx8775, nx8777, nx8779, nx8781, nx8783, nx8785, 
         nx8787, nx8789, nx8791, nx8793, nx8795, nx8797, nx8799, nx8801, nx8803, 
         nx8805, nx8807, nx8809, nx8811, nx8813, nx8815, nx8817, nx8819, nx8821, 
         nx8823, nx8825, nx8827, nx8833, nx8835, nx8837, nx8839, nx8841;
    wire [1701:0] \$dummy ;




    assign MemAddr[16] = MemWR ;
    fake_vcc ix502 (.Y (PWR)) ;
    or02 ix3 (.Y (CalcStartRST), .A0 (RST), .A1 (CalcStarted)) ;
    or02 ix1 (.Y (CacheRST), .A0 (RST), .A1 (FirstCycle)) ;
    fake_vcc CONTROLLER_ix522 (.Y (CONTROLLER_FilterAddr_17)) ;
    nor04_2x CONTROLLER_ix529 (.Y (CONTROLLER_NxtState_4), .A0 (CONTROLLER_nx561
             ), .A1 (CONTROLLER_nx563), .A2 (CONTROLLER_nx565), .A3 (
             CONTROLLER_nx567)) ;
    nand04 CONTROLLER_ix562 (.Y (CONTROLLER_nx561), .A0 (CONTROLLER_CurCol_2), .A1 (
           CONTROLLER_CurCol_3), .A2 (CONTROLLER_CurCol_4), .A3 (
           CONTROLLER_CurCol_5)) ;
    nor02_2x CONTROLLER_ix564 (.Y (CONTROLLER_nx563), .A0 (CONTROLLER_CurCol_1)
             , .A1 (FilterSize)) ;
    inv01 CONTROLLER_ix566 (.Y (CONTROLLER_nx565), .A (CONTROLLER_CurCol_6)) ;
    inv01 CONTROLLER_ix568 (.Y (CONTROLLER_nx567), .A (CONTROLLER_CurCol_7)) ;
    nor02_2x CONTROLLER_ix207 (.Y (MemAddr[17]), .A0 (CONTROLLER_nx795), .A1 (
             CONTROLLER_nx791)) ;
    xor2 CONTROLLER_ix121 (.Y (CONTROLLER_NxtCol_0), .A0 (CONTROLLER_nx571), .A1 (
         CONTROLLER_nx585)) ;
    nand02 CONTROLLER_ix572 (.Y (CONTROLLER_nx571), .A0 (CONTROLLER_CurRow_7), .A1 (
           CONTROLLER_nx12)) ;
    inv02 CONTROLLER_ix576 (.Y (CONTROLLER_nx575), .A (CONTROLLER_CurRow_6)) ;
    nand02 CONTROLLER_ix578 (.Y (CONTROLLER_nx577), .A0 (CONTROLLER_CurRow_5), .A1 (
           CONTROLLER_nx8)) ;
    inv01 CONTROLLER_ix582 (.Y (CONTROLLER_nx581), .A (CONTROLLER_CurRow_4)) ;
    nand04 CONTROLLER_ix584 (.Y (CONTROLLER_nx583), .A0 (CONTROLLER_CurRow_3), .A1 (
           CONTROLLER_CurRow_2), .A2 (CONTROLLER_nx799), .A3 (CONTROLLER_nx803)
           ) ;
    xnor2 CONTROLLER_ix586 (.Y (CONTROLLER_nx585), .A0 (CONTROLLER_CurCol_0), .A1 (
          CONTROLLER_nx58)) ;
    xnor2 CONTROLLER_ix119 (.Y (CONTROLLER_NxtCol_1), .A0 (CONTROLLER_CurCol_1)
          , .A1 (CONTROLLER_nx593)) ;
    oai21 CONTROLLER_ix594 (.Y (CONTROLLER_nx593), .A0 (CONTROLLER_CurCol_0), .A1 (
          Stride), .B0 (CONTROLLER_nx14)) ;
    xor2 CONTROLLER_ix113 (.Y (CONTROLLER_NxtCol_2), .A0 (CONTROLLER_CurCol_2), 
         .A1 (CONTROLLER_nx70)) ;
    inv01 CONTROLLER_ix600 (.Y (CONTROLLER_nx599), .A (CONTROLLER_CurCol_1)) ;
    xnor2 CONTROLLER_ix107 (.Y (CONTROLLER_NxtCol_3), .A0 (CONTROLLER_CurCol_3)
          , .A1 (CONTROLLER_nx602)) ;
    nand02 CONTROLLER_ix603 (.Y (CONTROLLER_nx602), .A0 (CONTROLLER_CurCol_2), .A1 (
           CONTROLLER_nx70)) ;
    xor2 CONTROLLER_ix101 (.Y (CONTROLLER_NxtCol_4), .A0 (CONTROLLER_CurCol_4), 
         .A1 (CONTROLLER_nx74)) ;
    inv01 CONTROLLER_ix607 (.Y (CONTROLLER_nx606), .A (CONTROLLER_CurCol_3)) ;
    xnor2 CONTROLLER_ix95 (.Y (CONTROLLER_NxtCol_5), .A0 (CONTROLLER_CurCol_5), 
          .A1 (CONTROLLER_nx609)) ;
    nand02 CONTROLLER_ix610 (.Y (CONTROLLER_nx609), .A0 (CONTROLLER_CurCol_4), .A1 (
           CONTROLLER_nx74)) ;
    xor2 CONTROLLER_ix89 (.Y (CONTROLLER_NxtCol_6), .A0 (CONTROLLER_CurCol_6), .A1 (
         CONTROLLER_nx78)) ;
    inv01 CONTROLLER_ix614 (.Y (CONTROLLER_nx613), .A (CONTROLLER_CurCol_5)) ;
    xnor2 CONTROLLER_ix83 (.Y (CONTROLLER_NxtCol_7), .A0 (CONTROLLER_nx616), .A1 (
          CONTROLLER_CurCol_7)) ;
    nand02 CONTROLLER_ix617 (.Y (CONTROLLER_nx616), .A0 (CONTROLLER_CurCol_6), .A1 (
           CONTROLLER_nx78)) ;
    inv01 CONTROLLER_ix619 (.Y (CONTROLLER_NxtRow_0), .A (CONTROLLER_CurRow_0)
          ) ;
    xnor2 CONTROLLER_ix51 (.Y (CONTROLLER_NxtRow_2), .A0 (CONTROLLER_CurRow_2), 
          .A1 (CONTROLLER_nx622)) ;
    xnor2 CONTROLLER_ix45 (.Y (CONTROLLER_NxtRow_3), .A0 (CONTROLLER_CurRow_3), 
          .A1 (CONTROLLER_nx625)) ;
    nand03 CONTROLLER_ix626 (.Y (CONTROLLER_nx625), .A0 (CONTROLLER_CurRow_2), .A1 (
           CONTROLLER_nx799), .A2 (CONTROLLER_nx803)) ;
    aoi21 CONTROLLER_ix39 (.Y (CONTROLLER_NxtRow_4), .A0 (CONTROLLER_nx583), .A1 (
          CONTROLLER_nx581), .B0 (CONTROLLER_nx8)) ;
    xor2 CONTROLLER_ix33 (.Y (CONTROLLER_NxtRow_5), .A0 (CONTROLLER_CurRow_5), .A1 (
         CONTROLLER_nx8)) ;
    aoi21 CONTROLLER_ix27 (.Y (CONTROLLER_NxtRow_6), .A0 (CONTROLLER_nx577), .A1 (
          CONTROLLER_nx575), .B0 (CONTROLLER_nx12)) ;
    xor2 CONTROLLER_ix21 (.Y (CONTROLLER_NxtRow_7), .A0 (CONTROLLER_CurRow_7), .A1 (
         CONTROLLER_nx12)) ;
    nand04 CONTROLLER_ix635 (.Y (CONTROLLER_nx634), .A0 (CONTROLLER_nx468), .A1 (
           CONTROLLER_nx482), .A2 (CONTROLLER_nx575), .A3 (CONTROLLER_nx640)) ;
    nor03_2x CONTROLLER_ix469 (.Y (CONTROLLER_nx468), .A0 (CONTROLLER_CurRow_5)
             , .A1 (CONTROLLER_CurRow_3), .A2 (CONTROLLER_CurRow_4)) ;
    aoi21 CONTROLLER_ix483 (.Y (CONTROLLER_nx482), .A0 (CONTROLLER_nx638), .A1 (
          CONTROLLER_nx799), .B0 (CONTROLLER_CurRow_2)) ;
    inv01 CONTROLLER_ix639 (.Y (CONTROLLER_nx638), .A (FilterSize)) ;
    inv01 CONTROLLER_ix641 (.Y (CONTROLLER_nx640), .A (CONTROLLER_CurRow_7)) ;
    or02 CONTROLLER_ix505 (.Y (MemRD), .A0 (CacheFilterWR), .A1 (
         CONTROLLER_nx795)) ;
    ao21 CONTROLLER_ix565 (.Y (CONTROLLER_CntRST), .A0 (CacheFilterWR), .A1 (
         CONTROLLER_NxtState_1), .B0 (nx7285)) ;
    aoi21 CONTROLLER_ix561 (.Y (CONTROLLER_NxtState_1), .A0 (CONTROLLER_nx645), 
          .A1 (CONTROLLER_nx647), .B0 (CONTROLLER_NxtState_4)) ;
    aoi21 CONTROLLER_ix646 (.Y (CONTROLLER_nx645), .A0 (CacheFilterWR), .A1 (
          CONTROLLER_nx634), .B0 (CONTROLLER_nx791)) ;
    aoi22 CONTROLLER_ix648 (.Y (CONTROLLER_nx647), .A0 (Instr), .A1 (FirstCycle)
          , .B0 (CONTROLLER_nx795), .B1 (CONTROLLER_nx632)) ;
    nor04 CONTROLLER_ix541 (.Y (FirstCycle), .A0 (CONTROLLER_nx650), .A1 (
          Calculating), .A2 (CONTROLLER_nx791), .A3 (MemRD)) ;
    inv01 CONTROLLER_ix651 (.Y (CONTROLLER_nx650), .A (Start)) ;
    ao21 CONTROLLER_ix515 (.Y (CONTROLLER_Restart), .A0 (Done), .A1 (Start), .B0 (
         RST)) ;
    nor02_2x CONTROLLER_ix595 (.Y (CONTROLLER_NxtState_0), .A0 (
             CONTROLLER_NxtState_4), .A1 (CONTROLLER_nx654)) ;
    aoi22 CONTROLLER_ix655 (.Y (CONTROLLER_nx654), .A0 (CONTROLLER_nx656), .A1 (
          FirstCycle), .B0 (CacheFilterWR), .B1 (CONTROLLER_nx492)) ;
    inv01 CONTROLLER_ix657 (.Y (CONTROLLER_nx656), .A (Instr)) ;
    nor02_2x CONTROLLER_ix571 (.Y (CONTROLLER_NxtState_2), .A0 (
             CONTROLLER_NxtState_4), .A1 (CONTROLLER_nx662)) ;
    nand02 CONTROLLER_ix663 (.Y (CONTROLLER_nx662), .A0 (Calculating), .A1 (
           AccFinishCalc)) ;
    nor02_2x CONTROLLER_ix583 (.Y (CONTROLLER_NxtState_3), .A0 (
             CONTROLLER_NxtState_4), .A1 (CONTROLLER_nx665)) ;
    aoi22 CONTROLLER_ix666 (.Y (CONTROLLER_nx665), .A0 (Calculating), .A1 (
          CONTROLLER_nx667), .B0 (CONTROLLER_nx795), .B1 (CONTROLLER_nx502)) ;
    inv01 CONTROLLER_ix668 (.Y (CONTROLLER_nx667), .A (AccFinishCalc)) ;
    aoi21 CONTROLLER_ix503 (.Y (CONTROLLER_nx502), .A0 (Stride), .A1 (
          CONTROLLER_nx803), .B0 (CONTROLLER_nx492)) ;
    oai221 CONTROLLER_ix157 (.Y (MemAddr[0]), .A0 (CONTROLLER_nx671), .A1 (
           CONTROLLER_nx807), .B0 (CONTROLLER_nx679), .B1 (nx7295), .C0 (
           CONTROLLER_nx685)) ;
    xnor2 CONTROLLER_ix672 (.Y (CONTROLLER_nx671), .A0 (CONTROLLER_nx673), .A1 (
          CONTROLLER_nx675)) ;
    nand02 CONTROLLER_ix674 (.Y (CONTROLLER_nx673), .A0 (CONTROLLER_nx638), .A1 (
           CONTROLLER_CurCol_0)) ;
    xnor2 CONTROLLER_ix676 (.Y (CONTROLLER_nx675), .A0 (FilterSize), .A1 (
          CONTROLLER_CurCol_1)) ;
    nand02 CONTROLLER_ix678 (.Y (CONTROLLER_nx677), .A0 (Stride), .A1 (
           CONTROLLER_nx791)) ;
    inv01 CONTROLLER_ix680 (.Y (CONTROLLER_nx679), .A (CONTROLLER_CurCol_0)) ;
    oai21 CONTROLLER_ix686 (.Y (CONTROLLER_nx685), .A0 (CONTROLLER_CurCol_0), .A1 (
          CONTROLLER_nx638), .B0 (CONTROLLER_nx142)) ;
    aoi21 CONTROLLER_ix143 (.Y (CONTROLLER_nx142), .A0 (CONTROLLER_nx638), .A1 (
          CONTROLLER_CurCol_0), .B0 (nx7297)) ;
    oai222 CONTROLLER_ix183 (.Y (MemAddr[1]), .A0 (CONTROLLER_nx691), .A1 (
           CONTROLLER_nx807), .B0 (CONTROLLER_nx599), .B1 (nx7295), .C0 (
           CONTROLLER_nx671), .C1 (nx7297)) ;
    xor2 CONTROLLER_ix692 (.Y (CONTROLLER_nx691), .A0 (CONTROLLER_CurCol_2), .A1 (
         CONTROLLER_nx693)) ;
    oai21 CONTROLLER_ix694 (.Y (CONTROLLER_nx693), .A0 (FilterSize), .A1 (
          CONTROLLER_CurCol_0), .B0 (CONTROLLER_CurCol_1)) ;
    oai222 CONTROLLER_ix201 (.Y (MemAddr[2]), .A0 (CONTROLLER_nx691), .A1 (
           nx7297), .B0 (CONTROLLER_nx696), .B1 (CONTROLLER_nx807), .C0 (
           CONTROLLER_nx699), .C1 (nx7295)) ;
    oai21 CONTROLLER_ix697 (.Y (CONTROLLER_nx696), .A0 (CONTROLLER_nx168), .A1 (
          CONTROLLER_CurCol_3), .B0 (CONTROLLER_nx701)) ;
    inv01 CONTROLLER_ix700 (.Y (CONTROLLER_nx699), .A (CONTROLLER_CurCol_2)) ;
    nand02 CONTROLLER_ix702 (.Y (CONTROLLER_nx701), .A0 (CONTROLLER_CurCol_3), .A1 (
           CONTROLLER_nx168)) ;
    oai221 CONTROLLER_ix229 (.Y (MemAddr[3]), .A0 (CONTROLLER_nx696), .A1 (
           nx7297), .B0 (CONTROLLER_nx606), .B1 (nx7295), .C0 (CONTROLLER_nx704)
           ) ;
    aoi22 CONTROLLER_ix705 (.Y (CONTROLLER_nx704), .A0 (CONTROLLER_nx803), .A1 (
          MemAddr[17]), .B0 (CONTROLLER_nx216), .B1 (CONTROLLER_nx150)) ;
    xnor2 CONTROLLER_ix217 (.Y (CONTROLLER_nx216), .A0 (CONTROLLER_CurCol_4), .A1 (
          CONTROLLER_nx701)) ;
    oai321 CONTROLLER_ix251 (.Y (MemAddr[4]), .A0 (CONTROLLER_nx709), .A1 (
           CONTROLLER_nx795), .A2 (CONTROLLER_nx791), .B0 (CONTROLLER_nx711), .B1 (
           CONTROLLER_nx807), .C0 (CONTROLLER_nx718)) ;
    inv02 CONTROLLER_ix710 (.Y (CONTROLLER_nx709), .A (CONTROLLER_CurRow_1)) ;
    oai21 CONTROLLER_ix712 (.Y (CONTROLLER_nx711), .A0 (CONTROLLER_nx210), .A1 (
          CONTROLLER_CurCol_5), .B0 (CONTROLLER_nx716)) ;
    nand02 CONTROLLER_ix717 (.Y (CONTROLLER_nx716), .A0 (CONTROLLER_CurCol_5), .A1 (
           CONTROLLER_nx210)) ;
    aoi22 CONTROLLER_ix719 (.Y (CONTROLLER_nx718), .A0 (CONTROLLER_CurCol_4), .A1 (
          CONTROLLER_nx823), .B0 (CONTROLLER_nx216), .B1 (CONTROLLER_nx829)) ;
    nor02ii CONTROLLER_ix125 (.Y (CONTROLLER_nx124), .A0 (CONTROLLER_nx793), .A1 (
            CONTROLLER_nx795)) ;
    oai221 CONTROLLER_ix273 (.Y (MemAddr[5]), .A0 (CONTROLLER_nx711), .A1 (
           nx7297), .B0 (CONTROLLER_nx613), .B1 (nx7295), .C0 (CONTROLLER_nx723)
           ) ;
    aoi22 CONTROLLER_ix724 (.Y (CONTROLLER_nx723), .A0 (CONTROLLER_CurRow_2), .A1 (
          MemAddr[17]), .B0 (CONTROLLER_nx260), .B1 (CONTROLLER_nx150)) ;
    xnor2 CONTROLLER_ix261 (.Y (CONTROLLER_nx260), .A0 (CONTROLLER_CurCol_6), .A1 (
          CONTROLLER_nx716)) ;
    oai321 CONTROLLER_ix289 (.Y (MemAddr[6]), .A0 (CONTROLLER_nx727), .A1 (
           CONTROLLER_nx795), .A2 (CONTROLLER_nx793), .B0 (CONTROLLER_nx729), .B1 (
           CONTROLLER_nx807), .C0 (CONTROLLER_nx732)) ;
    inv01 CONTROLLER_ix728 (.Y (CONTROLLER_nx727), .A (CONTROLLER_CurRow_3)) ;
    xnor2 CONTROLLER_ix730 (.Y (CONTROLLER_nx729), .A0 (CONTROLLER_nx254), .A1 (
          CONTROLLER_CurCol_7)) ;
    aoi22 CONTROLLER_ix733 (.Y (CONTROLLER_nx732), .A0 (CONTROLLER_CurCol_6), .A1 (
          CONTROLLER_nx823), .B0 (CONTROLLER_nx260), .B1 (CONTROLLER_nx829)) ;
    oai21 CONTROLLER_ix299 (.Y (MemAddr[7]), .A0 (CONTROLLER_nx729), .A1 (nx7297
          ), .B0 (CONTROLLER_nx735)) ;
    aoi22 CONTROLLER_ix736 (.Y (CONTROLLER_nx735), .A0 (CONTROLLER_CurRow_4), .A1 (
          MemAddr[17]), .B0 (CONTROLLER_CurCol_7), .B1 (CONTROLLER_nx823)) ;
    nand02 CONTROLLER_ix333 (.Y (MemAddr[8]), .A0 (CONTROLLER_nx738), .A1 (
           CONTROLLER_nx744)) ;
    aoi22 CONTROLLER_ix739 (.Y (CONTROLLER_nx738), .A0 (CONTROLLER_nx740), .A1 (
          CONTROLLER_nx829), .B0 (CONTROLLER_nx322), .B1 (CONTROLLER_nx150)) ;
    xnor2 CONTROLLER_ix323 (.Y (CONTROLLER_nx322), .A0 (CONTROLLER_nx740), .A1 (
          CONTROLLER_nx320)) ;
    aoi22 CONTROLLER_ix745 (.Y (CONTROLLER_nx744), .A0 (CONTROLLER_CurRow_5), .A1 (
          MemAddr[17]), .B0 (CONTROLLER_nx306), .B1 (CONTROLLER_nx310)) ;
    oai21 CONTROLLER_ix307 (.Y (CONTROLLER_nx306), .A0 (CONTROLLER_nx638), .A1 (
          Stride), .B0 (CONTROLLER_nx793)) ;
    oai321 CONTROLLER_ix365 (.Y (MemAddr[9]), .A0 (CONTROLLER_nx575), .A1 (
           CONTROLLER_nx797), .A2 (CONTROLLER_nx793), .B0 (CONTROLLER_nx749), .B1 (
           CONTROLLER_nx807), .C0 (CONTROLLER_nx753)) ;
    xnor2 CONTROLLER_ix750 (.Y (CONTROLLER_nx749), .A0 (CONTROLLER_CurRow_2), .A1 (
          CONTROLLER_nx751)) ;
    aoi21 CONTROLLER_ix752 (.Y (CONTROLLER_nx751), .A0 (CONTROLLER_nx805), .A1 (
          CONTROLLER_nx638), .B0 (CONTROLLER_nx799)) ;
    aoi22 CONTROLLER_ix754 (.Y (CONTROLLER_nx753), .A0 (CONTROLLER_nx801), .A1 (
          CONTROLLER_nx823), .B0 (CONTROLLER_nx322), .B1 (CONTROLLER_nx829)) ;
    oai221 CONTROLLER_ix387 (.Y (MemAddr[10]), .A0 (CONTROLLER_nx749), .A1 (
           nx7297), .B0 (CONTROLLER_nx756), .B1 (nx7295), .C0 (CONTROLLER_nx758)
           ) ;
    inv01 CONTROLLER_ix757 (.Y (CONTROLLER_nx756), .A (CONTROLLER_CurRow_2)) ;
    aoi22 CONTROLLER_ix759 (.Y (CONTROLLER_nx758), .A0 (CONTROLLER_CurRow_7), .A1 (
          MemAddr[17]), .B0 (CONTROLLER_nx374), .B1 (CONTROLLER_nx150)) ;
    nand02 CONTROLLER_ix347 (.Y (CONTROLLER_nx346), .A0 (CONTROLLER_nx751), .A1 (
           CONTROLLER_nx756)) ;
    oai222 CONTROLLER_ix405 (.Y (MemAddr[11]), .A0 (CONTROLLER_nx763), .A1 (
           CONTROLLER_nx817), .B0 (CONTROLLER_nx767), .B1 (CONTROLLER_nx807), .C0 (
           CONTROLLER_nx727), .C1 (nx7295)) ;
    aoi21 CONTROLLER_ix764 (.Y (CONTROLLER_nx763), .A0 (CONTROLLER_CurRow_3), .A1 (
          CONTROLLER_nx346), .B0 (CONTROLLER_nx765)) ;
    nor02_2x CONTROLLER_ix766 (.Y (CONTROLLER_nx765), .A0 (CONTROLLER_nx346), .A1 (
             CONTROLLER_CurRow_3)) ;
    xnor2 CONTROLLER_ix768 (.Y (CONTROLLER_nx767), .A0 (CONTROLLER_CurRow_4), .A1 (
          CONTROLLER_nx765)) ;
    oai222 CONTROLLER_ix423 (.Y (MemAddr[12]), .A0 (CONTROLLER_nx770), .A1 (
           CONTROLLER_nx809), .B0 (CONTROLLER_nx581), .B1 (CONTROLLER_nx813), .C0 (
           CONTROLLER_nx767), .C1 (CONTROLLER_nx817)) ;
    aoi21 CONTROLLER_ix771 (.Y (CONTROLLER_nx770), .A0 (CONTROLLER_CurRow_5), .A1 (
          CONTROLLER_nx390), .B0 (CONTROLLER_nx773)) ;
    nand02 CONTROLLER_ix391 (.Y (CONTROLLER_nx390), .A0 (CONTROLLER_nx765), .A1 (
           CONTROLLER_nx581)) ;
    nor02_2x CONTROLLER_ix774 (.Y (CONTROLLER_nx773), .A0 (CONTROLLER_nx390), .A1 (
             CONTROLLER_CurRow_5)) ;
    oai222 CONTROLLER_ix441 (.Y (MemAddr[13]), .A0 (CONTROLLER_nx770), .A1 (
           CONTROLLER_nx817), .B0 (CONTROLLER_nx776), .B1 (CONTROLLER_nx809), .C0 (
           CONTROLLER_nx778), .C1 (CONTROLLER_nx813)) ;
    xnor2 CONTROLLER_ix777 (.Y (CONTROLLER_nx776), .A0 (CONTROLLER_CurRow_6), .A1 (
          CONTROLLER_nx773)) ;
    inv01 CONTROLLER_ix779 (.Y (CONTROLLER_nx778), .A (CONTROLLER_CurRow_5)) ;
    oai222 CONTROLLER_ix453 (.Y (MemAddr[14]), .A0 (CONTROLLER_nx781), .A1 (
           CONTROLLER_nx809), .B0 (CONTROLLER_nx575), .B1 (CONTROLLER_nx813), .C0 (
           CONTROLLER_nx776), .C1 (CONTROLLER_nx817)) ;
    nand02 CONTROLLER_ix427 (.Y (CONTROLLER_nx426), .A0 (CONTROLLER_nx773), .A1 (
           CONTROLLER_nx575)) ;
    xnor2 CONTROLLER_ix445 (.Y (CONTROLLER_nx444), .A0 (CONTROLLER_CurRow_7), .A1 (
          CONTROLLER_nx426)) ;
    inv01 CONTROLLER_ix633 (.Y (CONTROLLER_nx632), .A (CONTROLLER_nx502)) ;
    inv01 CONTROLLER_ix493 (.Y (CONTROLLER_nx492), .A (CONTROLLER_nx634)) ;
    inv01 CONTROLLER_ix782 (.Y (CONTROLLER_nx781), .A (CONTROLLER_nx444)) ;
    inv01 CONTROLLER_ix375 (.Y (CONTROLLER_nx374), .A (CONTROLLER_nx763)) ;
    inv01 CONTROLLER_ix151 (.Y (CONTROLLER_nx150), .A (CONTROLLER_nx677)) ;
    inv01 CONTROLLER_ix15 (.Y (CONTROLLER_nx14), .A (CONTROLLER_nx571)) ;
    buf02 CONTROLLER_ix790 (.Y (CONTROLLER_nx791), .A (MemWR)) ;
    buf02 CONTROLLER_ix792 (.Y (CONTROLLER_nx793), .A (MemWR)) ;
    buf02 CONTROLLER_ix794 (.Y (CONTROLLER_nx795), .A (CacheWindowWR)) ;
    buf02 CONTROLLER_ix796 (.Y (CONTROLLER_nx797), .A (CacheWindowWR)) ;
    inv02 CONTROLLER_ix798 (.Y (CONTROLLER_nx799), .A (CONTROLLER_nx709)) ;
    inv02 CONTROLLER_ix800 (.Y (CONTROLLER_nx801), .A (CONTROLLER_nx709)) ;
    inv01 CONTROLLER_ix802 (.Y (CONTROLLER_nx803), .A (CONTROLLER_NxtRow_0)) ;
    inv01 CONTROLLER_ix804 (.Y (CONTROLLER_nx805), .A (CONTROLLER_NxtRow_0)) ;
    inv02 CONTROLLER_ix806 (.Y (CONTROLLER_nx807), .A (CONTROLLER_nx150)) ;
    inv02 CONTROLLER_ix808 (.Y (CONTROLLER_nx809), .A (CONTROLLER_nx150)) ;
    inv02 CONTROLLER_ix810 (.Y (CONTROLLER_nx811), .A (CONTROLLER_nx124)) ;
    inv02 CONTROLLER_ix812 (.Y (CONTROLLER_nx813), .A (CONTROLLER_nx823)) ;
    inv02 CONTROLLER_ix814 (.Y (CONTROLLER_nx815), .A (CONTROLLER_nx138)) ;
    inv02 CONTROLLER_ix816 (.Y (CONTROLLER_nx817), .A (CONTROLLER_nx829)) ;
    inv02 CONTROLLER_ix822 (.Y (CONTROLLER_nx823), .A (CONTROLLER_nx811)) ;
    nor02ii CONTROLLER_ix13 (.Y (CONTROLLER_nx12), .A0 (CONTROLLER_nx577), .A1 (
            CONTROLLER_CurRow_6)) ;
    nor02ii CONTROLLER_ix9 (.Y (CONTROLLER_nx8), .A0 (CONTROLLER_nx583), .A1 (
            CONTROLLER_CurRow_4)) ;
    nor02ii CONTROLLER_ix59 (.Y (CONTROLLER_nx58), .A0 (CONTROLLER_nx571), .A1 (
            Stride)) ;
    nor02ii CONTROLLER_ix71 (.Y (CONTROLLER_nx70), .A0 (CONTROLLER_nx593), .A1 (
            CONTROLLER_CurCol_1)) ;
    nor02ii CONTROLLER_ix75 (.Y (CONTROLLER_nx74), .A0 (CONTROLLER_nx602), .A1 (
            CONTROLLER_CurCol_3)) ;
    nor02ii CONTROLLER_ix79 (.Y (CONTROLLER_nx78), .A0 (CONTROLLER_nx609), .A1 (
            CONTROLLER_CurCol_5)) ;
    nor02ii CONTROLLER_ix689 (.Y (CONTROLLER_nx138), .A0 (Stride), .A1 (
            CONTROLLER_nx791)) ;
    nor02ii CONTROLLER_ix169 (.Y (CONTROLLER_nx168), .A0 (CONTROLLER_nx693), .A1 (
            CONTROLLER_CurCol_2)) ;
    nor02ii CONTROLLER_ix211 (.Y (CONTROLLER_nx210), .A0 (CONTROLLER_nx701), .A1 (
            CONTROLLER_CurCol_4)) ;
    nor02ii CONTROLLER_ix255 (.Y (CONTROLLER_nx254), .A0 (CONTROLLER_nx716), .A1 (
            CONTROLLER_CurCol_6)) ;
    nor02ii CONTROLLER_ix311 (.Y (CONTROLLER_nx310), .A0 (MemAddr[17]), .A1 (
            CONTROLLER_CurRow_0)) ;
    inv02 CONTROLLER_ix828 (.Y (CONTROLLER_nx829), .A (CONTROLLER_nx815)) ;
    dff CONTROLLER_STATE_reg_Dout_0 (.Q (CacheFilterWR), .QB (\$dummy [0]), .D (
        CONTROLLER_STATE_nx152), .CLK (CONTROLLER_STATE_NOT_CLK)) ;
    nor02_2x CONTROLLER_STATE_ix207 (.Y (CONTROLLER_STATE_nx206), .A0 (nx7285), 
             .A1 (CONTROLLER_FilterAddr_17)) ;
    inv01 CONTROLLER_STATE_ix209 (.Y (CONTROLLER_STATE_NOT_CLK), .A (CLK)) ;
    dff CONTROLLER_STATE_reg_Dout_1 (.Q (CacheWindowWR), .QB (\$dummy [1]), .D (
        CONTROLLER_STATE_nx162), .CLK (CONTROLLER_STATE_NOT_CLK)) ;
    dff CONTROLLER_STATE_reg_Dout_2 (.Q (MemWR), .QB (\$dummy [2]), .D (
        CONTROLLER_STATE_nx172), .CLK (CONTROLLER_STATE_NOT_CLK)) ;
    dff CONTROLLER_STATE_reg_Dout_3 (.Q (Calculating), .QB (\$dummy [3]), .D (
        CONTROLLER_STATE_nx182), .CLK (CONTROLLER_STATE_NOT_CLK)) ;
    dff CONTROLLER_STATE_reg_Dout_4 (.Q (Done), .QB (\$dummy [4]), .D (
        CONTROLLER_STATE_nx192), .CLK (CONTROLLER_STATE_NOT_CLK)) ;
    dff CONTROLLER_ROW_reg_Dout_0 (.Q (CONTROLLER_CurRow_0), .QB (\$dummy [5]), 
        .D (CONTROLLER_ROW_nx212), .CLK (CONTROLLER_ROW_nx327)) ;
    nor02_2x CONTROLLER_ROW_ix297 (.Y (CONTROLLER_ROW_nx296), .A0 (nx7289), .A1 (
             CONTROLLER_ROW_nx335)) ;
    inv01 CONTROLLER_ROW_ix299 (.Y (CONTROLLER_ROW_NOT_CLK), .A (CLK)) ;
    dff CONTROLLER_ROW_reg_Dout_1 (.Q (CONTROLLER_CurRow_1), .QB (\$dummy [6]), 
        .D (CONTROLLER_ROW_nx222), .CLK (CONTROLLER_ROW_nx327)) ;
    dff CONTROLLER_ROW_reg_Dout_2 (.Q (CONTROLLER_CurRow_2), .QB (\$dummy [7]), 
        .D (CONTROLLER_ROW_nx232), .CLK (CONTROLLER_ROW_nx327)) ;
    dff CONTROLLER_ROW_reg_Dout_3 (.Q (CONTROLLER_CurRow_3), .QB (\$dummy [8]), 
        .D (CONTROLLER_ROW_nx242), .CLK (CONTROLLER_ROW_nx327)) ;
    dff CONTROLLER_ROW_reg_Dout_4 (.Q (CONTROLLER_CurRow_4), .QB (\$dummy [9]), 
        .D (CONTROLLER_ROW_nx252), .CLK (CONTROLLER_ROW_nx327)) ;
    dff CONTROLLER_ROW_reg_Dout_5 (.Q (CONTROLLER_CurRow_5), .QB (\$dummy [10])
        , .D (CONTROLLER_ROW_nx262), .CLK (CONTROLLER_ROW_NOT_CLK)) ;
    dff CONTROLLER_ROW_reg_Dout_6 (.Q (CONTROLLER_CurRow_6), .QB (\$dummy [11])
        , .D (CONTROLLER_ROW_nx272), .CLK (CONTROLLER_ROW_NOT_CLK)) ;
    dff CONTROLLER_ROW_reg_Dout_7 (.Q (CONTROLLER_CurRow_7), .QB (\$dummy [12])
        , .D (CONTROLLER_ROW_nx282), .CLK (CONTROLLER_ROW_NOT_CLK)) ;
    inv01 CONTROLLER_ROW_ix326 (.Y (CONTROLLER_ROW_nx327), .A (CLK)) ;
    buf02 CONTROLLER_ROW_ix334 (.Y (CONTROLLER_ROW_nx335), .A (CONTROLLER_CntEN)
          ) ;
    buf02 CONTROLLER_ROW_ix336 (.Y (CONTROLLER_ROW_nx337), .A (CONTROLLER_CntEN)
          ) ;
    dff CONTROLLER_COL_reg_Dout_0 (.Q (CONTROLLER_CurCol_0), .QB (\$dummy [13])
        , .D (CONTROLLER_COL_nx212), .CLK (CONTROLLER_COL_nx327)) ;
    nor02_2x CONTROLLER_COL_ix297 (.Y (CONTROLLER_COL_nx296), .A0 (nx7289), .A1 (
             CONTROLLER_COL_nx335)) ;
    inv01 CONTROLLER_COL_ix299 (.Y (CONTROLLER_COL_NOT_CLK), .A (CLK)) ;
    dff CONTROLLER_COL_reg_Dout_1 (.Q (CONTROLLER_CurCol_1), .QB (\$dummy [14])
        , .D (CONTROLLER_COL_nx222), .CLK (CONTROLLER_COL_nx327)) ;
    dff CONTROLLER_COL_reg_Dout_2 (.Q (CONTROLLER_CurCol_2), .QB (\$dummy [15])
        , .D (CONTROLLER_COL_nx232), .CLK (CONTROLLER_COL_nx327)) ;
    dff CONTROLLER_COL_reg_Dout_3 (.Q (CONTROLLER_CurCol_3), .QB (\$dummy [16])
        , .D (CONTROLLER_COL_nx242), .CLK (CONTROLLER_COL_nx327)) ;
    dff CONTROLLER_COL_reg_Dout_4 (.Q (CONTROLLER_CurCol_4), .QB (\$dummy [17])
        , .D (CONTROLLER_COL_nx252), .CLK (CONTROLLER_COL_nx327)) ;
    dff CONTROLLER_COL_reg_Dout_5 (.Q (CONTROLLER_CurCol_5), .QB (\$dummy [18])
        , .D (CONTROLLER_COL_nx262), .CLK (CONTROLLER_COL_NOT_CLK)) ;
    dff CONTROLLER_COL_reg_Dout_6 (.Q (CONTROLLER_CurCol_6), .QB (\$dummy [19])
        , .D (CONTROLLER_COL_nx272), .CLK (CONTROLLER_COL_NOT_CLK)) ;
    dff CONTROLLER_COL_reg_Dout_7 (.Q (CONTROLLER_CurCol_7), .QB (\$dummy [20])
        , .D (CONTROLLER_COL_nx282), .CLK (CONTROLLER_COL_NOT_CLK)) ;
    inv01 CONTROLLER_COL_ix326 (.Y (CONTROLLER_COL_nx327), .A (CLK)) ;
    buf02 CONTROLLER_COL_ix334 (.Y (CONTROLLER_COL_nx335), .A (CONTROLLER_CntEN)
          ) ;
    buf02 CONTROLLER_COL_ix336 (.Y (CONTROLLER_COL_nx337), .A (CONTROLLER_CntEN)
          ) ;
    dffr CALC_FLIP_FLOP_1_reg_Dout (.Q (AccStartCalc), .QB (\$dummy [21]), .D (
         PWR), .CLK (Calculating), .R (CalcStartRST)) ;
    dffr CALC_FLIP_FLOP_2_reg_Dout (.Q (CalcStarted), .QB (\$dummy [22]), .D (
         nx8837), .CLK (CALC_FLIP_FLOP_2_NOT_CLK), .R (RST)) ;
    inv01 CALC_FLIP_FLOP_2_ix59 (.Y (CALC_FLIP_FLOP_2_NOT_CLK), .A (CLK)) ;
    nor02ii CALCULATOR_ix87 (.Y (CALCULATOR_CalculatingBooth), .A0 (
            CALCULATOR_nx990), .A1 (CALCULATOR_nx78)) ;
    nor04 CALCULATOR_ix991 (.Y (CALCULATOR_nx990), .A0 (CALCULATOR_CounterOut_0)
          , .A1 (CALCULATOR_CounterOut_1), .A2 (CALCULATOR_CounterOut_2), .A3 (
          CALCULATOR_CounterOut_3)) ;
    nand04 CALCULATOR_ix79 (.Y (CALCULATOR_nx78), .A0 (CALCULATOR_CounterOut_0)
           , .A1 (CALCULATOR_nx993), .A2 (CALCULATOR_nx995), .A3 (
           CALCULATOR_CounterOut_3)) ;
    inv01 CALCULATOR_ix994 (.Y (CALCULATOR_nx993), .A (CALCULATOR_CounterOut_1)
          ) ;
    inv01 CALCULATOR_ix996 (.Y (CALCULATOR_nx995), .A (CALCULATOR_CounterOut_2)
          ) ;
    nor02ii CALCULATOR_ix999 (.Y (CALCULATOR_CounterEN), .A0 (Instr), .A1 (
            CALCULATOR_nx78)) ;
    oai21 CALCULATOR_ix29 (.Y (MemDin[0]), .A0 (CALCULATOR_nx1001), .A1 (Instr)
          , .B0 (CALCULATOR_nx1003)) ;
    inv01 CALCULATOR_ix1002 (.Y (CALCULATOR_nx1001), .A (
          CALCULATOR_L5Results_1__0)) ;
    aoi32 CALCULATOR_ix1004 (.Y (CALCULATOR_nx1003), .A0 (
          CALCULATOR_L5Results_1__5), .A1 (FilterSize), .A2 (Instr), .B0 (
          CALCULATOR_L5Results_1__3), .B1 (CALCULATOR_nx22)) ;
    nor02ii CALCULATOR_ix23 (.Y (CALCULATOR_nx22), .A0 (FilterSize), .A1 (Instr)
            ) ;
    oai21 CALCULATOR_ix41 (.Y (MemDin[1]), .A0 (CALCULATOR_nx1007), .A1 (Instr)
          , .B0 (CALCULATOR_nx1009)) ;
    inv01 CALCULATOR_ix1008 (.Y (CALCULATOR_nx1007), .A (
          CALCULATOR_L5Results_1__1)) ;
    aoi32 CALCULATOR_ix1010 (.Y (CALCULATOR_nx1009), .A0 (
          CALCULATOR_L5Results_1__6), .A1 (FilterSize), .A2 (Instr), .B0 (
          CALCULATOR_L5Results_1__4), .B1 (CALCULATOR_nx22)) ;
    oai21 CALCULATOR_ix53 (.Y (MemDin[2]), .A0 (CALCULATOR_nx1012), .A1 (Instr)
          , .B0 (CALCULATOR_nx1014)) ;
    inv01 CALCULATOR_ix1013 (.Y (CALCULATOR_nx1012), .A (
          CALCULATOR_L5Results_1__2)) ;
    aoi32 CALCULATOR_ix1015 (.Y (CALCULATOR_nx1014), .A0 (
          CALCULATOR_L5Results_1__7), .A1 (FilterSize), .A2 (Instr), .B0 (
          CALCULATOR_L5Results_1__5), .B1 (CALCULATOR_nx22)) ;
    nor02ii CALCULATOR_ix3 (.Y (MemDin[5]), .A0 (Instr), .A1 (
            CALCULATOR_L5Results_1__5)) ;
    nor02ii CALCULATOR_ix7 (.Y (MemDin[6]), .A0 (Instr), .A1 (
            CALCULATOR_L5Results_1__6)) ;
    nor02ii CALCULATOR_ix11 (.Y (MemDin[7]), .A0 (Instr), .A1 (
            CALCULATOR_L5Results_1__7)) ;
    inv02 CALCULATOR_ix93 (.Y (AccFinishCalc), .A (CALCULATOR_CounterEN)) ;
    inv01 CALCULATOR_ix1042 (.Y (CALCULATOR_nx1043), .A (
          CALCULATOR_CalculatingBooth)) ;
    inv02 CALCULATOR_ix1044 (.Y (CALCULATOR_CalculatingBooth_dup_1146), .A (
          CALCULATOR_nx1043)) ;
    inv02 CALCULATOR_ix1046 (.Y (CALCULATOR_CalculatingBooth_dup_1181), .A (
          CALCULATOR_nx1043)) ;
    inv02 CALCULATOR_ix1048 (.Y (CALCULATOR_CalculatingBooth_dup_1224), .A (
          CALCULATOR_nx1043)) ;
    inv01 CALCULATOR_ix1050 (.Y (CALCULATOR_CalculatingBooth_dup_1315), .A (
          CALCULATOR_nx1043)) ;
    inv02 CALCULATOR_ix1060 (.Y (CALCULATOR_Start_dup_1144), .A (nx7303)) ;
    inv02 CALCULATOR_ix1062 (.Y (CALCULATOR_Start_dup_1149), .A (nx7303)) ;
    inv02 CALCULATOR_ix1064 (.Y (CALCULATOR_Start_dup_1154), .A (nx7303)) ;
    inv02 CALCULATOR_ix1066 (.Y (CALCULATOR_Start_dup_1159), .A (nx7303)) ;
    inv02 CALCULATOR_ix1068 (.Y (CALCULATOR_Start_dup_1164), .A (nx7303)) ;
    inv02 CALCULATOR_ix1070 (.Y (CALCULATOR_Start_dup_1169), .A (nx7303)) ;
    inv02 CALCULATOR_ix1072 (.Y (CALCULATOR_Start_dup_1174), .A (nx7303)) ;
    inv02 CALCULATOR_ix1074 (.Y (CALCULATOR_Start_dup_1179), .A (nx7307)) ;
    inv02 CALCULATOR_ix1076 (.Y (CALCULATOR_Start_dup_1184), .A (nx7307)) ;
    inv02 CALCULATOR_ix1078 (.Y (CALCULATOR_Start_dup_1189), .A (nx7307)) ;
    inv02 CALCULATOR_ix1080 (.Y (CALCULATOR_Start_dup_1194), .A (nx7307)) ;
    inv02 CALCULATOR_ix1082 (.Y (CALCULATOR_Start_dup_1199), .A (nx7307)) ;
    inv02 CALCULATOR_ix1084 (.Y (CALCULATOR_Start_dup_1204), .A (nx7307)) ;
    inv02 CALCULATOR_ix1086 (.Y (CALCULATOR_Start_dup_1209), .A (nx7307)) ;
    inv02 CALCULATOR_ix1088 (.Y (CALCULATOR_Start_dup_1222), .A (nx7311)) ;
    inv02 CALCULATOR_ix1090 (.Y (CALCULATOR_Start_dup_1235), .A (nx7311)) ;
    inv02 CALCULATOR_ix1092 (.Y (CALCULATOR_Start_dup_1248), .A (nx7311)) ;
    inv02 CALCULATOR_ix1094 (.Y (CALCULATOR_Start_dup_1261), .A (nx7311)) ;
    inv02 CALCULATOR_ix1096 (.Y (CALCULATOR_Start_dup_1274), .A (nx7311)) ;
    inv02 CALCULATOR_ix1098 (.Y (CALCULATOR_Start_dup_1287), .A (nx7311)) ;
    inv02 CALCULATOR_ix1100 (.Y (CALCULATOR_Start_dup_1300), .A (nx7311)) ;
    inv02 CALCULATOR_ix1102 (.Y (CALCULATOR_Start_dup_1313), .A (nx7299)) ;
    inv02 CALCULATOR_ix1104 (.Y (CALCULATOR_Start_dup_1326), .A (nx7299)) ;
    inv02 CALCULATOR_ix1106 (.Y (CALCULATOR_Start_dup_1339), .A (nx7299)) ;
    inv02 CALCULATOR_ix1108 (.Y (CALCULATOR_Start_dup_1352), .A (nx7299)) ;
    inv02 CALCULATOR_ix1110 (.Y (CALCULATOR_nx1111), .A (AccStartCalc)) ;
    dffr CALCULATOR_ACCELERATOR_COUNTER_reg_Dout_0 (.Q (CALCULATOR_CounterOut_0)
         , .QB (\$dummy [23]), .D (CALCULATOR_ACCELERATOR_COUNTER_nx81), .CLK (
         CLK), .R (CALCULATOR_CounterRST)) ;
    dffr CALCULATOR_ACCELERATOR_COUNTER_reg_Dout_1 (.Q (CALCULATOR_CounterOut_1)
         , .QB (\$dummy [24]), .D (CALCULATOR_ACCELERATOR_COUNTER_nx91), .CLK (
         CLK), .R (CALCULATOR_CounterRST)) ;
    xor2 CALCULATOR_ACCELERATOR_COUNTER_ix7 (.Y (
         CALCULATOR_ACCELERATOR_COUNTER_nx6), .A0 (CALCULATOR_CounterOut_1), .A1 (
         CALCULATOR_CounterOut_0)) ;
    dffr CALCULATOR_ACCELERATOR_COUNTER_reg_Dout_2 (.Q (CALCULATOR_CounterOut_2)
         , .QB (\$dummy [25]), .D (CALCULATOR_ACCELERATOR_COUNTER_nx101), .CLK (
         CLK), .R (CALCULATOR_CounterRST)) ;
    xnor2 CALCULATOR_ACCELERATOR_COUNTER_ix13 (.Y (
          CALCULATOR_ACCELERATOR_COUNTER_nx12), .A0 (CALCULATOR_CounterOut_2), .A1 (
          CALCULATOR_ACCELERATOR_COUNTER_nx133)) ;
    nand02 CALCULATOR_ACCELERATOR_COUNTER_ix134 (.Y (
           CALCULATOR_ACCELERATOR_COUNTER_nx133), .A0 (CALCULATOR_CounterOut_1)
           , .A1 (CALCULATOR_CounterOut_0)) ;
    dffr CALCULATOR_ACCELERATOR_COUNTER_reg_Dout_3 (.Q (CALCULATOR_CounterOut_3)
         , .QB (\$dummy [26]), .D (CALCULATOR_ACCELERATOR_COUNTER_nx111), .CLK (
         CLK), .R (CALCULATOR_CounterRST)) ;
    xnor2 CALCULATOR_ACCELERATOR_COUNTER_ix19 (.Y (
          CALCULATOR_ACCELERATOR_COUNTER_nx18), .A0 (CALCULATOR_CounterOut_3), .A1 (
          CALCULATOR_ACCELERATOR_COUNTER_nx139)) ;
    nand03 CALCULATOR_ACCELERATOR_COUNTER_ix140 (.Y (
           CALCULATOR_ACCELERATOR_COUNTER_nx139), .A0 (CALCULATOR_CounterOut_2)
           , .A1 (CALCULATOR_CounterOut_1), .A2 (CALCULATOR_CounterOut_0)) ;
    xor2 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix83 (.Y (CALCULATOR_L1Results_0__0), 
         .A0 (CALCULATOR_L1SecondOperands_0__0), .A1 (
         CALCULATOR_L1FirstOperands_0__0)) ;
    xnor2 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix380 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx379), .A0 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx381), .A1 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx383)) ;
    nand02 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix382 (.Y (
           CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx381), .A0 (
           CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothOperand_0), .A1 (nx7323)) ;
    xnor2 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix384 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx383), .A0 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothOperand_1), .A1 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_1)) ;
    inv01 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix388 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx387), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_2)) ;
    xnor2 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix390 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx389), .A0 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx391), .A1 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx395)) ;
    aoi32 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix392 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx391), .A0 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothOperand_0), .A1 (nx7323), .A2 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx154), .B0 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_1), .B1 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothOperand_1)) ;
    xnor2 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix396 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx395), .A0 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothOperand_2), .A1 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_2)) ;
    inv01 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix400 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx399), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_3)) ;
    xnor2 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix402 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx401), .A0 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx403), .A1 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx405)) ;
    xnor2 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix406 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx405), .A0 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothOperand_3), .A1 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_3)) ;
    inv01 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix410 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx409), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_4)) ;
    xnor2 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix412 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx411), .A0 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx413), .A1 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx415)) ;
    xnor2 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix416 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx415), .A0 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothOperand_4), .A1 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_4)) ;
    inv01 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix420 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx419), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_5)) ;
    xnor2 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix422 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx421), .A0 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx423), .A1 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx425)) ;
    xnor2 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix426 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx425), .A0 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothOperand_5), .A1 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_5)) ;
    inv01 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix430 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx429), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_6)) ;
    xnor2 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix432 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx431), .A0 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx433), .A1 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx435)) ;
    xnor2 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix436 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx435), .A0 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothOperand_6), .A1 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_6)) ;
    inv01 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix440 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx439), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_7)) ;
    xnor2 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix442 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx441), .A0 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx443), .A1 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx445)) ;
    xnor2 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix446 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx445), .A0 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothOperand_7), .A1 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_7)) ;
    inv01 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix450 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx449), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_8)) ;
    xnor2 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix452 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx451), .A0 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx453), .A1 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx455)) ;
    xnor2 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix456 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx455), .A0 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothOperand_8), .A1 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_8)) ;
    xor2 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix317 (.Y (
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx316), .A0 (
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx461), .A1 (
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx463)) ;
    xnor2 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix464 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx463), .A0 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothOperand_9), .A1 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_9)) ;
    xor2 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix337 (.Y (
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx336), .A0 (
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx467), .A1 (
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx471)) ;
    inv01 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix470 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx469), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_9)) ;
    xnor2 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix472 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx471), .A0 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothOperand_10), .A1 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_10)) ;
    xor2 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix357 (.Y (
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx356), .A0 (
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx475), .A1 (
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx479)) ;
    inv01 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix478 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx477), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_10)) ;
    xnor2 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix480 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx479), .A0 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothOperand_11), .A1 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_11)) ;
    xor2 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix377 (.Y (
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx376), .A0 (
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx483), .A1 (
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx487)) ;
    inv01 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix486 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx485), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_11)) ;
    xnor2 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix488 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx487), .A0 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothOperand_12), .A1 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_12)) ;
    xor2 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix397 (.Y (
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx396), .A0 (
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx491), .A1 (
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx495)) ;
    inv01 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix494 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx493), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_12)) ;
    xnor2 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix496 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx495), .A0 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothOperand_13), .A1 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_13)) ;
    xor2 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix417 (.Y (
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx416), .A0 (
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx499), .A1 (
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx503)) ;
    inv01 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix502 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx501), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_13)) ;
    xnor2 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix504 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx503), .A0 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothOperand_14), .A1 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_14)) ;
    xor2 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix437 (.Y (
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx436), .A0 (
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx507), .A1 (
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx511)) ;
    inv01 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix510 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx509), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_14)) ;
    xnor2 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix512 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx511), .A0 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothOperand_15), .A1 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_15)) ;
    xnor2 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix457 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx456), .A0 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx515), .A1 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx454)) ;
    inv01 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix518 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx517), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_15)) ;
    xor2 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix455 (.Y (
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx454), .A0 (
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothOperand_16), .A1 (
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_16)) ;
    mux21_ni CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix91 (.Y (
             CALCULATOR_L1SecondOperands_0__0), .A0 (
             CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_1), .A1 (
             CacheWindow_0__0__0), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix99 (.Y (
             CALCULATOR_L1SecondOperands_0__1), .A0 (
             CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_2), .A1 (
             CacheWindow_0__0__1), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix107 (.Y (
             CALCULATOR_L1SecondOperands_0__2), .A0 (
             CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_3), .A1 (
             CacheWindow_0__0__2), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix115 (.Y (
             CALCULATOR_L1SecondOperands_0__3), .A0 (
             CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_4), .A1 (
             CacheWindow_0__0__3), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix123 (.Y (
             CALCULATOR_L1SecondOperands_0__4), .A0 (
             CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_5), .A1 (
             CacheWindow_0__0__4), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix131 (.Y (
             CALCULATOR_L1SecondOperands_0__5), .A0 (
             CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_6), .A1 (
             CacheWindow_0__0__5), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix139 (.Y (
             CALCULATOR_L1SecondOperands_0__6), .A0 (
             CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_7), .A1 (
             CacheWindow_0__0__6), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix147 (.Y (
             CALCULATOR_L1SecondOperands_0__7), .A0 (
             CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_8), .A1 (
             CacheWindow_0__0__7), .S0 (Instr)) ;
    xor2 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix77 (.Y (CALCULATOR_L1Results_0__1), 
         .A0 (CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx529), .A1 (
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx531)) ;
    nand02 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix530 (.Y (
           CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx529), .A0 (
           CALCULATOR_L1SecondOperands_0__0), .A1 (
           CALCULATOR_L1FirstOperands_0__0)) ;
    xnor2 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix532 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx531), .A0 (
          CALCULATOR_L1SecondOperands_0__1), .A1 (
          CALCULATOR_L1FirstOperands_0__1)) ;
    xor2 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix75 (.Y (CALCULATOR_L1Results_0__2), 
         .A0 (CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx534), .A1 (
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx537)) ;
    aoi32 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix535 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx534), .A0 (
          CALCULATOR_L1SecondOperands_0__0), .A1 (
          CALCULATOR_L1FirstOperands_0__0), .A2 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx30), .B0 (
          CALCULATOR_L1FirstOperands_0__1), .B1 (
          CALCULATOR_L1SecondOperands_0__1)) ;
    xnor2 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix538 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx537), .A0 (
          CALCULATOR_L1SecondOperands_0__2), .A1 (
          CALCULATOR_L1FirstOperands_0__2)) ;
    xor2 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix73 (.Y (CALCULATOR_L1Results_0__3), 
         .A0 (CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx540), .A1 (
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx544)) ;
    aoi22 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix541 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx540), .A0 (
          CALCULATOR_L1FirstOperands_0__2), .A1 (
          CALCULATOR_L1SecondOperands_0__2), .B0 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx40), .B1 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx24)) ;
    xnor2 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix545 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx544), .A0 (
          CALCULATOR_L1SecondOperands_0__3), .A1 (
          CALCULATOR_L1FirstOperands_0__3)) ;
    xor2 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix71 (.Y (CALCULATOR_L1Results_0__4), 
         .A0 (CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx547), .A1 (
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx551)) ;
    aoi22 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix548 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx547), .A0 (
          CALCULATOR_L1FirstOperands_0__3), .A1 (
          CALCULATOR_L1SecondOperands_0__3), .B0 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx44), .B1 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx18)) ;
    xnor2 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix552 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx551), .A0 (
          CALCULATOR_L1SecondOperands_0__4), .A1 (
          CALCULATOR_L1FirstOperands_0__4)) ;
    xor2 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix69 (.Y (CALCULATOR_L1Results_0__5), 
         .A0 (CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx554), .A1 (
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx558)) ;
    aoi22 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix555 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx554), .A0 (
          CALCULATOR_L1FirstOperands_0__4), .A1 (
          CALCULATOR_L1SecondOperands_0__4), .B0 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx48), .B1 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx12)) ;
    xnor2 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix559 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx558), .A0 (
          CALCULATOR_L1SecondOperands_0__5), .A1 (
          CALCULATOR_L1FirstOperands_0__5)) ;
    xor2 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix67 (.Y (CALCULATOR_L1Results_0__6), 
         .A0 (CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx561), .A1 (
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx565)) ;
    aoi22 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix562 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx561), .A0 (
          CALCULATOR_L1FirstOperands_0__5), .A1 (
          CALCULATOR_L1SecondOperands_0__5), .B0 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx52), .B1 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx6)) ;
    xnor2 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix566 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx565), .A0 (
          CALCULATOR_L1SecondOperands_0__6), .A1 (
          CALCULATOR_L1FirstOperands_0__6)) ;
    xnor2 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix65 (.Y (CALCULATOR_L1Results_0__7)
          , .A0 (CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx568), .A1 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx62)) ;
    aoi22 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix569 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx568), .A0 (
          CALCULATOR_L1FirstOperands_0__6), .A1 (
          CALCULATOR_L1SecondOperands_0__6), .B0 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx56), .B1 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx0)) ;
    xor2 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix63 (.Y (
         CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx62), .A0 (
         CALCULATOR_L1SecondOperands_0__7), .A1 (CALCULATOR_L1FirstOperands_0__7
         )) ;
    inv01 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix155 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx154), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx383)) ;
    inv01 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix57 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx56), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx561)) ;
    inv01 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix53 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx52), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx554)) ;
    inv01 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix49 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx48), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx547)) ;
    inv01 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix45 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx44), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx540)) ;
    inv01 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix41 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx40), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx534)) ;
    inv01 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix31 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx30), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx531)) ;
    inv01 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix25 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx24), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx537)) ;
    inv01 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix19 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx18), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx544)) ;
    inv01 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix13 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx12), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx551)) ;
    inv01 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix7 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx6), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx558)) ;
    inv01 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix1 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx0), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx565)) ;
    fake_gnd CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix216 (.Y (
             CALCULATOR_L1_0_L2_0_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    aoi21 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix77 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_10), .A0 (
          CacheFilter_0__0__1), .A1 (CacheFilter_0__0__0), .B0 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx4)) ;
    nor02_2x CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix5 (.Y (
             CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx4), .A0 (
             CacheFilter_0__0__0), .A1 (CacheFilter_0__0__1)) ;
    aoi21 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix67 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_11), .A0 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx328), .A1 (
          CacheFilter_0__0__2), .B0 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx8)) ;
    nor03_2x CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix9 (.Y (
             CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx8), .A0 (
             CacheFilter_0__0__2), .A1 (CacheFilter_0__0__0), .A2 (
             CacheFilter_0__0__1)) ;
    xnor2 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix59 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_12), .A0 (
          CacheFilter_0__0__3), .A1 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx8)) ;
    xnor2 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix51 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_13), .A0 (
          CacheFilter_0__0__4), .A1 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx12)) ;
    nor04 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix13 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx12), .A0 (
          CacheFilter_0__0__3), .A1 (CacheFilter_0__0__2), .A2 (
          CacheFilter_0__0__0), .A3 (CacheFilter_0__0__1)) ;
    xnor2 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix43 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_14), .A0 (
          CacheFilter_0__0__5), .A1 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx16)) ;
    nor02ii CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix17 (.Y (
            CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx16), .A0 (
            CacheFilter_0__0__4), .A1 (
            CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx12)) ;
    xnor2 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix35 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_15), .A0 (
          CacheFilter_0__0__6), .A1 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx20)) ;
    nor02ii CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix21 (.Y (
            CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx20), .A0 (
            CacheFilter_0__0__5), .A1 (
            CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx16)) ;
    xnor2 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix27 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_16), .A0 (
          CacheFilter_0__0__7), .A1 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx24)) ;
    nor02ii CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix25 (.Y (
            CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx24), .A0 (
            CacheFilter_0__0__6), .A1 (
            CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx20)) ;
    inv01 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix329 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx328), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx4)) ;
    inv02 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix383 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx384), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_0)) ;
    dff CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_0 (.Q (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_0), .QB (
        \$dummy [27]), .D (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .CLK (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    inv01 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix565 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx564), .A (RST
          )) ;
    nor02_2x CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix567 (.Y (
             CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566), .A0 (
             RST), .A1 (
             CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644)) ;
    dff CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_1 (.Q (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_1), .QB (
        \$dummy [28]), .D (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .CLK (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_2 (.Q (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_2), .QB (
        \$dummy [29]), .D (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .CLK (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_3 (.Q (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_3), .QB (
        \$dummy [30]), .D (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .CLK (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_4 (.Q (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_4), .QB (
        \$dummy [31]), .D (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .CLK (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_5 (.Q (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_5), .QB (
        \$dummy [32]), .D (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .CLK (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_6 (.Q (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_6), .QB (
        \$dummy [33]), .D (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .CLK (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_7 (.Q (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_7), .QB (
        \$dummy [34]), .D (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .CLK (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_8 (.Q (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_8), .QB (
        \$dummy [35]), .D (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .CLK (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_9 (.Q (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_9), .QB (
        \$dummy [36]), .D (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .CLK (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_10 (.Q (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_10), .QB (
        \$dummy [37]), .D (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .CLK (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_11 (.Q (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_11), .QB (
        \$dummy [38]), .D (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .CLK (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_12 (.Q (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_12), .QB (
        \$dummy [39]), .D (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .CLK (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_13 (.Q (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_13), .QB (
        \$dummy [40]), .D (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .CLK (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_14 (.Q (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_14), .QB (
        \$dummy [41]), .D (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .CLK (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_15 (.Q (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_15), .QB (
        \$dummy [42]), .D (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .CLK (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_16 (.Q (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_16), .QB (
        \$dummy [43]), .D (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .CLK (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    inv02 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix623 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix625 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix627 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix643 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644), .A (
          nx7379)) ;
    dff CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_0 (.Q (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_0), .QB (
        \$dummy [44]), .D (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .CLK (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    nor02_2x CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix567 (.Y (
             CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566), .A0 (
             RST), .A1 (
             CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644)) ;
    dff CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_1 (.Q (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_1), .QB (
        \$dummy [45]), .D (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .CLK (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_2 (.Q (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_2), .QB (
        \$dummy [46]), .D (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .CLK (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_3 (.Q (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_3), .QB (
        \$dummy [47]), .D (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .CLK (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_4 (.Q (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_4), .QB (
        \$dummy [48]), .D (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .CLK (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_5 (.Q (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_5), .QB (
        \$dummy [49]), .D (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .CLK (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_6 (.Q (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_6), .QB (
        \$dummy [50]), .D (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .CLK (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_7 (.Q (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_7), .QB (
        \$dummy [51]), .D (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .CLK (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_8 (.Q (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_8), .QB (
        \$dummy [52]), .D (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .CLK (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_9 (.Q (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_9), .QB (
        \$dummy [53]), .D (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .CLK (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_10 (.Q (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_10), .QB (
        \$dummy [54]), .D (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .CLK (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_11 (.Q (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_11), .QB (
        \$dummy [55]), .D (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .CLK (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_12 (.Q (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_12), .QB (
        \$dummy [56]), .D (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .CLK (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_13 (.Q (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_13), .QB (
        \$dummy [57]), .D (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .CLK (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_14 (.Q (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_14), .QB (
        \$dummy [58]), .D (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .CLK (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_15 (.Q (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_15), .QB (
        \$dummy [59]), .D (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .CLK (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_16 (.Q (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_16), .QB (
        \$dummy [60]), .D (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .CLK (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    inv02 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix623 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix625 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix627 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix643 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644), .A (
          nx7385)) ;
    dff CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_0 (.Q (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_0), .QB (\$dummy [61]), .D (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .CLK (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    nor02_2x CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix567 (.Y (
             CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566), .A0 (
             RST), .A1 (
             CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    dff CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_1 (.Q (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_1), .QB (\$dummy [62]), .D (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .CLK (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_2 (.Q (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_2), .QB (\$dummy [63]), .D (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .CLK (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_3 (.Q (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_3), .QB (\$dummy [64]), .D (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .CLK (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_4 (.Q (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_4), .QB (\$dummy [65]), .D (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .CLK (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_5 (.Q (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_5), .QB (\$dummy [66]), .D (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .CLK (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_6 (.Q (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_6), .QB (\$dummy [67]), .D (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .CLK (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_7 (.Q (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_7), .QB (\$dummy [68]), .D (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .CLK (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_8 (.Q (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_8), .QB (\$dummy [69]), .D (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .CLK (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_9 (.Q (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_9), .QB (\$dummy [70]), .D (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .CLK (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_10 (.Q (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_10), .QB (\$dummy [71]), .D (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .CLK (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_11 (.Q (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_11), .QB (\$dummy [72]), .D (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .CLK (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_12 (.Q (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_12), .QB (\$dummy [73]), .D (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .CLK (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_13 (.Q (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_13), .QB (\$dummy [74]), .D (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .CLK (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_14 (.Q (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_14), .QB (\$dummy [75]), .D (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .CLK (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_15 (.Q (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_15), .QB (\$dummy [76]), .D (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .CLK (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_16 (.Q (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_16), .QB (\$dummy [77]), .D (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .CLK (
        CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    inv02 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix623 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix625 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix627 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix643 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642)) ;
    xor2 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix83 (.Y (CALCULATOR_L1Results_1__0), 
         .A0 (CALCULATOR_L1SecondOperands_1__0), .A1 (
         CALCULATOR_L1FirstOperands_1__0)) ;
    xnor2 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix380 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx379), .A0 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx381), .A1 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx383)) ;
    nand02 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix382 (.Y (
           CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx381), .A0 (
           CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothOperand_0), .A1 (nx7405)) ;
    xnor2 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix384 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx383), .A0 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothOperand_1), .A1 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_1)) ;
    inv01 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix388 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx387), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_2)) ;
    xnor2 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix390 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx389), .A0 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx391), .A1 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx395)) ;
    aoi32 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix392 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx391), .A0 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothOperand_0), .A1 (nx7405), .A2 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx154), .B0 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_1), .B1 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothOperand_1)) ;
    xnor2 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix396 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx395), .A0 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothOperand_2), .A1 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_2)) ;
    inv01 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix400 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx399), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_3)) ;
    xnor2 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix402 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx401), .A0 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx403), .A1 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx405)) ;
    xnor2 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix406 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx405), .A0 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothOperand_3), .A1 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_3)) ;
    inv01 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix410 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx409), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_4)) ;
    xnor2 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix412 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx411), .A0 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx413), .A1 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx415)) ;
    xnor2 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix416 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx415), .A0 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothOperand_4), .A1 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_4)) ;
    inv01 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix420 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx419), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_5)) ;
    xnor2 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix422 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx421), .A0 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx423), .A1 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx425)) ;
    xnor2 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix426 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx425), .A0 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothOperand_5), .A1 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_5)) ;
    inv01 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix430 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx429), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_6)) ;
    xnor2 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix432 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx431), .A0 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx433), .A1 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx435)) ;
    xnor2 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix436 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx435), .A0 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothOperand_6), .A1 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_6)) ;
    inv01 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix440 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx439), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_7)) ;
    xnor2 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix442 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx441), .A0 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx443), .A1 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx445)) ;
    xnor2 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix446 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx445), .A0 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothOperand_7), .A1 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_7)) ;
    inv01 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix450 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx449), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_8)) ;
    xnor2 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix452 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx451), .A0 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx453), .A1 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx455)) ;
    xnor2 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix456 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx455), .A0 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothOperand_8), .A1 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_8)) ;
    xor2 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix317 (.Y (
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx316), .A0 (
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx461), .A1 (
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx463)) ;
    xnor2 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix464 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx463), .A0 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothOperand_9), .A1 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_9)) ;
    xor2 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix337 (.Y (
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx336), .A0 (
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx467), .A1 (
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx471)) ;
    inv01 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix470 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx469), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_9)) ;
    xnor2 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix472 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx471), .A0 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothOperand_10), .A1 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_10)) ;
    xor2 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix357 (.Y (
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx356), .A0 (
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx475), .A1 (
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx479)) ;
    inv01 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix478 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx477), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_10)) ;
    xnor2 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix480 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx479), .A0 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothOperand_11), .A1 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_11)) ;
    xor2 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix377 (.Y (
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx376), .A0 (
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx483), .A1 (
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx487)) ;
    inv01 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix486 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx485), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_11)) ;
    xnor2 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix488 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx487), .A0 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothOperand_12), .A1 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_12)) ;
    xor2 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix397 (.Y (
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx396), .A0 (
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx491), .A1 (
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx495)) ;
    inv01 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix494 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx493), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_12)) ;
    xnor2 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix496 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx495), .A0 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothOperand_13), .A1 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_13)) ;
    xor2 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix417 (.Y (
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx416), .A0 (
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx499), .A1 (
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx503)) ;
    inv01 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix502 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx501), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_13)) ;
    xnor2 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix504 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx503), .A0 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothOperand_14), .A1 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_14)) ;
    xor2 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix437 (.Y (
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx436), .A0 (
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx507), .A1 (
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx511)) ;
    inv01 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix510 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx509), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_14)) ;
    xnor2 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix512 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx511), .A0 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothOperand_15), .A1 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_15)) ;
    xnor2 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix457 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx456), .A0 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx515), .A1 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx454)) ;
    inv01 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix518 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx517), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_15)) ;
    xor2 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix455 (.Y (
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx454), .A0 (
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothOperand_16), .A1 (
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_16)) ;
    mux21_ni CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix91 (.Y (
             CALCULATOR_L1SecondOperands_1__0), .A0 (
             CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_1), .A1 (
             CacheWindow_0__1__0), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix99 (.Y (
             CALCULATOR_L1SecondOperands_1__1), .A0 (
             CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_2), .A1 (
             CacheWindow_0__1__1), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix107 (.Y (
             CALCULATOR_L1SecondOperands_1__2), .A0 (
             CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_3), .A1 (
             CacheWindow_0__1__2), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix115 (.Y (
             CALCULATOR_L1SecondOperands_1__3), .A0 (
             CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_4), .A1 (
             CacheWindow_0__1__3), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix123 (.Y (
             CALCULATOR_L1SecondOperands_1__4), .A0 (
             CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_5), .A1 (
             CacheWindow_0__1__4), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix131 (.Y (
             CALCULATOR_L1SecondOperands_1__5), .A0 (
             CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_6), .A1 (
             CacheWindow_0__1__5), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix139 (.Y (
             CALCULATOR_L1SecondOperands_1__6), .A0 (
             CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_7), .A1 (
             CacheWindow_0__1__6), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix147 (.Y (
             CALCULATOR_L1SecondOperands_1__7), .A0 (
             CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_8), .A1 (
             CacheWindow_0__1__7), .S0 (Instr)) ;
    xor2 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix77 (.Y (CALCULATOR_L1Results_1__1), 
         .A0 (CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx529), .A1 (
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx531)) ;
    nand02 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix530 (.Y (
           CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx529), .A0 (
           CALCULATOR_L1SecondOperands_1__0), .A1 (
           CALCULATOR_L1FirstOperands_1__0)) ;
    xnor2 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix532 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx531), .A0 (
          CALCULATOR_L1SecondOperands_1__1), .A1 (
          CALCULATOR_L1FirstOperands_1__1)) ;
    xor2 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix75 (.Y (CALCULATOR_L1Results_1__2), 
         .A0 (CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx534), .A1 (
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx537)) ;
    aoi32 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix535 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx534), .A0 (
          CALCULATOR_L1SecondOperands_1__0), .A1 (
          CALCULATOR_L1FirstOperands_1__0), .A2 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx30), .B0 (
          CALCULATOR_L1FirstOperands_1__1), .B1 (
          CALCULATOR_L1SecondOperands_1__1)) ;
    xnor2 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix538 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx537), .A0 (
          CALCULATOR_L1SecondOperands_1__2), .A1 (
          CALCULATOR_L1FirstOperands_1__2)) ;
    xor2 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix73 (.Y (CALCULATOR_L1Results_1__3), 
         .A0 (CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx540), .A1 (
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx544)) ;
    aoi22 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix541 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx540), .A0 (
          CALCULATOR_L1FirstOperands_1__2), .A1 (
          CALCULATOR_L1SecondOperands_1__2), .B0 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx40), .B1 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx24)) ;
    xnor2 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix545 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx544), .A0 (
          CALCULATOR_L1SecondOperands_1__3), .A1 (
          CALCULATOR_L1FirstOperands_1__3)) ;
    xor2 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix71 (.Y (CALCULATOR_L1Results_1__4), 
         .A0 (CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx547), .A1 (
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx551)) ;
    aoi22 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix548 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx547), .A0 (
          CALCULATOR_L1FirstOperands_1__3), .A1 (
          CALCULATOR_L1SecondOperands_1__3), .B0 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx44), .B1 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx18)) ;
    xnor2 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix552 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx551), .A0 (
          CALCULATOR_L1SecondOperands_1__4), .A1 (
          CALCULATOR_L1FirstOperands_1__4)) ;
    xor2 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix69 (.Y (CALCULATOR_L1Results_1__5), 
         .A0 (CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx554), .A1 (
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx558)) ;
    aoi22 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix555 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx554), .A0 (
          CALCULATOR_L1FirstOperands_1__4), .A1 (
          CALCULATOR_L1SecondOperands_1__4), .B0 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx48), .B1 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx12)) ;
    xnor2 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix559 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx558), .A0 (
          CALCULATOR_L1SecondOperands_1__5), .A1 (
          CALCULATOR_L1FirstOperands_1__5)) ;
    xor2 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix67 (.Y (CALCULATOR_L1Results_1__6), 
         .A0 (CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx561), .A1 (
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx565)) ;
    aoi22 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix562 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx561), .A0 (
          CALCULATOR_L1FirstOperands_1__5), .A1 (
          CALCULATOR_L1SecondOperands_1__5), .B0 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx52), .B1 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx6)) ;
    xnor2 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix566 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx565), .A0 (
          CALCULATOR_L1SecondOperands_1__6), .A1 (
          CALCULATOR_L1FirstOperands_1__6)) ;
    xnor2 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix65 (.Y (CALCULATOR_L1Results_1__7)
          , .A0 (CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx568), .A1 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx62)) ;
    aoi22 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix569 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx568), .A0 (
          CALCULATOR_L1FirstOperands_1__6), .A1 (
          CALCULATOR_L1SecondOperands_1__6), .B0 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx56), .B1 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx0)) ;
    xor2 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix63 (.Y (
         CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx62), .A0 (
         CALCULATOR_L1SecondOperands_1__7), .A1 (CALCULATOR_L1FirstOperands_1__7
         )) ;
    inv01 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix155 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx154), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx383)) ;
    inv01 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix57 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx56), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx561)) ;
    inv01 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix53 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx52), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx554)) ;
    inv01 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix49 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx48), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx547)) ;
    inv01 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix45 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx44), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx540)) ;
    inv01 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix41 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx40), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx534)) ;
    inv01 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix31 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx30), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx531)) ;
    inv01 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix25 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx24), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx537)) ;
    inv01 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix19 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx18), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx544)) ;
    inv01 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix13 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx12), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx551)) ;
    inv01 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix7 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx6), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx558)) ;
    inv01 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix1 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx0), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx565)) ;
    fake_gnd CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix216 (.Y (
             CALCULATOR_L1_0_L2_1_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    aoi21 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix77 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_10), .A0 (
          CacheFilter_0__1__1), .A1 (CacheFilter_0__1__0), .B0 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx4)) ;
    nor02_2x CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix5 (.Y (
             CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx4), .A0 (
             CacheFilter_0__1__0), .A1 (CacheFilter_0__1__1)) ;
    aoi21 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix67 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_11), .A0 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx328), .A1 (
          CacheFilter_0__1__2), .B0 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx8)) ;
    nor03_2x CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix9 (.Y (
             CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx8), .A0 (
             CacheFilter_0__1__2), .A1 (CacheFilter_0__1__0), .A2 (
             CacheFilter_0__1__1)) ;
    xnor2 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix59 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_12), .A0 (
          CacheFilter_0__1__3), .A1 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx8)) ;
    xnor2 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix51 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_13), .A0 (
          CacheFilter_0__1__4), .A1 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx12)) ;
    nor04 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix13 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx12), .A0 (
          CacheFilter_0__1__3), .A1 (CacheFilter_0__1__2), .A2 (
          CacheFilter_0__1__0), .A3 (CacheFilter_0__1__1)) ;
    xnor2 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix43 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_14), .A0 (
          CacheFilter_0__1__5), .A1 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx16)) ;
    nor02ii CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix17 (.Y (
            CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx16), .A0 (
            CacheFilter_0__1__4), .A1 (
            CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx12)) ;
    xnor2 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix35 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_15), .A0 (
          CacheFilter_0__1__6), .A1 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx20)) ;
    nor02ii CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix21 (.Y (
            CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx20), .A0 (
            CacheFilter_0__1__5), .A1 (
            CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx16)) ;
    xnor2 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix27 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_16), .A0 (
          CacheFilter_0__1__7), .A1 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx24)) ;
    nor02ii CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix25 (.Y (
            CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx24), .A0 (
            CacheFilter_0__1__6), .A1 (
            CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx20)) ;
    inv01 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix329 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx328), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx4)) ;
    inv02 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix383 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx384), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_0)) ;
    dff CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_0 (.Q (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_0), .QB (
        \$dummy [78]), .D (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .CLK (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    nor02_2x CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix567 (.Y (
             CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566), .A0 (
             RST), .A1 (
             CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644)) ;
    dff CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_1 (.Q (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_1), .QB (
        \$dummy [79]), .D (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .CLK (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_2 (.Q (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_2), .QB (
        \$dummy [80]), .D (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .CLK (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_3 (.Q (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_3), .QB (
        \$dummy [81]), .D (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .CLK (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_4 (.Q (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_4), .QB (
        \$dummy [82]), .D (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .CLK (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_5 (.Q (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_5), .QB (
        \$dummy [83]), .D (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .CLK (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_6 (.Q (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_6), .QB (
        \$dummy [84]), .D (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .CLK (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_7 (.Q (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_7), .QB (
        \$dummy [85]), .D (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .CLK (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_8 (.Q (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_8), .QB (
        \$dummy [86]), .D (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .CLK (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_9 (.Q (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_9), .QB (
        \$dummy [87]), .D (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .CLK (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_10 (.Q (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_10), .QB (
        \$dummy [88]), .D (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .CLK (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_11 (.Q (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_11), .QB (
        \$dummy [89]), .D (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .CLK (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_12 (.Q (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_12), .QB (
        \$dummy [90]), .D (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .CLK (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_13 (.Q (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_13), .QB (
        \$dummy [91]), .D (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .CLK (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_14 (.Q (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_14), .QB (
        \$dummy [92]), .D (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .CLK (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_15 (.Q (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_15), .QB (
        \$dummy [93]), .D (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .CLK (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_16 (.Q (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_16), .QB (
        \$dummy [94]), .D (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .CLK (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    inv02 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix623 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix625 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix627 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix643 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644), .A (
          nx7419)) ;
    dff CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_0 (.Q (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_0), .QB (
        \$dummy [95]), .D (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .CLK (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    nor02_2x CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix567 (.Y (
             CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566), .A0 (
             RST), .A1 (
             CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644)) ;
    dff CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_1 (.Q (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_1), .QB (
        \$dummy [96]), .D (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .CLK (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_2 (.Q (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_2), .QB (
        \$dummy [97]), .D (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .CLK (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_3 (.Q (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_3), .QB (
        \$dummy [98]), .D (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .CLK (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_4 (.Q (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_4), .QB (
        \$dummy [99]), .D (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .CLK (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_5 (.Q (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_5), .QB (
        \$dummy [100]), .D (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .CLK (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_6 (.Q (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_6), .QB (
        \$dummy [101]), .D (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .CLK (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_7 (.Q (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_7), .QB (
        \$dummy [102]), .D (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .CLK (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_8 (.Q (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_8), .QB (
        \$dummy [103]), .D (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .CLK (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_9 (.Q (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_9), .QB (
        \$dummy [104]), .D (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .CLK (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_10 (.Q (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_10), .QB (
        \$dummy [105]), .D (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .CLK (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_11 (.Q (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_11), .QB (
        \$dummy [106]), .D (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .CLK (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_12 (.Q (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_12), .QB (
        \$dummy [107]), .D (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .CLK (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_13 (.Q (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_13), .QB (
        \$dummy [108]), .D (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .CLK (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_14 (.Q (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_14), .QB (
        \$dummy [109]), .D (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .CLK (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_15 (.Q (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_15), .QB (
        \$dummy [110]), .D (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .CLK (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_16 (.Q (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_16), .QB (
        \$dummy [111]), .D (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .CLK (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    inv02 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix623 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix625 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix627 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix643 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644), .A (
          nx7425)) ;
    dff CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_0 (.Q (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_0), .QB (\$dummy [112]), .D (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .CLK (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    nor02_2x CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix567 (.Y (
             CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566), .A0 (
             RST), .A1 (
             CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    dff CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_1 (.Q (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_1), .QB (\$dummy [113]), .D (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .CLK (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_2 (.Q (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_2), .QB (\$dummy [114]), .D (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .CLK (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_3 (.Q (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_3), .QB (\$dummy [115]), .D (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .CLK (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_4 (.Q (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_4), .QB (\$dummy [116]), .D (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .CLK (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_5 (.Q (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_5), .QB (\$dummy [117]), .D (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .CLK (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_6 (.Q (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_6), .QB (\$dummy [118]), .D (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .CLK (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_7 (.Q (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_7), .QB (\$dummy [119]), .D (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .CLK (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_8 (.Q (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_8), .QB (\$dummy [120]), .D (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .CLK (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_9 (.Q (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_9), .QB (\$dummy [121]), .D (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .CLK (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_10 (.Q (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_10), .QB (\$dummy [122]), .D (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .CLK (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_11 (.Q (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_11), .QB (\$dummy [123]), .D (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .CLK (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_12 (.Q (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_12), .QB (\$dummy [124]), .D (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .CLK (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_13 (.Q (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_13), .QB (\$dummy [125]), .D (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .CLK (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_14 (.Q (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_14), .QB (\$dummy [126]), .D (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .CLK (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_15 (.Q (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_15), .QB (\$dummy [127]), .D (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .CLK (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_16 (.Q (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_16), .QB (\$dummy [128]), .D (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .CLK (
        CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    inv02 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix623 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix625 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix627 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix643 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642)) ;
    xor2 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix83 (.Y (CALCULATOR_L1Results_2__0), 
         .A0 (CALCULATOR_L1SecondOperands_2__0), .A1 (
         CALCULATOR_L1FirstOperands_2__0)) ;
    xnor2 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix380 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx379), .A0 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx381), .A1 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx383)) ;
    nand02 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix382 (.Y (
           CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx381), .A0 (
           CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothOperand_0), .A1 (nx7445)) ;
    xnor2 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix384 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx383), .A0 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothOperand_1), .A1 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_1)) ;
    inv01 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix388 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx387), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_2)) ;
    xnor2 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix390 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx389), .A0 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx391), .A1 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx395)) ;
    aoi32 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix392 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx391), .A0 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothOperand_0), .A1 (nx7445), .A2 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx154), .B0 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_1), .B1 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothOperand_1)) ;
    xnor2 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix396 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx395), .A0 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothOperand_2), .A1 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_2)) ;
    inv01 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix400 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx399), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_3)) ;
    xnor2 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix402 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx401), .A0 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx403), .A1 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx405)) ;
    xnor2 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix406 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx405), .A0 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothOperand_3), .A1 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_3)) ;
    inv01 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix410 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx409), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_4)) ;
    xnor2 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix412 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx411), .A0 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx413), .A1 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx415)) ;
    xnor2 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix416 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx415), .A0 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothOperand_4), .A1 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_4)) ;
    inv01 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix420 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx419), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_5)) ;
    xnor2 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix422 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx421), .A0 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx423), .A1 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx425)) ;
    xnor2 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix426 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx425), .A0 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothOperand_5), .A1 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_5)) ;
    inv01 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix430 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx429), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_6)) ;
    xnor2 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix432 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx431), .A0 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx433), .A1 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx435)) ;
    xnor2 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix436 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx435), .A0 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothOperand_6), .A1 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_6)) ;
    inv01 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix440 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx439), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_7)) ;
    xnor2 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix442 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx441), .A0 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx443), .A1 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx445)) ;
    xnor2 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix446 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx445), .A0 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothOperand_7), .A1 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_7)) ;
    inv01 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix450 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx449), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_8)) ;
    xnor2 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix452 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx451), .A0 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx453), .A1 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx455)) ;
    xnor2 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix456 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx455), .A0 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothOperand_8), .A1 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_8)) ;
    xor2 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix317 (.Y (
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx316), .A0 (
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx461), .A1 (
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx463)) ;
    xnor2 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix464 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx463), .A0 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothOperand_9), .A1 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_9)) ;
    xor2 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix337 (.Y (
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx336), .A0 (
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx467), .A1 (
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx471)) ;
    inv01 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix470 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx469), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_9)) ;
    xnor2 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix472 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx471), .A0 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothOperand_10), .A1 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_10)) ;
    xor2 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix357 (.Y (
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx356), .A0 (
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx475), .A1 (
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx479)) ;
    inv01 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix478 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx477), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_10)) ;
    xnor2 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix480 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx479), .A0 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothOperand_11), .A1 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_11)) ;
    xor2 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix377 (.Y (
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx376), .A0 (
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx483), .A1 (
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx487)) ;
    inv01 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix486 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx485), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_11)) ;
    xnor2 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix488 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx487), .A0 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothOperand_12), .A1 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_12)) ;
    xor2 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix397 (.Y (
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx396), .A0 (
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx491), .A1 (
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx495)) ;
    inv01 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix494 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx493), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_12)) ;
    xnor2 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix496 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx495), .A0 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothOperand_13), .A1 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_13)) ;
    xor2 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix417 (.Y (
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx416), .A0 (
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx499), .A1 (
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx503)) ;
    inv01 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix502 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx501), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_13)) ;
    xnor2 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix504 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx503), .A0 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothOperand_14), .A1 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_14)) ;
    xor2 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix437 (.Y (
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx436), .A0 (
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx507), .A1 (
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx511)) ;
    inv01 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix510 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx509), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_14)) ;
    xnor2 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix512 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx511), .A0 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothOperand_15), .A1 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_15)) ;
    xnor2 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix457 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx456), .A0 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx515), .A1 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx454)) ;
    inv01 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix518 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx517), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_15)) ;
    xor2 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix455 (.Y (
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx454), .A0 (
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothOperand_16), .A1 (
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_16)) ;
    mux21_ni CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix91 (.Y (
             CALCULATOR_L1SecondOperands_2__0), .A0 (
             CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_1), .A1 (
             CacheWindow_0__2__0), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix99 (.Y (
             CALCULATOR_L1SecondOperands_2__1), .A0 (
             CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_2), .A1 (
             CacheWindow_0__2__1), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix107 (.Y (
             CALCULATOR_L1SecondOperands_2__2), .A0 (
             CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_3), .A1 (
             CacheWindow_0__2__2), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix115 (.Y (
             CALCULATOR_L1SecondOperands_2__3), .A0 (
             CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_4), .A1 (
             CacheWindow_0__2__3), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix123 (.Y (
             CALCULATOR_L1SecondOperands_2__4), .A0 (
             CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_5), .A1 (
             CacheWindow_0__2__4), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix131 (.Y (
             CALCULATOR_L1SecondOperands_2__5), .A0 (
             CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_6), .A1 (
             CacheWindow_0__2__5), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix139 (.Y (
             CALCULATOR_L1SecondOperands_2__6), .A0 (
             CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_7), .A1 (
             CacheWindow_0__2__6), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix147 (.Y (
             CALCULATOR_L1SecondOperands_2__7), .A0 (
             CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_8), .A1 (
             CacheWindow_0__2__7), .S0 (Instr)) ;
    xor2 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix77 (.Y (CALCULATOR_L1Results_2__1), 
         .A0 (CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx529), .A1 (
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx531)) ;
    nand02 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix530 (.Y (
           CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx529), .A0 (
           CALCULATOR_L1SecondOperands_2__0), .A1 (
           CALCULATOR_L1FirstOperands_2__0)) ;
    xnor2 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix532 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx531), .A0 (
          CALCULATOR_L1SecondOperands_2__1), .A1 (
          CALCULATOR_L1FirstOperands_2__1)) ;
    xor2 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix75 (.Y (CALCULATOR_L1Results_2__2), 
         .A0 (CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx534), .A1 (
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx537)) ;
    aoi32 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix535 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx534), .A0 (
          CALCULATOR_L1SecondOperands_2__0), .A1 (
          CALCULATOR_L1FirstOperands_2__0), .A2 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx30), .B0 (
          CALCULATOR_L1FirstOperands_2__1), .B1 (
          CALCULATOR_L1SecondOperands_2__1)) ;
    xnor2 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix538 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx537), .A0 (
          CALCULATOR_L1SecondOperands_2__2), .A1 (
          CALCULATOR_L1FirstOperands_2__2)) ;
    xor2 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix73 (.Y (CALCULATOR_L1Results_2__3), 
         .A0 (CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx540), .A1 (
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx544)) ;
    aoi22 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix541 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx540), .A0 (
          CALCULATOR_L1FirstOperands_2__2), .A1 (
          CALCULATOR_L1SecondOperands_2__2), .B0 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx40), .B1 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx24)) ;
    xnor2 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix545 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx544), .A0 (
          CALCULATOR_L1SecondOperands_2__3), .A1 (
          CALCULATOR_L1FirstOperands_2__3)) ;
    xor2 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix71 (.Y (CALCULATOR_L1Results_2__4), 
         .A0 (CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx547), .A1 (
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx551)) ;
    aoi22 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix548 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx547), .A0 (
          CALCULATOR_L1FirstOperands_2__3), .A1 (
          CALCULATOR_L1SecondOperands_2__3), .B0 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx44), .B1 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx18)) ;
    xnor2 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix552 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx551), .A0 (
          CALCULATOR_L1SecondOperands_2__4), .A1 (
          CALCULATOR_L1FirstOperands_2__4)) ;
    xor2 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix69 (.Y (CALCULATOR_L1Results_2__5), 
         .A0 (CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx554), .A1 (
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx558)) ;
    aoi22 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix555 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx554), .A0 (
          CALCULATOR_L1FirstOperands_2__4), .A1 (
          CALCULATOR_L1SecondOperands_2__4), .B0 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx48), .B1 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx12)) ;
    xnor2 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix559 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx558), .A0 (
          CALCULATOR_L1SecondOperands_2__5), .A1 (
          CALCULATOR_L1FirstOperands_2__5)) ;
    xor2 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix67 (.Y (CALCULATOR_L1Results_2__6), 
         .A0 (CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx561), .A1 (
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx565)) ;
    aoi22 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix562 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx561), .A0 (
          CALCULATOR_L1FirstOperands_2__5), .A1 (
          CALCULATOR_L1SecondOperands_2__5), .B0 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx52), .B1 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx6)) ;
    xnor2 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix566 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx565), .A0 (
          CALCULATOR_L1SecondOperands_2__6), .A1 (
          CALCULATOR_L1FirstOperands_2__6)) ;
    xnor2 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix65 (.Y (CALCULATOR_L1Results_2__7)
          , .A0 (CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx568), .A1 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx62)) ;
    aoi22 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix569 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx568), .A0 (
          CALCULATOR_L1FirstOperands_2__6), .A1 (
          CALCULATOR_L1SecondOperands_2__6), .B0 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx56), .B1 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx0)) ;
    xor2 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix63 (.Y (
         CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx62), .A0 (
         CALCULATOR_L1SecondOperands_2__7), .A1 (CALCULATOR_L1FirstOperands_2__7
         )) ;
    inv01 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix155 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx154), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx383)) ;
    inv01 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix57 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx56), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx561)) ;
    inv01 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix53 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx52), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx554)) ;
    inv01 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix49 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx48), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx547)) ;
    inv01 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix45 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx44), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx540)) ;
    inv01 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix41 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx40), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx534)) ;
    inv01 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix31 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx30), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx531)) ;
    inv01 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix25 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx24), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx537)) ;
    inv01 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix19 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx18), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx544)) ;
    inv01 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix13 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx12), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx551)) ;
    inv01 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix7 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx6), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx558)) ;
    inv01 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix1 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx0), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx565)) ;
    fake_gnd CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix216 (.Y (
             CALCULATOR_L1_0_L2_2_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    aoi21 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix77 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_10), .A0 (
          CacheFilter_0__2__1), .A1 (CacheFilter_0__2__0), .B0 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx4)) ;
    nor02_2x CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix5 (.Y (
             CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx4), .A0 (
             CacheFilter_0__2__0), .A1 (CacheFilter_0__2__1)) ;
    aoi21 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix67 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_11), .A0 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx328), .A1 (
          CacheFilter_0__2__2), .B0 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx8)) ;
    nor03_2x CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix9 (.Y (
             CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx8), .A0 (
             CacheFilter_0__2__2), .A1 (CacheFilter_0__2__0), .A2 (
             CacheFilter_0__2__1)) ;
    xnor2 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix59 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_12), .A0 (
          CacheFilter_0__2__3), .A1 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx8)) ;
    xnor2 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix51 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_13), .A0 (
          CacheFilter_0__2__4), .A1 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx12)) ;
    nor04 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix13 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx12), .A0 (
          CacheFilter_0__2__3), .A1 (CacheFilter_0__2__2), .A2 (
          CacheFilter_0__2__0), .A3 (CacheFilter_0__2__1)) ;
    xnor2 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix43 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_14), .A0 (
          CacheFilter_0__2__5), .A1 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx16)) ;
    nor02ii CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix17 (.Y (
            CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx16), .A0 (
            CacheFilter_0__2__4), .A1 (
            CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx12)) ;
    xnor2 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix35 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_15), .A0 (
          CacheFilter_0__2__6), .A1 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx20)) ;
    nor02ii CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix21 (.Y (
            CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx20), .A0 (
            CacheFilter_0__2__5), .A1 (
            CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx16)) ;
    xnor2 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix27 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_16), .A0 (
          CacheFilter_0__2__7), .A1 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx24)) ;
    nor02ii CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix25 (.Y (
            CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx24), .A0 (
            CacheFilter_0__2__6), .A1 (
            CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx20)) ;
    inv01 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix329 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx328), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx4)) ;
    inv02 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix383 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx384), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_0)) ;
    dff CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_0 (.Q (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_0), .QB (
        \$dummy [129]), .D (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .CLK (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    nor02_2x CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix567 (.Y (
             CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566), .A0 (
             RST), .A1 (
             CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644)) ;
    dff CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_1 (.Q (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_1), .QB (
        \$dummy [130]), .D (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .CLK (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_2 (.Q (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_2), .QB (
        \$dummy [131]), .D (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .CLK (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_3 (.Q (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_3), .QB (
        \$dummy [132]), .D (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .CLK (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_4 (.Q (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_4), .QB (
        \$dummy [133]), .D (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .CLK (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_5 (.Q (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_5), .QB (
        \$dummy [134]), .D (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .CLK (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_6 (.Q (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_6), .QB (
        \$dummy [135]), .D (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .CLK (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_7 (.Q (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_7), .QB (
        \$dummy [136]), .D (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .CLK (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_8 (.Q (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_8), .QB (
        \$dummy [137]), .D (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .CLK (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_9 (.Q (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_9), .QB (
        \$dummy [138]), .D (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .CLK (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_10 (.Q (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_10), .QB (
        \$dummy [139]), .D (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .CLK (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_11 (.Q (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_11), .QB (
        \$dummy [140]), .D (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .CLK (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_12 (.Q (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_12), .QB (
        \$dummy [141]), .D (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .CLK (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_13 (.Q (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_13), .QB (
        \$dummy [142]), .D (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .CLK (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_14 (.Q (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_14), .QB (
        \$dummy [143]), .D (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .CLK (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_15 (.Q (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_15), .QB (
        \$dummy [144]), .D (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .CLK (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_16 (.Q (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_16), .QB (
        \$dummy [145]), .D (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .CLK (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    inv02 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix623 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix625 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix627 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix643 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644), .A (
          nx7459)) ;
    dff CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_0 (.Q (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_0), .QB (
        \$dummy [146]), .D (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .CLK (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    nor02_2x CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix567 (.Y (
             CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566), .A0 (
             RST), .A1 (
             CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644)) ;
    dff CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_1 (.Q (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_1), .QB (
        \$dummy [147]), .D (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .CLK (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_2 (.Q (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_2), .QB (
        \$dummy [148]), .D (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .CLK (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_3 (.Q (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_3), .QB (
        \$dummy [149]), .D (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .CLK (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_4 (.Q (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_4), .QB (
        \$dummy [150]), .D (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .CLK (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_5 (.Q (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_5), .QB (
        \$dummy [151]), .D (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .CLK (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_6 (.Q (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_6), .QB (
        \$dummy [152]), .D (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .CLK (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_7 (.Q (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_7), .QB (
        \$dummy [153]), .D (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .CLK (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_8 (.Q (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_8), .QB (
        \$dummy [154]), .D (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .CLK (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_9 (.Q (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_9), .QB (
        \$dummy [155]), .D (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .CLK (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_10 (.Q (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_10), .QB (
        \$dummy [156]), .D (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .CLK (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_11 (.Q (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_11), .QB (
        \$dummy [157]), .D (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .CLK (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_12 (.Q (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_12), .QB (
        \$dummy [158]), .D (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .CLK (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_13 (.Q (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_13), .QB (
        \$dummy [159]), .D (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .CLK (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_14 (.Q (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_14), .QB (
        \$dummy [160]), .D (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .CLK (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_15 (.Q (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_15), .QB (
        \$dummy [161]), .D (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .CLK (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_16 (.Q (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_16), .QB (
        \$dummy [162]), .D (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .CLK (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    inv02 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix623 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix625 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix627 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix643 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644), .A (
          nx7465)) ;
    dff CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_0 (.Q (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_0), .QB (\$dummy [163]), .D (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .CLK (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    nor02_2x CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix567 (.Y (
             CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566), .A0 (
             RST), .A1 (
             CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    dff CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_1 (.Q (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_1), .QB (\$dummy [164]), .D (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .CLK (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_2 (.Q (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_2), .QB (\$dummy [165]), .D (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .CLK (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_3 (.Q (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_3), .QB (\$dummy [166]), .D (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .CLK (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_4 (.Q (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_4), .QB (\$dummy [167]), .D (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .CLK (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_5 (.Q (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_5), .QB (\$dummy [168]), .D (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .CLK (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_6 (.Q (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_6), .QB (\$dummy [169]), .D (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .CLK (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_7 (.Q (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_7), .QB (\$dummy [170]), .D (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .CLK (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_8 (.Q (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_8), .QB (\$dummy [171]), .D (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .CLK (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_9 (.Q (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_9), .QB (\$dummy [172]), .D (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .CLK (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_10 (.Q (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_10), .QB (\$dummy [173]), .D (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .CLK (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_11 (.Q (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_11), .QB (\$dummy [174]), .D (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .CLK (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_12 (.Q (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_12), .QB (\$dummy [175]), .D (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .CLK (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_13 (.Q (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_13), .QB (\$dummy [176]), .D (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .CLK (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_14 (.Q (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_14), .QB (\$dummy [177]), .D (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .CLK (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_15 (.Q (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_15), .QB (\$dummy [178]), .D (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .CLK (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_16 (.Q (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_16), .QB (\$dummy [179]), .D (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .CLK (
        CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    inv02 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix623 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix625 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix627 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix643 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642)) ;
    xor2 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix83 (.Y (CALCULATOR_L1Results_3__0), 
         .A0 (CALCULATOR_L1SecondOperands_3__0), .A1 (
         CALCULATOR_L1FirstOperands_3__0)) ;
    xnor2 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix380 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx379), .A0 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx381), .A1 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx383)) ;
    nand02 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix382 (.Y (
           CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx381), .A0 (
           CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothOperand_0), .A1 (nx7485)) ;
    xnor2 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix384 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx383), .A0 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothOperand_1), .A1 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_1)) ;
    inv01 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix388 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx387), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_2)) ;
    xnor2 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix390 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx389), .A0 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx391), .A1 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx395)) ;
    aoi32 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix392 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx391), .A0 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothOperand_0), .A1 (nx7485), .A2 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx154), .B0 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_1), .B1 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothOperand_1)) ;
    xnor2 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix396 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx395), .A0 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothOperand_2), .A1 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_2)) ;
    inv01 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix400 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx399), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_3)) ;
    xnor2 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix402 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx401), .A0 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx403), .A1 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx405)) ;
    xnor2 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix406 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx405), .A0 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothOperand_3), .A1 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_3)) ;
    inv01 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix410 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx409), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_4)) ;
    xnor2 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix412 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx411), .A0 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx413), .A1 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx415)) ;
    xnor2 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix416 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx415), .A0 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothOperand_4), .A1 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_4)) ;
    inv01 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix420 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx419), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_5)) ;
    xnor2 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix422 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx421), .A0 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx423), .A1 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx425)) ;
    xnor2 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix426 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx425), .A0 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothOperand_5), .A1 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_5)) ;
    inv01 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix430 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx429), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_6)) ;
    xnor2 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix432 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx431), .A0 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx433), .A1 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx435)) ;
    xnor2 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix436 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx435), .A0 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothOperand_6), .A1 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_6)) ;
    inv01 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix440 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx439), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_7)) ;
    xnor2 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix442 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx441), .A0 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx443), .A1 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx445)) ;
    xnor2 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix446 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx445), .A0 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothOperand_7), .A1 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_7)) ;
    inv01 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix450 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx449), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_8)) ;
    xnor2 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix452 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx451), .A0 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx453), .A1 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx455)) ;
    xnor2 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix456 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx455), .A0 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothOperand_8), .A1 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_8)) ;
    xor2 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix317 (.Y (
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx316), .A0 (
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx461), .A1 (
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx463)) ;
    xnor2 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix464 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx463), .A0 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothOperand_9), .A1 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_9)) ;
    xor2 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix337 (.Y (
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx336), .A0 (
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx467), .A1 (
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx471)) ;
    inv01 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix470 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx469), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_9)) ;
    xnor2 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix472 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx471), .A0 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothOperand_10), .A1 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_10)) ;
    xor2 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix357 (.Y (
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx356), .A0 (
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx475), .A1 (
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx479)) ;
    inv01 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix478 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx477), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_10)) ;
    xnor2 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix480 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx479), .A0 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothOperand_11), .A1 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_11)) ;
    xor2 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix377 (.Y (
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx376), .A0 (
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx483), .A1 (
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx487)) ;
    inv01 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix486 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx485), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_11)) ;
    xnor2 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix488 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx487), .A0 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothOperand_12), .A1 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_12)) ;
    xor2 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix397 (.Y (
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx396), .A0 (
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx491), .A1 (
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx495)) ;
    inv01 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix494 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx493), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_12)) ;
    xnor2 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix496 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx495), .A0 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothOperand_13), .A1 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_13)) ;
    xor2 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix417 (.Y (
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx416), .A0 (
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx499), .A1 (
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx503)) ;
    inv01 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix502 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx501), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_13)) ;
    xnor2 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix504 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx503), .A0 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothOperand_14), .A1 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_14)) ;
    xor2 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix437 (.Y (
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx436), .A0 (
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx507), .A1 (
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx511)) ;
    inv01 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix510 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx509), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_14)) ;
    xnor2 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix512 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx511), .A0 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothOperand_15), .A1 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_15)) ;
    xnor2 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix457 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx456), .A0 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx515), .A1 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx454)) ;
    inv01 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix518 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx517), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_15)) ;
    xor2 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix455 (.Y (
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx454), .A0 (
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothOperand_16), .A1 (
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_16)) ;
    mux21_ni CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix91 (.Y (
             CALCULATOR_L1SecondOperands_3__0), .A0 (
             CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_1), .A1 (
             CacheWindow_0__3__0), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix99 (.Y (
             CALCULATOR_L1SecondOperands_3__1), .A0 (
             CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_2), .A1 (
             CacheWindow_0__3__1), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix107 (.Y (
             CALCULATOR_L1SecondOperands_3__2), .A0 (
             CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_3), .A1 (
             CacheWindow_0__3__2), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix115 (.Y (
             CALCULATOR_L1SecondOperands_3__3), .A0 (
             CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_4), .A1 (
             CacheWindow_0__3__3), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix123 (.Y (
             CALCULATOR_L1SecondOperands_3__4), .A0 (
             CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_5), .A1 (
             CacheWindow_0__3__4), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix131 (.Y (
             CALCULATOR_L1SecondOperands_3__5), .A0 (
             CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_6), .A1 (
             CacheWindow_0__3__5), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix139 (.Y (
             CALCULATOR_L1SecondOperands_3__6), .A0 (
             CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_7), .A1 (
             CacheWindow_0__3__6), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix147 (.Y (
             CALCULATOR_L1SecondOperands_3__7), .A0 (
             CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_8), .A1 (
             CacheWindow_0__3__7), .S0 (Instr)) ;
    xor2 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix77 (.Y (CALCULATOR_L1Results_3__1), 
         .A0 (CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx529), .A1 (
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx531)) ;
    nand02 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix530 (.Y (
           CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx529), .A0 (
           CALCULATOR_L1SecondOperands_3__0), .A1 (
           CALCULATOR_L1FirstOperands_3__0)) ;
    xnor2 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix532 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx531), .A0 (
          CALCULATOR_L1SecondOperands_3__1), .A1 (
          CALCULATOR_L1FirstOperands_3__1)) ;
    xor2 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix75 (.Y (CALCULATOR_L1Results_3__2), 
         .A0 (CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx534), .A1 (
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx537)) ;
    aoi32 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix535 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx534), .A0 (
          CALCULATOR_L1SecondOperands_3__0), .A1 (
          CALCULATOR_L1FirstOperands_3__0), .A2 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx30), .B0 (
          CALCULATOR_L1FirstOperands_3__1), .B1 (
          CALCULATOR_L1SecondOperands_3__1)) ;
    xnor2 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix538 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx537), .A0 (
          CALCULATOR_L1SecondOperands_3__2), .A1 (
          CALCULATOR_L1FirstOperands_3__2)) ;
    xor2 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix73 (.Y (CALCULATOR_L1Results_3__3), 
         .A0 (CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx540), .A1 (
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx544)) ;
    aoi22 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix541 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx540), .A0 (
          CALCULATOR_L1FirstOperands_3__2), .A1 (
          CALCULATOR_L1SecondOperands_3__2), .B0 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx40), .B1 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx24)) ;
    xnor2 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix545 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx544), .A0 (
          CALCULATOR_L1SecondOperands_3__3), .A1 (
          CALCULATOR_L1FirstOperands_3__3)) ;
    xor2 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix71 (.Y (CALCULATOR_L1Results_3__4), 
         .A0 (CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx547), .A1 (
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx551)) ;
    aoi22 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix548 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx547), .A0 (
          CALCULATOR_L1FirstOperands_3__3), .A1 (
          CALCULATOR_L1SecondOperands_3__3), .B0 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx44), .B1 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx18)) ;
    xnor2 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix552 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx551), .A0 (
          CALCULATOR_L1SecondOperands_3__4), .A1 (
          CALCULATOR_L1FirstOperands_3__4)) ;
    xor2 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix69 (.Y (CALCULATOR_L1Results_3__5), 
         .A0 (CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx554), .A1 (
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx558)) ;
    aoi22 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix555 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx554), .A0 (
          CALCULATOR_L1FirstOperands_3__4), .A1 (
          CALCULATOR_L1SecondOperands_3__4), .B0 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx48), .B1 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx12)) ;
    xnor2 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix559 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx558), .A0 (
          CALCULATOR_L1SecondOperands_3__5), .A1 (
          CALCULATOR_L1FirstOperands_3__5)) ;
    xor2 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix67 (.Y (CALCULATOR_L1Results_3__6), 
         .A0 (CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx561), .A1 (
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx565)) ;
    aoi22 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix562 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx561), .A0 (
          CALCULATOR_L1FirstOperands_3__5), .A1 (
          CALCULATOR_L1SecondOperands_3__5), .B0 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx52), .B1 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx6)) ;
    xnor2 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix566 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx565), .A0 (
          CALCULATOR_L1SecondOperands_3__6), .A1 (
          CALCULATOR_L1FirstOperands_3__6)) ;
    xnor2 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix65 (.Y (CALCULATOR_L1Results_3__7)
          , .A0 (CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx568), .A1 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx62)) ;
    aoi22 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix569 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx568), .A0 (
          CALCULATOR_L1FirstOperands_3__6), .A1 (
          CALCULATOR_L1SecondOperands_3__6), .B0 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx56), .B1 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx0)) ;
    xor2 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix63 (.Y (
         CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx62), .A0 (
         CALCULATOR_L1SecondOperands_3__7), .A1 (CALCULATOR_L1FirstOperands_3__7
         )) ;
    inv01 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix155 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx154), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx383)) ;
    inv01 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix57 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx56), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx561)) ;
    inv01 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix53 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx52), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx554)) ;
    inv01 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix49 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx48), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx547)) ;
    inv01 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix45 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx44), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx540)) ;
    inv01 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix41 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx40), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx534)) ;
    inv01 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix31 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx30), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx531)) ;
    inv01 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix25 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx24), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx537)) ;
    inv01 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix19 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx18), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx544)) ;
    inv01 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix13 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx12), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx551)) ;
    inv01 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix7 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx6), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx558)) ;
    inv01 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix1 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx0), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx565)) ;
    fake_gnd CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix216 (.Y (
             CALCULATOR_L1_0_L2_3_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    aoi21 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix77 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_10), .A0 (
          CacheFilter_0__3__1), .A1 (CacheFilter_0__3__0), .B0 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx4)) ;
    nor02_2x CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix5 (.Y (
             CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx4), .A0 (
             CacheFilter_0__3__0), .A1 (CacheFilter_0__3__1)) ;
    aoi21 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix67 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_11), .A0 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx328), .A1 (
          CacheFilter_0__3__2), .B0 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx8)) ;
    nor03_2x CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix9 (.Y (
             CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx8), .A0 (
             CacheFilter_0__3__2), .A1 (CacheFilter_0__3__0), .A2 (
             CacheFilter_0__3__1)) ;
    xnor2 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix59 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_12), .A0 (
          CacheFilter_0__3__3), .A1 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx8)) ;
    xnor2 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix51 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_13), .A0 (
          CacheFilter_0__3__4), .A1 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx12)) ;
    nor04 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix13 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx12), .A0 (
          CacheFilter_0__3__3), .A1 (CacheFilter_0__3__2), .A2 (
          CacheFilter_0__3__0), .A3 (CacheFilter_0__3__1)) ;
    xnor2 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix43 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_14), .A0 (
          CacheFilter_0__3__5), .A1 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx16)) ;
    nor02ii CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix17 (.Y (
            CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx16), .A0 (
            CacheFilter_0__3__4), .A1 (
            CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx12)) ;
    xnor2 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix35 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_15), .A0 (
          CacheFilter_0__3__6), .A1 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx20)) ;
    nor02ii CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix21 (.Y (
            CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx20), .A0 (
            CacheFilter_0__3__5), .A1 (
            CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx16)) ;
    xnor2 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix27 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_16), .A0 (
          CacheFilter_0__3__7), .A1 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx24)) ;
    nor02ii CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix25 (.Y (
            CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx24), .A0 (
            CacheFilter_0__3__6), .A1 (
            CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx20)) ;
    inv01 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix329 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx328), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx4)) ;
    inv02 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix383 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx384), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_0)) ;
    dff CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_0 (.Q (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_0), .QB (
        \$dummy [180]), .D (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .CLK (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    nor02_2x CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix567 (.Y (
             CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566), .A0 (
             RST), .A1 (
             CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644)) ;
    dff CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_1 (.Q (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_1), .QB (
        \$dummy [181]), .D (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .CLK (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_2 (.Q (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_2), .QB (
        \$dummy [182]), .D (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .CLK (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_3 (.Q (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_3), .QB (
        \$dummy [183]), .D (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .CLK (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_4 (.Q (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_4), .QB (
        \$dummy [184]), .D (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .CLK (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_5 (.Q (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_5), .QB (
        \$dummy [185]), .D (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .CLK (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_6 (.Q (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_6), .QB (
        \$dummy [186]), .D (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .CLK (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_7 (.Q (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_7), .QB (
        \$dummy [187]), .D (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .CLK (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_8 (.Q (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_8), .QB (
        \$dummy [188]), .D (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .CLK (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_9 (.Q (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_9), .QB (
        \$dummy [189]), .D (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .CLK (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_10 (.Q (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_10), .QB (
        \$dummy [190]), .D (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .CLK (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_11 (.Q (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_11), .QB (
        \$dummy [191]), .D (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .CLK (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_12 (.Q (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_12), .QB (
        \$dummy [192]), .D (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .CLK (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_13 (.Q (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_13), .QB (
        \$dummy [193]), .D (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .CLK (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_14 (.Q (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_14), .QB (
        \$dummy [194]), .D (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .CLK (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_15 (.Q (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_15), .QB (
        \$dummy [195]), .D (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .CLK (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_16 (.Q (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_16), .QB (
        \$dummy [196]), .D (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .CLK (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    inv02 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix623 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix625 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix627 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix643 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644), .A (
          nx7499)) ;
    dff CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_0 (.Q (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_0), .QB (
        \$dummy [197]), .D (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .CLK (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    nor02_2x CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix567 (.Y (
             CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566), .A0 (
             RST), .A1 (
             CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644)) ;
    dff CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_1 (.Q (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_1), .QB (
        \$dummy [198]), .D (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .CLK (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_2 (.Q (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_2), .QB (
        \$dummy [199]), .D (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .CLK (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_3 (.Q (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_3), .QB (
        \$dummy [200]), .D (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .CLK (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_4 (.Q (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_4), .QB (
        \$dummy [201]), .D (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .CLK (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_5 (.Q (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_5), .QB (
        \$dummy [202]), .D (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .CLK (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_6 (.Q (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_6), .QB (
        \$dummy [203]), .D (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .CLK (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_7 (.Q (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_7), .QB (
        \$dummy [204]), .D (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .CLK (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_8 (.Q (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_8), .QB (
        \$dummy [205]), .D (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .CLK (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_9 (.Q (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_9), .QB (
        \$dummy [206]), .D (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .CLK (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_10 (.Q (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_10), .QB (
        \$dummy [207]), .D (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .CLK (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_11 (.Q (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_11), .QB (
        \$dummy [208]), .D (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .CLK (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_12 (.Q (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_12), .QB (
        \$dummy [209]), .D (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .CLK (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_13 (.Q (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_13), .QB (
        \$dummy [210]), .D (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .CLK (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_14 (.Q (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_14), .QB (
        \$dummy [211]), .D (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .CLK (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_15 (.Q (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_15), .QB (
        \$dummy [212]), .D (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .CLK (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_16 (.Q (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_16), .QB (
        \$dummy [213]), .D (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .CLK (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    inv02 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix623 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix625 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix627 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix643 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644), .A (
          nx7505)) ;
    dff CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_0 (.Q (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_0), .QB (\$dummy [214]), .D (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .CLK (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    nor02_2x CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix567 (.Y (
             CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566), .A0 (
             RST), .A1 (
             CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    dff CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_1 (.Q (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_1), .QB (\$dummy [215]), .D (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .CLK (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_2 (.Q (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_2), .QB (\$dummy [216]), .D (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .CLK (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_3 (.Q (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_3), .QB (\$dummy [217]), .D (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .CLK (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_4 (.Q (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_4), .QB (\$dummy [218]), .D (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .CLK (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_5 (.Q (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_5), .QB (\$dummy [219]), .D (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .CLK (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_6 (.Q (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_6), .QB (\$dummy [220]), .D (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .CLK (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_7 (.Q (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_7), .QB (\$dummy [221]), .D (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .CLK (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_8 (.Q (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_8), .QB (\$dummy [222]), .D (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .CLK (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_9 (.Q (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_9), .QB (\$dummy [223]), .D (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .CLK (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_10 (.Q (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_10), .QB (\$dummy [224]), .D (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .CLK (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_11 (.Q (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_11), .QB (\$dummy [225]), .D (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .CLK (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_12 (.Q (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_12), .QB (\$dummy [226]), .D (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .CLK (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_13 (.Q (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_13), .QB (\$dummy [227]), .D (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .CLK (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_14 (.Q (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_14), .QB (\$dummy [228]), .D (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .CLK (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_15 (.Q (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_15), .QB (\$dummy [229]), .D (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .CLK (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_16 (.Q (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_16), .QB (\$dummy [230]), .D (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .CLK (
        CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    inv02 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix623 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix625 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix627 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix643 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642)) ;
    xor2 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix83 (.Y (CALCULATOR_L1Results_4__0), 
         .A0 (CALCULATOR_L1SecondOperands_4__0), .A1 (
         CALCULATOR_L1FirstOperands_4__0)) ;
    xnor2 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix380 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx379), .A0 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx381), .A1 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx383)) ;
    nand02 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix382 (.Y (
           CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx381), .A0 (
           CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothOperand_0), .A1 (nx7525)) ;
    xnor2 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix384 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx383), .A0 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothOperand_1), .A1 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_1)) ;
    inv01 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix388 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx387), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_2)) ;
    xnor2 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix390 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx389), .A0 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx391), .A1 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx395)) ;
    aoi32 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix392 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx391), .A0 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothOperand_0), .A1 (nx7525), .A2 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx154), .B0 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_1), .B1 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothOperand_1)) ;
    xnor2 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix396 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx395), .A0 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothOperand_2), .A1 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_2)) ;
    inv01 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix400 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx399), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_3)) ;
    xnor2 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix402 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx401), .A0 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx403), .A1 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx405)) ;
    xnor2 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix406 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx405), .A0 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothOperand_3), .A1 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_3)) ;
    inv01 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix410 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx409), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_4)) ;
    xnor2 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix412 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx411), .A0 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx413), .A1 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx415)) ;
    xnor2 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix416 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx415), .A0 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothOperand_4), .A1 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_4)) ;
    inv01 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix420 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx419), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_5)) ;
    xnor2 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix422 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx421), .A0 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx423), .A1 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx425)) ;
    xnor2 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix426 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx425), .A0 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothOperand_5), .A1 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_5)) ;
    inv01 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix430 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx429), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_6)) ;
    xnor2 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix432 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx431), .A0 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx433), .A1 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx435)) ;
    xnor2 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix436 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx435), .A0 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothOperand_6), .A1 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_6)) ;
    inv01 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix440 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx439), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_7)) ;
    xnor2 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix442 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx441), .A0 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx443), .A1 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx445)) ;
    xnor2 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix446 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx445), .A0 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothOperand_7), .A1 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_7)) ;
    inv01 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix450 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx449), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_8)) ;
    xnor2 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix452 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx451), .A0 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx453), .A1 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx455)) ;
    xnor2 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix456 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx455), .A0 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothOperand_8), .A1 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_8)) ;
    xor2 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix317 (.Y (
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx316), .A0 (
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx461), .A1 (
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx463)) ;
    xnor2 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix464 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx463), .A0 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothOperand_9), .A1 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_9)) ;
    xor2 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix337 (.Y (
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx336), .A0 (
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx467), .A1 (
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx471)) ;
    inv01 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix470 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx469), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_9)) ;
    xnor2 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix472 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx471), .A0 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothOperand_10), .A1 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_10)) ;
    xor2 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix357 (.Y (
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx356), .A0 (
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx475), .A1 (
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx479)) ;
    inv01 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix478 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx477), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_10)) ;
    xnor2 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix480 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx479), .A0 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothOperand_11), .A1 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_11)) ;
    xor2 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix377 (.Y (
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx376), .A0 (
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx483), .A1 (
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx487)) ;
    inv01 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix486 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx485), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_11)) ;
    xnor2 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix488 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx487), .A0 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothOperand_12), .A1 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_12)) ;
    xor2 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix397 (.Y (
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx396), .A0 (
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx491), .A1 (
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx495)) ;
    inv01 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix494 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx493), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_12)) ;
    xnor2 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix496 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx495), .A0 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothOperand_13), .A1 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_13)) ;
    xor2 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix417 (.Y (
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx416), .A0 (
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx499), .A1 (
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx503)) ;
    inv01 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix502 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx501), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_13)) ;
    xnor2 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix504 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx503), .A0 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothOperand_14), .A1 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_14)) ;
    xor2 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix437 (.Y (
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx436), .A0 (
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx507), .A1 (
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx511)) ;
    inv01 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix510 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx509), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_14)) ;
    xnor2 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix512 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx511), .A0 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothOperand_15), .A1 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_15)) ;
    xnor2 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix457 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx456), .A0 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx515), .A1 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx454)) ;
    inv01 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix518 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx517), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_15)) ;
    xor2 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix455 (.Y (
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx454), .A0 (
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothOperand_16), .A1 (
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_16)) ;
    mux21_ni CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix91 (.Y (
             CALCULATOR_L1SecondOperands_4__0), .A0 (
             CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_1), .A1 (
             CacheWindow_0__4__0), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix99 (.Y (
             CALCULATOR_L1SecondOperands_4__1), .A0 (
             CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_2), .A1 (
             CacheWindow_0__4__1), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix107 (.Y (
             CALCULATOR_L1SecondOperands_4__2), .A0 (
             CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_3), .A1 (
             CacheWindow_0__4__2), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix115 (.Y (
             CALCULATOR_L1SecondOperands_4__3), .A0 (
             CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_4), .A1 (
             CacheWindow_0__4__3), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix123 (.Y (
             CALCULATOR_L1SecondOperands_4__4), .A0 (
             CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_5), .A1 (
             CacheWindow_0__4__4), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix131 (.Y (
             CALCULATOR_L1SecondOperands_4__5), .A0 (
             CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_6), .A1 (
             CacheWindow_0__4__5), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix139 (.Y (
             CALCULATOR_L1SecondOperands_4__6), .A0 (
             CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_7), .A1 (
             CacheWindow_0__4__6), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix147 (.Y (
             CALCULATOR_L1SecondOperands_4__7), .A0 (
             CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_8), .A1 (
             CacheWindow_0__4__7), .S0 (Instr)) ;
    xor2 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix77 (.Y (CALCULATOR_L1Results_4__1), 
         .A0 (CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx529), .A1 (
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx531)) ;
    nand02 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix530 (.Y (
           CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx529), .A0 (
           CALCULATOR_L1SecondOperands_4__0), .A1 (
           CALCULATOR_L1FirstOperands_4__0)) ;
    xnor2 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix532 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx531), .A0 (
          CALCULATOR_L1SecondOperands_4__1), .A1 (
          CALCULATOR_L1FirstOperands_4__1)) ;
    xor2 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix75 (.Y (CALCULATOR_L1Results_4__2), 
         .A0 (CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx534), .A1 (
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx537)) ;
    aoi32 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix535 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx534), .A0 (
          CALCULATOR_L1SecondOperands_4__0), .A1 (
          CALCULATOR_L1FirstOperands_4__0), .A2 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx30), .B0 (
          CALCULATOR_L1FirstOperands_4__1), .B1 (
          CALCULATOR_L1SecondOperands_4__1)) ;
    xnor2 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix538 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx537), .A0 (
          CALCULATOR_L1SecondOperands_4__2), .A1 (
          CALCULATOR_L1FirstOperands_4__2)) ;
    xor2 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix73 (.Y (CALCULATOR_L1Results_4__3), 
         .A0 (CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx540), .A1 (
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx544)) ;
    aoi22 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix541 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx540), .A0 (
          CALCULATOR_L1FirstOperands_4__2), .A1 (
          CALCULATOR_L1SecondOperands_4__2), .B0 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx40), .B1 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx24)) ;
    xnor2 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix545 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx544), .A0 (
          CALCULATOR_L1SecondOperands_4__3), .A1 (
          CALCULATOR_L1FirstOperands_4__3)) ;
    xor2 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix71 (.Y (CALCULATOR_L1Results_4__4), 
         .A0 (CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx547), .A1 (
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx551)) ;
    aoi22 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix548 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx547), .A0 (
          CALCULATOR_L1FirstOperands_4__3), .A1 (
          CALCULATOR_L1SecondOperands_4__3), .B0 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx44), .B1 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx18)) ;
    xnor2 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix552 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx551), .A0 (
          CALCULATOR_L1SecondOperands_4__4), .A1 (
          CALCULATOR_L1FirstOperands_4__4)) ;
    xor2 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix69 (.Y (CALCULATOR_L1Results_4__5), 
         .A0 (CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx554), .A1 (
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx558)) ;
    aoi22 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix555 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx554), .A0 (
          CALCULATOR_L1FirstOperands_4__4), .A1 (
          CALCULATOR_L1SecondOperands_4__4), .B0 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx48), .B1 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx12)) ;
    xnor2 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix559 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx558), .A0 (
          CALCULATOR_L1SecondOperands_4__5), .A1 (
          CALCULATOR_L1FirstOperands_4__5)) ;
    xor2 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix67 (.Y (CALCULATOR_L1Results_4__6), 
         .A0 (CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx561), .A1 (
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx565)) ;
    aoi22 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix562 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx561), .A0 (
          CALCULATOR_L1FirstOperands_4__5), .A1 (
          CALCULATOR_L1SecondOperands_4__5), .B0 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx52), .B1 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx6)) ;
    xnor2 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix566 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx565), .A0 (
          CALCULATOR_L1SecondOperands_4__6), .A1 (
          CALCULATOR_L1FirstOperands_4__6)) ;
    xnor2 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix65 (.Y (CALCULATOR_L1Results_4__7)
          , .A0 (CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx568), .A1 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx62)) ;
    aoi22 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix569 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx568), .A0 (
          CALCULATOR_L1FirstOperands_4__6), .A1 (
          CALCULATOR_L1SecondOperands_4__6), .B0 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx56), .B1 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx0)) ;
    xor2 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix63 (.Y (
         CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx62), .A0 (
         CALCULATOR_L1SecondOperands_4__7), .A1 (CALCULATOR_L1FirstOperands_4__7
         )) ;
    inv01 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix155 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx154), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx383)) ;
    inv01 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix57 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx56), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx561)) ;
    inv01 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix53 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx52), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx554)) ;
    inv01 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix49 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx48), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx547)) ;
    inv01 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix45 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx44), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx540)) ;
    inv01 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix41 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx40), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx534)) ;
    inv01 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix31 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx30), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx531)) ;
    inv01 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix25 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx24), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx537)) ;
    inv01 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix19 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx18), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx544)) ;
    inv01 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix13 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx12), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx551)) ;
    inv01 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix7 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx6), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx558)) ;
    inv01 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix1 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx0), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx565)) ;
    fake_gnd CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix216 (.Y (
             CALCULATOR_L1_0_L2_4_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    aoi21 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix77 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_10), .A0 (
          CacheFilter_0__4__1), .A1 (CacheFilter_0__4__0), .B0 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx4)) ;
    nor02_2x CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix5 (.Y (
             CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx4), .A0 (
             CacheFilter_0__4__0), .A1 (CacheFilter_0__4__1)) ;
    aoi21 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix67 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_11), .A0 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx328), .A1 (
          CacheFilter_0__4__2), .B0 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx8)) ;
    nor03_2x CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix9 (.Y (
             CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx8), .A0 (
             CacheFilter_0__4__2), .A1 (CacheFilter_0__4__0), .A2 (
             CacheFilter_0__4__1)) ;
    xnor2 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix59 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_12), .A0 (
          CacheFilter_0__4__3), .A1 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx8)) ;
    xnor2 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix51 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_13), .A0 (
          CacheFilter_0__4__4), .A1 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx12)) ;
    nor04 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix13 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx12), .A0 (
          CacheFilter_0__4__3), .A1 (CacheFilter_0__4__2), .A2 (
          CacheFilter_0__4__0), .A3 (CacheFilter_0__4__1)) ;
    xnor2 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix43 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_14), .A0 (
          CacheFilter_0__4__5), .A1 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx16)) ;
    nor02ii CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix17 (.Y (
            CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx16), .A0 (
            CacheFilter_0__4__4), .A1 (
            CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx12)) ;
    xnor2 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix35 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_15), .A0 (
          CacheFilter_0__4__6), .A1 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx20)) ;
    nor02ii CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix21 (.Y (
            CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx20), .A0 (
            CacheFilter_0__4__5), .A1 (
            CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx16)) ;
    xnor2 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix27 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_16), .A0 (
          CacheFilter_0__4__7), .A1 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx24)) ;
    nor02ii CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix25 (.Y (
            CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx24), .A0 (
            CacheFilter_0__4__6), .A1 (
            CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx20)) ;
    inv01 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix329 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx328), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx4)) ;
    inv02 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix383 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx384), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_0)) ;
    dff CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_0 (.Q (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_0), .QB (
        \$dummy [231]), .D (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .CLK (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    nor02_2x CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix567 (.Y (
             CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566), .A0 (
             RST), .A1 (
             CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644)) ;
    dff CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_1 (.Q (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_1), .QB (
        \$dummy [232]), .D (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .CLK (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_2 (.Q (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_2), .QB (
        \$dummy [233]), .D (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .CLK (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_3 (.Q (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_3), .QB (
        \$dummy [234]), .D (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .CLK (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_4 (.Q (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_4), .QB (
        \$dummy [235]), .D (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .CLK (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_5 (.Q (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_5), .QB (
        \$dummy [236]), .D (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .CLK (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_6 (.Q (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_6), .QB (
        \$dummy [237]), .D (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .CLK (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_7 (.Q (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_7), .QB (
        \$dummy [238]), .D (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .CLK (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_8 (.Q (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_8), .QB (
        \$dummy [239]), .D (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .CLK (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_9 (.Q (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_9), .QB (
        \$dummy [240]), .D (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .CLK (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_10 (.Q (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_10), .QB (
        \$dummy [241]), .D (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .CLK (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_11 (.Q (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_11), .QB (
        \$dummy [242]), .D (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .CLK (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_12 (.Q (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_12), .QB (
        \$dummy [243]), .D (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .CLK (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_13 (.Q (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_13), .QB (
        \$dummy [244]), .D (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .CLK (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_14 (.Q (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_14), .QB (
        \$dummy [245]), .D (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .CLK (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_15 (.Q (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_15), .QB (
        \$dummy [246]), .D (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .CLK (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_16 (.Q (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_16), .QB (
        \$dummy [247]), .D (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .CLK (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    inv02 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix623 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix625 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix627 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix643 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644), .A (
          nx7539)) ;
    dff CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_0 (.Q (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_0), .QB (
        \$dummy [248]), .D (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .CLK (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    nor02_2x CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix567 (.Y (
             CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566), .A0 (
             RST), .A1 (
             CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644)) ;
    dff CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_1 (.Q (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_1), .QB (
        \$dummy [249]), .D (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .CLK (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_2 (.Q (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_2), .QB (
        \$dummy [250]), .D (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .CLK (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_3 (.Q (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_3), .QB (
        \$dummy [251]), .D (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .CLK (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_4 (.Q (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_4), .QB (
        \$dummy [252]), .D (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .CLK (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_5 (.Q (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_5), .QB (
        \$dummy [253]), .D (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .CLK (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_6 (.Q (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_6), .QB (
        \$dummy [254]), .D (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .CLK (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_7 (.Q (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_7), .QB (
        \$dummy [255]), .D (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .CLK (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_8 (.Q (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_8), .QB (
        \$dummy [256]), .D (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .CLK (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_9 (.Q (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_9), .QB (
        \$dummy [257]), .D (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .CLK (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_10 (.Q (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_10), .QB (
        \$dummy [258]), .D (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .CLK (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_11 (.Q (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_11), .QB (
        \$dummy [259]), .D (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .CLK (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_12 (.Q (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_12), .QB (
        \$dummy [260]), .D (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .CLK (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_13 (.Q (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_13), .QB (
        \$dummy [261]), .D (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .CLK (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_14 (.Q (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_14), .QB (
        \$dummy [262]), .D (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .CLK (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_15 (.Q (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_15), .QB (
        \$dummy [263]), .D (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .CLK (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_16 (.Q (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_16), .QB (
        \$dummy [264]), .D (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .CLK (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    inv02 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix623 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix625 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix627 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix643 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644), .A (
          nx7545)) ;
    dff CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_0 (.Q (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_0), .QB (\$dummy [265]), .D (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .CLK (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    nor02_2x CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix567 (.Y (
             CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566), .A0 (
             RST), .A1 (
             CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    dff CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_1 (.Q (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_1), .QB (\$dummy [266]), .D (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .CLK (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_2 (.Q (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_2), .QB (\$dummy [267]), .D (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .CLK (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_3 (.Q (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_3), .QB (\$dummy [268]), .D (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .CLK (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_4 (.Q (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_4), .QB (\$dummy [269]), .D (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .CLK (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_5 (.Q (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_5), .QB (\$dummy [270]), .D (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .CLK (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_6 (.Q (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_6), .QB (\$dummy [271]), .D (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .CLK (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_7 (.Q (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_7), .QB (\$dummy [272]), .D (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .CLK (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_8 (.Q (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_8), .QB (\$dummy [273]), .D (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .CLK (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_9 (.Q (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_9), .QB (\$dummy [274]), .D (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .CLK (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_10 (.Q (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_10), .QB (\$dummy [275]), .D (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .CLK (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_11 (.Q (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_11), .QB (\$dummy [276]), .D (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .CLK (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_12 (.Q (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_12), .QB (\$dummy [277]), .D (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .CLK (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_13 (.Q (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_13), .QB (\$dummy [278]), .D (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .CLK (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_14 (.Q (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_14), .QB (\$dummy [279]), .D (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .CLK (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_15 (.Q (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_15), .QB (\$dummy [280]), .D (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .CLK (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_16 (.Q (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_16), .QB (\$dummy [281]), .D (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .CLK (
        CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    inv02 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix623 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix625 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix627 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix643 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642)) ;
    xor2 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix83 (.Y (CALCULATOR_L1Results_5__0), 
         .A0 (CALCULATOR_L1SecondOperands_5__0), .A1 (
         CALCULATOR_L1FirstOperands_5__0)) ;
    xnor2 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix380 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx379), .A0 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx381), .A1 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx383)) ;
    nand02 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix382 (.Y (
           CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx381), .A0 (
           CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothOperand_0), .A1 (nx7565)) ;
    xnor2 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix384 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx383), .A0 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothOperand_1), .A1 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_1)) ;
    inv01 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix388 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx387), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_2)) ;
    xnor2 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix390 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx389), .A0 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx391), .A1 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx395)) ;
    aoi32 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix392 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx391), .A0 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothOperand_0), .A1 (nx7565), .A2 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx154), .B0 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_1), .B1 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothOperand_1)) ;
    xnor2 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix396 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx395), .A0 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothOperand_2), .A1 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_2)) ;
    inv01 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix400 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx399), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_3)) ;
    xnor2 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix402 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx401), .A0 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx403), .A1 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx405)) ;
    xnor2 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix406 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx405), .A0 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothOperand_3), .A1 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_3)) ;
    inv01 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix410 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx409), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_4)) ;
    xnor2 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix412 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx411), .A0 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx413), .A1 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx415)) ;
    xnor2 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix416 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx415), .A0 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothOperand_4), .A1 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_4)) ;
    inv01 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix420 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx419), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_5)) ;
    xnor2 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix422 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx421), .A0 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx423), .A1 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx425)) ;
    xnor2 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix426 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx425), .A0 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothOperand_5), .A1 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_5)) ;
    inv01 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix430 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx429), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_6)) ;
    xnor2 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix432 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx431), .A0 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx433), .A1 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx435)) ;
    xnor2 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix436 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx435), .A0 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothOperand_6), .A1 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_6)) ;
    inv01 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix440 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx439), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_7)) ;
    xnor2 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix442 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx441), .A0 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx443), .A1 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx445)) ;
    xnor2 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix446 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx445), .A0 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothOperand_7), .A1 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_7)) ;
    inv01 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix450 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx449), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_8)) ;
    xnor2 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix452 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx451), .A0 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx453), .A1 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx455)) ;
    xnor2 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix456 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx455), .A0 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothOperand_8), .A1 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_8)) ;
    xor2 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix317 (.Y (
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx316), .A0 (
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx461), .A1 (
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx463)) ;
    xnor2 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix464 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx463), .A0 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothOperand_9), .A1 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_9)) ;
    xor2 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix337 (.Y (
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx336), .A0 (
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx467), .A1 (
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx471)) ;
    inv01 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix470 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx469), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_9)) ;
    xnor2 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix472 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx471), .A0 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothOperand_10), .A1 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_10)) ;
    xor2 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix357 (.Y (
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx356), .A0 (
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx475), .A1 (
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx479)) ;
    inv01 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix478 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx477), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_10)) ;
    xnor2 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix480 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx479), .A0 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothOperand_11), .A1 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_11)) ;
    xor2 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix377 (.Y (
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx376), .A0 (
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx483), .A1 (
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx487)) ;
    inv01 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix486 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx485), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_11)) ;
    xnor2 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix488 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx487), .A0 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothOperand_12), .A1 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_12)) ;
    xor2 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix397 (.Y (
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx396), .A0 (
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx491), .A1 (
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx495)) ;
    inv01 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix494 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx493), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_12)) ;
    xnor2 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix496 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx495), .A0 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothOperand_13), .A1 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_13)) ;
    xor2 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix417 (.Y (
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx416), .A0 (
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx499), .A1 (
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx503)) ;
    inv01 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix502 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx501), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_13)) ;
    xnor2 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix504 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx503), .A0 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothOperand_14), .A1 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_14)) ;
    xor2 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix437 (.Y (
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx436), .A0 (
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx507), .A1 (
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx511)) ;
    inv01 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix510 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx509), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_14)) ;
    xnor2 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix512 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx511), .A0 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothOperand_15), .A1 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_15)) ;
    xnor2 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix457 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx456), .A0 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx515), .A1 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx454)) ;
    inv01 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix518 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx517), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_15)) ;
    xor2 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix455 (.Y (
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx454), .A0 (
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothOperand_16), .A1 (
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_16)) ;
    mux21_ni CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix91 (.Y (
             CALCULATOR_L1SecondOperands_5__0), .A0 (
             CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_1), .A1 (
             CacheWindow_1__0__0), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix99 (.Y (
             CALCULATOR_L1SecondOperands_5__1), .A0 (
             CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_2), .A1 (
             CacheWindow_1__0__1), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix107 (.Y (
             CALCULATOR_L1SecondOperands_5__2), .A0 (
             CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_3), .A1 (
             CacheWindow_1__0__2), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix115 (.Y (
             CALCULATOR_L1SecondOperands_5__3), .A0 (
             CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_4), .A1 (
             CacheWindow_1__0__3), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix123 (.Y (
             CALCULATOR_L1SecondOperands_5__4), .A0 (
             CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_5), .A1 (
             CacheWindow_1__0__4), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix131 (.Y (
             CALCULATOR_L1SecondOperands_5__5), .A0 (
             CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_6), .A1 (
             CacheWindow_1__0__5), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix139 (.Y (
             CALCULATOR_L1SecondOperands_5__6), .A0 (
             CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_7), .A1 (
             CacheWindow_1__0__6), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix147 (.Y (
             CALCULATOR_L1SecondOperands_5__7), .A0 (
             CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_8), .A1 (
             CacheWindow_1__0__7), .S0 (Instr)) ;
    xor2 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix77 (.Y (CALCULATOR_L1Results_5__1), 
         .A0 (CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx529), .A1 (
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx531)) ;
    nand02 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix530 (.Y (
           CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx529), .A0 (
           CALCULATOR_L1SecondOperands_5__0), .A1 (
           CALCULATOR_L1FirstOperands_5__0)) ;
    xnor2 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix532 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx531), .A0 (
          CALCULATOR_L1SecondOperands_5__1), .A1 (
          CALCULATOR_L1FirstOperands_5__1)) ;
    xor2 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix75 (.Y (CALCULATOR_L1Results_5__2), 
         .A0 (CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx534), .A1 (
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx537)) ;
    aoi32 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix535 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx534), .A0 (
          CALCULATOR_L1SecondOperands_5__0), .A1 (
          CALCULATOR_L1FirstOperands_5__0), .A2 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx30), .B0 (
          CALCULATOR_L1FirstOperands_5__1), .B1 (
          CALCULATOR_L1SecondOperands_5__1)) ;
    xnor2 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix538 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx537), .A0 (
          CALCULATOR_L1SecondOperands_5__2), .A1 (
          CALCULATOR_L1FirstOperands_5__2)) ;
    xor2 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix73 (.Y (CALCULATOR_L1Results_5__3), 
         .A0 (CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx540), .A1 (
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx544)) ;
    aoi22 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix541 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx540), .A0 (
          CALCULATOR_L1FirstOperands_5__2), .A1 (
          CALCULATOR_L1SecondOperands_5__2), .B0 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx40), .B1 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx24)) ;
    xnor2 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix545 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx544), .A0 (
          CALCULATOR_L1SecondOperands_5__3), .A1 (
          CALCULATOR_L1FirstOperands_5__3)) ;
    xor2 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix71 (.Y (CALCULATOR_L1Results_5__4), 
         .A0 (CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx547), .A1 (
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx551)) ;
    aoi22 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix548 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx547), .A0 (
          CALCULATOR_L1FirstOperands_5__3), .A1 (
          CALCULATOR_L1SecondOperands_5__3), .B0 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx44), .B1 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx18)) ;
    xnor2 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix552 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx551), .A0 (
          CALCULATOR_L1SecondOperands_5__4), .A1 (
          CALCULATOR_L1FirstOperands_5__4)) ;
    xor2 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix69 (.Y (CALCULATOR_L1Results_5__5), 
         .A0 (CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx554), .A1 (
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx558)) ;
    aoi22 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix555 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx554), .A0 (
          CALCULATOR_L1FirstOperands_5__4), .A1 (
          CALCULATOR_L1SecondOperands_5__4), .B0 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx48), .B1 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx12)) ;
    xnor2 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix559 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx558), .A0 (
          CALCULATOR_L1SecondOperands_5__5), .A1 (
          CALCULATOR_L1FirstOperands_5__5)) ;
    xor2 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix67 (.Y (CALCULATOR_L1Results_5__6), 
         .A0 (CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx561), .A1 (
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx565)) ;
    aoi22 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix562 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx561), .A0 (
          CALCULATOR_L1FirstOperands_5__5), .A1 (
          CALCULATOR_L1SecondOperands_5__5), .B0 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx52), .B1 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx6)) ;
    xnor2 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix566 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx565), .A0 (
          CALCULATOR_L1SecondOperands_5__6), .A1 (
          CALCULATOR_L1FirstOperands_5__6)) ;
    xnor2 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix65 (.Y (CALCULATOR_L1Results_5__7)
          , .A0 (CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx568), .A1 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx62)) ;
    aoi22 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix569 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx568), .A0 (
          CALCULATOR_L1FirstOperands_5__6), .A1 (
          CALCULATOR_L1SecondOperands_5__6), .B0 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx56), .B1 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx0)) ;
    xor2 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix63 (.Y (
         CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx62), .A0 (
         CALCULATOR_L1SecondOperands_5__7), .A1 (CALCULATOR_L1FirstOperands_5__7
         )) ;
    inv01 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix155 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx154), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx383)) ;
    inv01 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix57 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx56), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx561)) ;
    inv01 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix53 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx52), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx554)) ;
    inv01 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix49 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx48), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx547)) ;
    inv01 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix45 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx44), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx540)) ;
    inv01 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix41 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx40), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx534)) ;
    inv01 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix31 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx30), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx531)) ;
    inv01 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix25 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx24), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx537)) ;
    inv01 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix19 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx18), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx544)) ;
    inv01 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix13 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx12), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx551)) ;
    inv01 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix7 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx6), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx558)) ;
    inv01 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix1 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx0), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx565)) ;
    fake_gnd CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix216 (.Y (
             CALCULATOR_L1_1_L2_0_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    aoi21 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix77 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_10), .A0 (
          CacheFilter_1__0__1), .A1 (CacheFilter_1__0__0), .B0 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx4)) ;
    nor02_2x CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix5 (.Y (
             CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx4), .A0 (
             CacheFilter_1__0__0), .A1 (CacheFilter_1__0__1)) ;
    aoi21 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix67 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_11), .A0 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx328), .A1 (
          CacheFilter_1__0__2), .B0 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx8)) ;
    nor03_2x CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix9 (.Y (
             CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx8), .A0 (
             CacheFilter_1__0__2), .A1 (CacheFilter_1__0__0), .A2 (
             CacheFilter_1__0__1)) ;
    xnor2 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix59 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_12), .A0 (
          CacheFilter_1__0__3), .A1 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx8)) ;
    xnor2 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix51 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_13), .A0 (
          CacheFilter_1__0__4), .A1 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx12)) ;
    nor04 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix13 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx12), .A0 (
          CacheFilter_1__0__3), .A1 (CacheFilter_1__0__2), .A2 (
          CacheFilter_1__0__0), .A3 (CacheFilter_1__0__1)) ;
    xnor2 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix43 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_14), .A0 (
          CacheFilter_1__0__5), .A1 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx16)) ;
    nor02ii CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix17 (.Y (
            CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx16), .A0 (
            CacheFilter_1__0__4), .A1 (
            CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx12)) ;
    xnor2 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix35 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_15), .A0 (
          CacheFilter_1__0__6), .A1 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx20)) ;
    nor02ii CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix21 (.Y (
            CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx20), .A0 (
            CacheFilter_1__0__5), .A1 (
            CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx16)) ;
    xnor2 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix27 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_16), .A0 (
          CacheFilter_1__0__7), .A1 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx24)) ;
    nor02ii CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix25 (.Y (
            CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx24), .A0 (
            CacheFilter_1__0__6), .A1 (
            CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx20)) ;
    inv01 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix329 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx328), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx4)) ;
    inv02 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix383 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx384), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_0)) ;
    dff CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_0 (.Q (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_0), .QB (
        \$dummy [282]), .D (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .CLK (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    nor02_2x CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix567 (.Y (
             CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566), .A0 (
             RST), .A1 (
             CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644)) ;
    dff CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_1 (.Q (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_1), .QB (
        \$dummy [283]), .D (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .CLK (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_2 (.Q (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_2), .QB (
        \$dummy [284]), .D (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .CLK (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_3 (.Q (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_3), .QB (
        \$dummy [285]), .D (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .CLK (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_4 (.Q (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_4), .QB (
        \$dummy [286]), .D (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .CLK (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_5 (.Q (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_5), .QB (
        \$dummy [287]), .D (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .CLK (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_6 (.Q (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_6), .QB (
        \$dummy [288]), .D (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .CLK (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_7 (.Q (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_7), .QB (
        \$dummy [289]), .D (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .CLK (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_8 (.Q (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_8), .QB (
        \$dummy [290]), .D (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .CLK (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_9 (.Q (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_9), .QB (
        \$dummy [291]), .D (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .CLK (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_10 (.Q (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_10), .QB (
        \$dummy [292]), .D (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .CLK (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_11 (.Q (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_11), .QB (
        \$dummy [293]), .D (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .CLK (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_12 (.Q (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_12), .QB (
        \$dummy [294]), .D (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .CLK (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_13 (.Q (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_13), .QB (
        \$dummy [295]), .D (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .CLK (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_14 (.Q (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_14), .QB (
        \$dummy [296]), .D (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .CLK (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_15 (.Q (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_15), .QB (
        \$dummy [297]), .D (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .CLK (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_16 (.Q (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_16), .QB (
        \$dummy [298]), .D (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .CLK (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    inv02 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix623 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix625 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix627 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix643 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644), .A (
          nx7579)) ;
    dff CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_0 (.Q (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_0), .QB (
        \$dummy [299]), .D (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .CLK (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    nor02_2x CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix567 (.Y (
             CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566), .A0 (
             RST), .A1 (
             CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644)) ;
    dff CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_1 (.Q (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_1), .QB (
        \$dummy [300]), .D (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .CLK (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_2 (.Q (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_2), .QB (
        \$dummy [301]), .D (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .CLK (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_3 (.Q (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_3), .QB (
        \$dummy [302]), .D (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .CLK (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_4 (.Q (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_4), .QB (
        \$dummy [303]), .D (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .CLK (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_5 (.Q (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_5), .QB (
        \$dummy [304]), .D (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .CLK (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_6 (.Q (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_6), .QB (
        \$dummy [305]), .D (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .CLK (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_7 (.Q (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_7), .QB (
        \$dummy [306]), .D (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .CLK (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_8 (.Q (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_8), .QB (
        \$dummy [307]), .D (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .CLK (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_9 (.Q (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_9), .QB (
        \$dummy [308]), .D (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .CLK (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_10 (.Q (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_10), .QB (
        \$dummy [309]), .D (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .CLK (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_11 (.Q (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_11), .QB (
        \$dummy [310]), .D (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .CLK (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_12 (.Q (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_12), .QB (
        \$dummy [311]), .D (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .CLK (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_13 (.Q (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_13), .QB (
        \$dummy [312]), .D (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .CLK (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_14 (.Q (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_14), .QB (
        \$dummy [313]), .D (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .CLK (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_15 (.Q (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_15), .QB (
        \$dummy [314]), .D (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .CLK (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_16 (.Q (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_16), .QB (
        \$dummy [315]), .D (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .CLK (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    inv02 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix623 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix625 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix627 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix643 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644), .A (
          nx7585)) ;
    dff CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_0 (.Q (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_0), .QB (\$dummy [316]), .D (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .CLK (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    nor02_2x CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix567 (.Y (
             CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566), .A0 (
             RST), .A1 (
             CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    dff CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_1 (.Q (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_1), .QB (\$dummy [317]), .D (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .CLK (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_2 (.Q (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_2), .QB (\$dummy [318]), .D (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .CLK (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_3 (.Q (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_3), .QB (\$dummy [319]), .D (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .CLK (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_4 (.Q (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_4), .QB (\$dummy [320]), .D (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .CLK (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_5 (.Q (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_5), .QB (\$dummy [321]), .D (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .CLK (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_6 (.Q (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_6), .QB (\$dummy [322]), .D (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .CLK (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_7 (.Q (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_7), .QB (\$dummy [323]), .D (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .CLK (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_8 (.Q (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_8), .QB (\$dummy [324]), .D (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .CLK (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_9 (.Q (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_9), .QB (\$dummy [325]), .D (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .CLK (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_10 (.Q (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_10), .QB (\$dummy [326]), .D (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .CLK (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_11 (.Q (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_11), .QB (\$dummy [327]), .D (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .CLK (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_12 (.Q (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_12), .QB (\$dummy [328]), .D (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .CLK (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_13 (.Q (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_13), .QB (\$dummy [329]), .D (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .CLK (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_14 (.Q (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_14), .QB (\$dummy [330]), .D (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .CLK (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_15 (.Q (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_15), .QB (\$dummy [331]), .D (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .CLK (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_16 (.Q (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_16), .QB (\$dummy [332]), .D (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .CLK (
        CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    inv02 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix623 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix625 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix627 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix643 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642)) ;
    xor2 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix83 (.Y (CALCULATOR_L1Results_6__0), 
         .A0 (CALCULATOR_L1SecondOperands_6__0), .A1 (
         CALCULATOR_L1FirstOperands_6__0)) ;
    xnor2 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix380 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx379), .A0 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx381), .A1 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx383)) ;
    nand02 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix382 (.Y (
           CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx381), .A0 (
           CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothOperand_0), .A1 (nx7605)) ;
    xnor2 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix384 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx383), .A0 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothOperand_1), .A1 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_1)) ;
    inv01 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix388 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx387), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_2)) ;
    xnor2 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix390 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx389), .A0 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx391), .A1 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx395)) ;
    aoi32 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix392 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx391), .A0 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothOperand_0), .A1 (nx7605), .A2 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx154), .B0 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_1), .B1 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothOperand_1)) ;
    xnor2 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix396 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx395), .A0 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothOperand_2), .A1 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_2)) ;
    inv01 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix400 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx399), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_3)) ;
    xnor2 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix402 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx401), .A0 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx403), .A1 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx405)) ;
    xnor2 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix406 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx405), .A0 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothOperand_3), .A1 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_3)) ;
    inv01 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix410 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx409), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_4)) ;
    xnor2 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix412 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx411), .A0 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx413), .A1 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx415)) ;
    xnor2 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix416 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx415), .A0 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothOperand_4), .A1 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_4)) ;
    inv01 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix420 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx419), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_5)) ;
    xnor2 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix422 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx421), .A0 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx423), .A1 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx425)) ;
    xnor2 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix426 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx425), .A0 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothOperand_5), .A1 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_5)) ;
    inv01 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix430 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx429), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_6)) ;
    xnor2 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix432 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx431), .A0 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx433), .A1 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx435)) ;
    xnor2 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix436 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx435), .A0 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothOperand_6), .A1 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_6)) ;
    inv01 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix440 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx439), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_7)) ;
    xnor2 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix442 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx441), .A0 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx443), .A1 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx445)) ;
    xnor2 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix446 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx445), .A0 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothOperand_7), .A1 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_7)) ;
    inv01 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix450 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx449), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_8)) ;
    xnor2 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix452 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx451), .A0 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx453), .A1 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx455)) ;
    xnor2 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix456 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx455), .A0 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothOperand_8), .A1 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_8)) ;
    xor2 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix317 (.Y (
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx316), .A0 (
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx461), .A1 (
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx463)) ;
    xnor2 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix464 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx463), .A0 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothOperand_9), .A1 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_9)) ;
    xor2 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix337 (.Y (
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx336), .A0 (
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx467), .A1 (
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx471)) ;
    inv01 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix470 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx469), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_9)) ;
    xnor2 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix472 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx471), .A0 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothOperand_10), .A1 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_10)) ;
    xor2 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix357 (.Y (
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx356), .A0 (
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx475), .A1 (
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx479)) ;
    inv01 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix478 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx477), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_10)) ;
    xnor2 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix480 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx479), .A0 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothOperand_11), .A1 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_11)) ;
    xor2 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix377 (.Y (
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx376), .A0 (
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx483), .A1 (
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx487)) ;
    inv01 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix486 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx485), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_11)) ;
    xnor2 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix488 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx487), .A0 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothOperand_12), .A1 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_12)) ;
    xor2 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix397 (.Y (
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx396), .A0 (
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx491), .A1 (
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx495)) ;
    inv01 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix494 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx493), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_12)) ;
    xnor2 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix496 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx495), .A0 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothOperand_13), .A1 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_13)) ;
    xor2 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix417 (.Y (
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx416), .A0 (
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx499), .A1 (
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx503)) ;
    inv01 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix502 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx501), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_13)) ;
    xnor2 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix504 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx503), .A0 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothOperand_14), .A1 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_14)) ;
    xor2 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix437 (.Y (
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx436), .A0 (
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx507), .A1 (
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx511)) ;
    inv01 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix510 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx509), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_14)) ;
    xnor2 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix512 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx511), .A0 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothOperand_15), .A1 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_15)) ;
    xnor2 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix457 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx456), .A0 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx515), .A1 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx454)) ;
    inv01 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix518 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx517), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_15)) ;
    xor2 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix455 (.Y (
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx454), .A0 (
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothOperand_16), .A1 (
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_16)) ;
    mux21_ni CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix91 (.Y (
             CALCULATOR_L1SecondOperands_6__0), .A0 (
             CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_1), .A1 (
             CacheWindow_1__1__0), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix99 (.Y (
             CALCULATOR_L1SecondOperands_6__1), .A0 (
             CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_2), .A1 (
             CacheWindow_1__1__1), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix107 (.Y (
             CALCULATOR_L1SecondOperands_6__2), .A0 (
             CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_3), .A1 (
             CacheWindow_1__1__2), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix115 (.Y (
             CALCULATOR_L1SecondOperands_6__3), .A0 (
             CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_4), .A1 (
             CacheWindow_1__1__3), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix123 (.Y (
             CALCULATOR_L1SecondOperands_6__4), .A0 (
             CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_5), .A1 (
             CacheWindow_1__1__4), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix131 (.Y (
             CALCULATOR_L1SecondOperands_6__5), .A0 (
             CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_6), .A1 (
             CacheWindow_1__1__5), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix139 (.Y (
             CALCULATOR_L1SecondOperands_6__6), .A0 (
             CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_7), .A1 (
             CacheWindow_1__1__6), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix147 (.Y (
             CALCULATOR_L1SecondOperands_6__7), .A0 (
             CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_8), .A1 (
             CacheWindow_1__1__7), .S0 (Instr)) ;
    xor2 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix77 (.Y (CALCULATOR_L1Results_6__1), 
         .A0 (CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx529), .A1 (
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx531)) ;
    nand02 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix530 (.Y (
           CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx529), .A0 (
           CALCULATOR_L1SecondOperands_6__0), .A1 (
           CALCULATOR_L1FirstOperands_6__0)) ;
    xnor2 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix532 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx531), .A0 (
          CALCULATOR_L1SecondOperands_6__1), .A1 (
          CALCULATOR_L1FirstOperands_6__1)) ;
    xor2 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix75 (.Y (CALCULATOR_L1Results_6__2), 
         .A0 (CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx534), .A1 (
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx537)) ;
    aoi32 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix535 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx534), .A0 (
          CALCULATOR_L1SecondOperands_6__0), .A1 (
          CALCULATOR_L1FirstOperands_6__0), .A2 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx30), .B0 (
          CALCULATOR_L1FirstOperands_6__1), .B1 (
          CALCULATOR_L1SecondOperands_6__1)) ;
    xnor2 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix538 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx537), .A0 (
          CALCULATOR_L1SecondOperands_6__2), .A1 (
          CALCULATOR_L1FirstOperands_6__2)) ;
    xor2 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix73 (.Y (CALCULATOR_L1Results_6__3), 
         .A0 (CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx540), .A1 (
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx544)) ;
    aoi22 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix541 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx540), .A0 (
          CALCULATOR_L1FirstOperands_6__2), .A1 (
          CALCULATOR_L1SecondOperands_6__2), .B0 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx40), .B1 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx24)) ;
    xnor2 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix545 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx544), .A0 (
          CALCULATOR_L1SecondOperands_6__3), .A1 (
          CALCULATOR_L1FirstOperands_6__3)) ;
    xor2 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix71 (.Y (CALCULATOR_L1Results_6__4), 
         .A0 (CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx547), .A1 (
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx551)) ;
    aoi22 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix548 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx547), .A0 (
          CALCULATOR_L1FirstOperands_6__3), .A1 (
          CALCULATOR_L1SecondOperands_6__3), .B0 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx44), .B1 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx18)) ;
    xnor2 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix552 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx551), .A0 (
          CALCULATOR_L1SecondOperands_6__4), .A1 (
          CALCULATOR_L1FirstOperands_6__4)) ;
    xor2 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix69 (.Y (CALCULATOR_L1Results_6__5), 
         .A0 (CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx554), .A1 (
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx558)) ;
    aoi22 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix555 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx554), .A0 (
          CALCULATOR_L1FirstOperands_6__4), .A1 (
          CALCULATOR_L1SecondOperands_6__4), .B0 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx48), .B1 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx12)) ;
    xnor2 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix559 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx558), .A0 (
          CALCULATOR_L1SecondOperands_6__5), .A1 (
          CALCULATOR_L1FirstOperands_6__5)) ;
    xor2 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix67 (.Y (CALCULATOR_L1Results_6__6), 
         .A0 (CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx561), .A1 (
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx565)) ;
    aoi22 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix562 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx561), .A0 (
          CALCULATOR_L1FirstOperands_6__5), .A1 (
          CALCULATOR_L1SecondOperands_6__5), .B0 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx52), .B1 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx6)) ;
    xnor2 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix566 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx565), .A0 (
          CALCULATOR_L1SecondOperands_6__6), .A1 (
          CALCULATOR_L1FirstOperands_6__6)) ;
    xnor2 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix65 (.Y (CALCULATOR_L1Results_6__7)
          , .A0 (CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx568), .A1 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx62)) ;
    aoi22 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix569 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx568), .A0 (
          CALCULATOR_L1FirstOperands_6__6), .A1 (
          CALCULATOR_L1SecondOperands_6__6), .B0 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx56), .B1 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx0)) ;
    xor2 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix63 (.Y (
         CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx62), .A0 (
         CALCULATOR_L1SecondOperands_6__7), .A1 (CALCULATOR_L1FirstOperands_6__7
         )) ;
    inv01 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix155 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx154), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx383)) ;
    inv01 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix57 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx56), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx561)) ;
    inv01 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix53 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx52), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx554)) ;
    inv01 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix49 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx48), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx547)) ;
    inv01 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix45 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx44), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx540)) ;
    inv01 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix41 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx40), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx534)) ;
    inv01 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix31 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx30), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx531)) ;
    inv01 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix25 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx24), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx537)) ;
    inv01 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix19 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx18), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx544)) ;
    inv01 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix13 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx12), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx551)) ;
    inv01 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix7 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx6), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx558)) ;
    inv01 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix1 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx0), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx565)) ;
    fake_gnd CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix216 (.Y (
             CALCULATOR_L1_1_L2_1_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    aoi21 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix77 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_10), .A0 (
          CacheFilter_1__1__1), .A1 (CacheFilter_1__1__0), .B0 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx4)) ;
    nor02_2x CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix5 (.Y (
             CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx4), .A0 (
             CacheFilter_1__1__0), .A1 (CacheFilter_1__1__1)) ;
    aoi21 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix67 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_11), .A0 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx328), .A1 (
          CacheFilter_1__1__2), .B0 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx8)) ;
    nor03_2x CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix9 (.Y (
             CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx8), .A0 (
             CacheFilter_1__1__2), .A1 (CacheFilter_1__1__0), .A2 (
             CacheFilter_1__1__1)) ;
    xnor2 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix59 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_12), .A0 (
          CacheFilter_1__1__3), .A1 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx8)) ;
    xnor2 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix51 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_13), .A0 (
          CacheFilter_1__1__4), .A1 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx12)) ;
    nor04 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix13 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx12), .A0 (
          CacheFilter_1__1__3), .A1 (CacheFilter_1__1__2), .A2 (
          CacheFilter_1__1__0), .A3 (CacheFilter_1__1__1)) ;
    xnor2 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix43 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_14), .A0 (
          CacheFilter_1__1__5), .A1 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx16)) ;
    nor02ii CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix17 (.Y (
            CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx16), .A0 (
            CacheFilter_1__1__4), .A1 (
            CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx12)) ;
    xnor2 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix35 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_15), .A0 (
          CacheFilter_1__1__6), .A1 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx20)) ;
    nor02ii CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix21 (.Y (
            CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx20), .A0 (
            CacheFilter_1__1__5), .A1 (
            CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx16)) ;
    xnor2 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix27 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_16), .A0 (
          CacheFilter_1__1__7), .A1 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx24)) ;
    nor02ii CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix25 (.Y (
            CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx24), .A0 (
            CacheFilter_1__1__6), .A1 (
            CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx20)) ;
    inv01 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix329 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx328), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx4)) ;
    inv02 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix383 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx384), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_0)) ;
    dff CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_0 (.Q (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_0), .QB (
        \$dummy [333]), .D (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .CLK (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    nor02_2x CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix567 (.Y (
             CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566), .A0 (
             RST), .A1 (
             CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644)) ;
    dff CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_1 (.Q (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_1), .QB (
        \$dummy [334]), .D (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .CLK (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_2 (.Q (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_2), .QB (
        \$dummy [335]), .D (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .CLK (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_3 (.Q (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_3), .QB (
        \$dummy [336]), .D (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .CLK (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_4 (.Q (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_4), .QB (
        \$dummy [337]), .D (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .CLK (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_5 (.Q (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_5), .QB (
        \$dummy [338]), .D (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .CLK (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_6 (.Q (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_6), .QB (
        \$dummy [339]), .D (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .CLK (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_7 (.Q (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_7), .QB (
        \$dummy [340]), .D (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .CLK (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_8 (.Q (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_8), .QB (
        \$dummy [341]), .D (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .CLK (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_9 (.Q (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_9), .QB (
        \$dummy [342]), .D (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .CLK (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_10 (.Q (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_10), .QB (
        \$dummy [343]), .D (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .CLK (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_11 (.Q (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_11), .QB (
        \$dummy [344]), .D (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .CLK (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_12 (.Q (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_12), .QB (
        \$dummy [345]), .D (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .CLK (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_13 (.Q (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_13), .QB (
        \$dummy [346]), .D (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .CLK (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_14 (.Q (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_14), .QB (
        \$dummy [347]), .D (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .CLK (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_15 (.Q (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_15), .QB (
        \$dummy [348]), .D (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .CLK (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_16 (.Q (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_16), .QB (
        \$dummy [349]), .D (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .CLK (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    inv02 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix623 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix625 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix627 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix643 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644), .A (
          nx7619)) ;
    dff CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_0 (.Q (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_0), .QB (
        \$dummy [350]), .D (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .CLK (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    nor02_2x CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix567 (.Y (
             CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566), .A0 (
             RST), .A1 (
             CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644)) ;
    dff CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_1 (.Q (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_1), .QB (
        \$dummy [351]), .D (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .CLK (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_2 (.Q (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_2), .QB (
        \$dummy [352]), .D (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .CLK (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_3 (.Q (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_3), .QB (
        \$dummy [353]), .D (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .CLK (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_4 (.Q (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_4), .QB (
        \$dummy [354]), .D (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .CLK (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_5 (.Q (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_5), .QB (
        \$dummy [355]), .D (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .CLK (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_6 (.Q (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_6), .QB (
        \$dummy [356]), .D (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .CLK (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_7 (.Q (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_7), .QB (
        \$dummy [357]), .D (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .CLK (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_8 (.Q (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_8), .QB (
        \$dummy [358]), .D (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .CLK (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_9 (.Q (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_9), .QB (
        \$dummy [359]), .D (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .CLK (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_10 (.Q (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_10), .QB (
        \$dummy [360]), .D (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .CLK (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_11 (.Q (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_11), .QB (
        \$dummy [361]), .D (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .CLK (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_12 (.Q (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_12), .QB (
        \$dummy [362]), .D (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .CLK (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_13 (.Q (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_13), .QB (
        \$dummy [363]), .D (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .CLK (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_14 (.Q (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_14), .QB (
        \$dummy [364]), .D (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .CLK (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_15 (.Q (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_15), .QB (
        \$dummy [365]), .D (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .CLK (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_16 (.Q (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_16), .QB (
        \$dummy [366]), .D (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .CLK (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    inv02 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix623 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix625 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix627 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix643 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644), .A (
          nx7625)) ;
    dff CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_0 (.Q (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_0), .QB (\$dummy [367]), .D (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .CLK (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    nor02_2x CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix567 (.Y (
             CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566), .A0 (
             RST), .A1 (
             CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    dff CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_1 (.Q (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_1), .QB (\$dummy [368]), .D (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .CLK (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_2 (.Q (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_2), .QB (\$dummy [369]), .D (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .CLK (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_3 (.Q (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_3), .QB (\$dummy [370]), .D (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .CLK (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_4 (.Q (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_4), .QB (\$dummy [371]), .D (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .CLK (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_5 (.Q (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_5), .QB (\$dummy [372]), .D (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .CLK (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_6 (.Q (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_6), .QB (\$dummy [373]), .D (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .CLK (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_7 (.Q (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_7), .QB (\$dummy [374]), .D (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .CLK (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_8 (.Q (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_8), .QB (\$dummy [375]), .D (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .CLK (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_9 (.Q (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_9), .QB (\$dummy [376]), .D (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .CLK (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_10 (.Q (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_10), .QB (\$dummy [377]), .D (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .CLK (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_11 (.Q (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_11), .QB (\$dummy [378]), .D (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .CLK (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_12 (.Q (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_12), .QB (\$dummy [379]), .D (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .CLK (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_13 (.Q (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_13), .QB (\$dummy [380]), .D (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .CLK (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_14 (.Q (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_14), .QB (\$dummy [381]), .D (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .CLK (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_15 (.Q (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_15), .QB (\$dummy [382]), .D (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .CLK (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_16 (.Q (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_16), .QB (\$dummy [383]), .D (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .CLK (
        CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    inv02 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix623 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix625 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix627 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix643 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642)) ;
    xor2 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix83 (.Y (CALCULATOR_L1Results_7__0), 
         .A0 (CALCULATOR_L1SecondOperands_7__0), .A1 (
         CALCULATOR_L1FirstOperands_7__0)) ;
    xnor2 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix380 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx379), .A0 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx381), .A1 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx383)) ;
    nand02 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix382 (.Y (
           CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx381), .A0 (
           CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothOperand_0), .A1 (nx7645)) ;
    xnor2 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix384 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx383), .A0 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothOperand_1), .A1 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_1)) ;
    inv01 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix388 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx387), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_2)) ;
    xnor2 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix390 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx389), .A0 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx391), .A1 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx395)) ;
    aoi32 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix392 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx391), .A0 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothOperand_0), .A1 (nx7645), .A2 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx154), .B0 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_1), .B1 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothOperand_1)) ;
    xnor2 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix396 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx395), .A0 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothOperand_2), .A1 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_2)) ;
    inv01 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix400 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx399), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_3)) ;
    xnor2 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix402 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx401), .A0 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx403), .A1 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx405)) ;
    xnor2 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix406 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx405), .A0 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothOperand_3), .A1 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_3)) ;
    inv01 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix410 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx409), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_4)) ;
    xnor2 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix412 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx411), .A0 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx413), .A1 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx415)) ;
    xnor2 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix416 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx415), .A0 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothOperand_4), .A1 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_4)) ;
    inv01 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix420 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx419), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_5)) ;
    xnor2 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix422 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx421), .A0 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx423), .A1 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx425)) ;
    xnor2 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix426 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx425), .A0 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothOperand_5), .A1 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_5)) ;
    inv01 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix430 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx429), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_6)) ;
    xnor2 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix432 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx431), .A0 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx433), .A1 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx435)) ;
    xnor2 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix436 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx435), .A0 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothOperand_6), .A1 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_6)) ;
    inv01 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix440 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx439), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_7)) ;
    xnor2 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix442 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx441), .A0 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx443), .A1 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx445)) ;
    xnor2 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix446 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx445), .A0 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothOperand_7), .A1 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_7)) ;
    inv01 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix450 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx449), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_8)) ;
    xnor2 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix452 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx451), .A0 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx453), .A1 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx455)) ;
    xnor2 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix456 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx455), .A0 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothOperand_8), .A1 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_8)) ;
    xor2 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix317 (.Y (
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx316), .A0 (
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx461), .A1 (
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx463)) ;
    xnor2 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix464 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx463), .A0 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothOperand_9), .A1 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_9)) ;
    xor2 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix337 (.Y (
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx336), .A0 (
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx467), .A1 (
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx471)) ;
    inv01 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix470 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx469), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_9)) ;
    xnor2 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix472 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx471), .A0 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothOperand_10), .A1 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_10)) ;
    xor2 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix357 (.Y (
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx356), .A0 (
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx475), .A1 (
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx479)) ;
    inv01 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix478 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx477), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_10)) ;
    xnor2 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix480 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx479), .A0 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothOperand_11), .A1 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_11)) ;
    xor2 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix377 (.Y (
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx376), .A0 (
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx483), .A1 (
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx487)) ;
    inv01 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix486 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx485), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_11)) ;
    xnor2 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix488 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx487), .A0 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothOperand_12), .A1 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_12)) ;
    xor2 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix397 (.Y (
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx396), .A0 (
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx491), .A1 (
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx495)) ;
    inv01 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix494 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx493), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_12)) ;
    xnor2 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix496 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx495), .A0 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothOperand_13), .A1 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_13)) ;
    xor2 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix417 (.Y (
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx416), .A0 (
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx499), .A1 (
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx503)) ;
    inv01 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix502 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx501), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_13)) ;
    xnor2 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix504 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx503), .A0 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothOperand_14), .A1 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_14)) ;
    xor2 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix437 (.Y (
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx436), .A0 (
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx507), .A1 (
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx511)) ;
    inv01 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix510 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx509), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_14)) ;
    xnor2 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix512 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx511), .A0 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothOperand_15), .A1 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_15)) ;
    xnor2 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix457 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx456), .A0 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx515), .A1 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx454)) ;
    inv01 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix518 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx517), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_15)) ;
    xor2 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix455 (.Y (
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx454), .A0 (
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothOperand_16), .A1 (
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_16)) ;
    mux21_ni CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix91 (.Y (
             CALCULATOR_L1SecondOperands_7__0), .A0 (
             CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_1), .A1 (
             CacheWindow_1__2__0), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix99 (.Y (
             CALCULATOR_L1SecondOperands_7__1), .A0 (
             CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_2), .A1 (
             CacheWindow_1__2__1), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix107 (.Y (
             CALCULATOR_L1SecondOperands_7__2), .A0 (
             CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_3), .A1 (
             CacheWindow_1__2__2), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix115 (.Y (
             CALCULATOR_L1SecondOperands_7__3), .A0 (
             CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_4), .A1 (
             CacheWindow_1__2__3), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix123 (.Y (
             CALCULATOR_L1SecondOperands_7__4), .A0 (
             CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_5), .A1 (
             CacheWindow_1__2__4), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix131 (.Y (
             CALCULATOR_L1SecondOperands_7__5), .A0 (
             CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_6), .A1 (
             CacheWindow_1__2__5), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix139 (.Y (
             CALCULATOR_L1SecondOperands_7__6), .A0 (
             CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_7), .A1 (
             CacheWindow_1__2__6), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix147 (.Y (
             CALCULATOR_L1SecondOperands_7__7), .A0 (
             CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_8), .A1 (
             CacheWindow_1__2__7), .S0 (Instr)) ;
    xor2 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix77 (.Y (CALCULATOR_L1Results_7__1), 
         .A0 (CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx529), .A1 (
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx531)) ;
    nand02 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix530 (.Y (
           CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx529), .A0 (
           CALCULATOR_L1SecondOperands_7__0), .A1 (
           CALCULATOR_L1FirstOperands_7__0)) ;
    xnor2 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix532 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx531), .A0 (
          CALCULATOR_L1SecondOperands_7__1), .A1 (
          CALCULATOR_L1FirstOperands_7__1)) ;
    xor2 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix75 (.Y (CALCULATOR_L1Results_7__2), 
         .A0 (CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx534), .A1 (
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx537)) ;
    aoi32 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix535 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx534), .A0 (
          CALCULATOR_L1SecondOperands_7__0), .A1 (
          CALCULATOR_L1FirstOperands_7__0), .A2 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx30), .B0 (
          CALCULATOR_L1FirstOperands_7__1), .B1 (
          CALCULATOR_L1SecondOperands_7__1)) ;
    xnor2 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix538 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx537), .A0 (
          CALCULATOR_L1SecondOperands_7__2), .A1 (
          CALCULATOR_L1FirstOperands_7__2)) ;
    xor2 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix73 (.Y (CALCULATOR_L1Results_7__3), 
         .A0 (CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx540), .A1 (
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx544)) ;
    aoi22 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix541 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx540), .A0 (
          CALCULATOR_L1FirstOperands_7__2), .A1 (
          CALCULATOR_L1SecondOperands_7__2), .B0 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx40), .B1 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx24)) ;
    xnor2 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix545 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx544), .A0 (
          CALCULATOR_L1SecondOperands_7__3), .A1 (
          CALCULATOR_L1FirstOperands_7__3)) ;
    xor2 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix71 (.Y (CALCULATOR_L1Results_7__4), 
         .A0 (CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx547), .A1 (
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx551)) ;
    aoi22 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix548 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx547), .A0 (
          CALCULATOR_L1FirstOperands_7__3), .A1 (
          CALCULATOR_L1SecondOperands_7__3), .B0 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx44), .B1 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx18)) ;
    xnor2 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix552 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx551), .A0 (
          CALCULATOR_L1SecondOperands_7__4), .A1 (
          CALCULATOR_L1FirstOperands_7__4)) ;
    xor2 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix69 (.Y (CALCULATOR_L1Results_7__5), 
         .A0 (CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx554), .A1 (
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx558)) ;
    aoi22 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix555 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx554), .A0 (
          CALCULATOR_L1FirstOperands_7__4), .A1 (
          CALCULATOR_L1SecondOperands_7__4), .B0 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx48), .B1 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx12)) ;
    xnor2 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix559 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx558), .A0 (
          CALCULATOR_L1SecondOperands_7__5), .A1 (
          CALCULATOR_L1FirstOperands_7__5)) ;
    xor2 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix67 (.Y (CALCULATOR_L1Results_7__6), 
         .A0 (CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx561), .A1 (
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx565)) ;
    aoi22 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix562 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx561), .A0 (
          CALCULATOR_L1FirstOperands_7__5), .A1 (
          CALCULATOR_L1SecondOperands_7__5), .B0 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx52), .B1 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx6)) ;
    xnor2 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix566 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx565), .A0 (
          CALCULATOR_L1SecondOperands_7__6), .A1 (
          CALCULATOR_L1FirstOperands_7__6)) ;
    xnor2 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix65 (.Y (CALCULATOR_L1Results_7__7)
          , .A0 (CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx568), .A1 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx62)) ;
    aoi22 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix569 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx568), .A0 (
          CALCULATOR_L1FirstOperands_7__6), .A1 (
          CALCULATOR_L1SecondOperands_7__6), .B0 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx56), .B1 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx0)) ;
    xor2 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix63 (.Y (
         CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx62), .A0 (
         CALCULATOR_L1SecondOperands_7__7), .A1 (CALCULATOR_L1FirstOperands_7__7
         )) ;
    inv01 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix155 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx154), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx383)) ;
    inv01 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix57 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx56), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx561)) ;
    inv01 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix53 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx52), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx554)) ;
    inv01 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix49 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx48), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx547)) ;
    inv01 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix45 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx44), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx540)) ;
    inv01 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix41 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx40), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx534)) ;
    inv01 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix31 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx30), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx531)) ;
    inv01 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix25 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx24), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx537)) ;
    inv01 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix19 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx18), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx544)) ;
    inv01 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix13 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx12), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx551)) ;
    inv01 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix7 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx6), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx558)) ;
    inv01 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix1 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx0), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx565)) ;
    fake_gnd CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix216 (.Y (
             CALCULATOR_L1_1_L2_2_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    aoi21 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix77 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_10), .A0 (
          CacheFilter_1__2__1), .A1 (CacheFilter_1__2__0), .B0 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx4)) ;
    nor02_2x CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix5 (.Y (
             CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx4), .A0 (
             CacheFilter_1__2__0), .A1 (CacheFilter_1__2__1)) ;
    aoi21 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix67 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_11), .A0 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx328), .A1 (
          CacheFilter_1__2__2), .B0 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx8)) ;
    nor03_2x CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix9 (.Y (
             CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx8), .A0 (
             CacheFilter_1__2__2), .A1 (CacheFilter_1__2__0), .A2 (
             CacheFilter_1__2__1)) ;
    xnor2 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix59 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_12), .A0 (
          CacheFilter_1__2__3), .A1 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx8)) ;
    xnor2 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix51 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_13), .A0 (
          CacheFilter_1__2__4), .A1 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx12)) ;
    nor04 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix13 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx12), .A0 (
          CacheFilter_1__2__3), .A1 (CacheFilter_1__2__2), .A2 (
          CacheFilter_1__2__0), .A3 (CacheFilter_1__2__1)) ;
    xnor2 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix43 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_14), .A0 (
          CacheFilter_1__2__5), .A1 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx16)) ;
    nor02ii CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix17 (.Y (
            CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx16), .A0 (
            CacheFilter_1__2__4), .A1 (
            CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx12)) ;
    xnor2 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix35 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_15), .A0 (
          CacheFilter_1__2__6), .A1 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx20)) ;
    nor02ii CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix21 (.Y (
            CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx20), .A0 (
            CacheFilter_1__2__5), .A1 (
            CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx16)) ;
    xnor2 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix27 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_16), .A0 (
          CacheFilter_1__2__7), .A1 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx24)) ;
    nor02ii CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix25 (.Y (
            CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx24), .A0 (
            CacheFilter_1__2__6), .A1 (
            CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx20)) ;
    inv01 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix329 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx328), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx4)) ;
    inv02 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix383 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx384), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_0)) ;
    dff CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_0 (.Q (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_0), .QB (
        \$dummy [384]), .D (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .CLK (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    nor02_2x CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix567 (.Y (
             CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566), .A0 (
             RST), .A1 (
             CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644)) ;
    dff CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_1 (.Q (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_1), .QB (
        \$dummy [385]), .D (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .CLK (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_2 (.Q (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_2), .QB (
        \$dummy [386]), .D (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .CLK (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_3 (.Q (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_3), .QB (
        \$dummy [387]), .D (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .CLK (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_4 (.Q (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_4), .QB (
        \$dummy [388]), .D (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .CLK (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_5 (.Q (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_5), .QB (
        \$dummy [389]), .D (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .CLK (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_6 (.Q (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_6), .QB (
        \$dummy [390]), .D (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .CLK (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_7 (.Q (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_7), .QB (
        \$dummy [391]), .D (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .CLK (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_8 (.Q (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_8), .QB (
        \$dummy [392]), .D (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .CLK (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_9 (.Q (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_9), .QB (
        \$dummy [393]), .D (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .CLK (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_10 (.Q (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_10), .QB (
        \$dummy [394]), .D (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .CLK (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_11 (.Q (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_11), .QB (
        \$dummy [395]), .D (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .CLK (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_12 (.Q (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_12), .QB (
        \$dummy [396]), .D (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .CLK (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_13 (.Q (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_13), .QB (
        \$dummy [397]), .D (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .CLK (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_14 (.Q (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_14), .QB (
        \$dummy [398]), .D (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .CLK (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_15 (.Q (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_15), .QB (
        \$dummy [399]), .D (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .CLK (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_16 (.Q (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_16), .QB (
        \$dummy [400]), .D (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .CLK (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    inv02 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix623 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix625 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix627 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix643 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644), .A (
          nx7659)) ;
    dff CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_0 (.Q (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_0), .QB (
        \$dummy [401]), .D (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .CLK (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    nor02_2x CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix567 (.Y (
             CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566), .A0 (
             RST), .A1 (
             CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644)) ;
    dff CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_1 (.Q (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_1), .QB (
        \$dummy [402]), .D (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .CLK (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_2 (.Q (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_2), .QB (
        \$dummy [403]), .D (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .CLK (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_3 (.Q (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_3), .QB (
        \$dummy [404]), .D (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .CLK (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_4 (.Q (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_4), .QB (
        \$dummy [405]), .D (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .CLK (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_5 (.Q (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_5), .QB (
        \$dummy [406]), .D (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .CLK (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_6 (.Q (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_6), .QB (
        \$dummy [407]), .D (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .CLK (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_7 (.Q (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_7), .QB (
        \$dummy [408]), .D (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .CLK (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_8 (.Q (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_8), .QB (
        \$dummy [409]), .D (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .CLK (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_9 (.Q (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_9), .QB (
        \$dummy [410]), .D (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .CLK (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_10 (.Q (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_10), .QB (
        \$dummy [411]), .D (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .CLK (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_11 (.Q (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_11), .QB (
        \$dummy [412]), .D (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .CLK (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_12 (.Q (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_12), .QB (
        \$dummy [413]), .D (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .CLK (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_13 (.Q (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_13), .QB (
        \$dummy [414]), .D (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .CLK (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_14 (.Q (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_14), .QB (
        \$dummy [415]), .D (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .CLK (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_15 (.Q (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_15), .QB (
        \$dummy [416]), .D (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .CLK (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_16 (.Q (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_16), .QB (
        \$dummy [417]), .D (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .CLK (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    inv02 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix623 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix625 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix627 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix643 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644), .A (
          nx7665)) ;
    dff CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_0 (.Q (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_0), .QB (\$dummy [418]), .D (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .CLK (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    nor02_2x CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix567 (.Y (
             CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566), .A0 (
             RST), .A1 (
             CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    dff CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_1 (.Q (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_1), .QB (\$dummy [419]), .D (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .CLK (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_2 (.Q (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_2), .QB (\$dummy [420]), .D (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .CLK (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_3 (.Q (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_3), .QB (\$dummy [421]), .D (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .CLK (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_4 (.Q (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_4), .QB (\$dummy [422]), .D (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .CLK (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_5 (.Q (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_5), .QB (\$dummy [423]), .D (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .CLK (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_6 (.Q (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_6), .QB (\$dummy [424]), .D (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .CLK (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_7 (.Q (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_7), .QB (\$dummy [425]), .D (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .CLK (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_8 (.Q (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_8), .QB (\$dummy [426]), .D (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .CLK (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_9 (.Q (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_9), .QB (\$dummy [427]), .D (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .CLK (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_10 (.Q (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_10), .QB (\$dummy [428]), .D (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .CLK (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_11 (.Q (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_11), .QB (\$dummy [429]), .D (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .CLK (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_12 (.Q (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_12), .QB (\$dummy [430]), .D (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .CLK (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_13 (.Q (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_13), .QB (\$dummy [431]), .D (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .CLK (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_14 (.Q (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_14), .QB (\$dummy [432]), .D (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .CLK (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_15 (.Q (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_15), .QB (\$dummy [433]), .D (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .CLK (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_16 (.Q (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_16), .QB (\$dummy [434]), .D (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .CLK (
        CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    inv02 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix623 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix625 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix627 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix643 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642)) ;
    xor2 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix83 (.Y (CALCULATOR_L1Results_8__0), 
         .A0 (CALCULATOR_L1SecondOperands_8__0), .A1 (
         CALCULATOR_L1FirstOperands_8__0)) ;
    xnor2 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix380 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx379), .A0 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx381), .A1 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx383)) ;
    nand02 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix382 (.Y (
           CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx381), .A0 (
           CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothOperand_0), .A1 (nx7685)) ;
    xnor2 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix384 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx383), .A0 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothOperand_1), .A1 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_1)) ;
    inv01 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix388 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx387), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_2)) ;
    xnor2 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix390 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx389), .A0 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx391), .A1 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx395)) ;
    aoi32 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix392 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx391), .A0 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothOperand_0), .A1 (nx7685), .A2 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx154), .B0 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_1), .B1 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothOperand_1)) ;
    xnor2 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix396 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx395), .A0 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothOperand_2), .A1 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_2)) ;
    inv01 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix400 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx399), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_3)) ;
    xnor2 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix402 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx401), .A0 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx403), .A1 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx405)) ;
    xnor2 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix406 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx405), .A0 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothOperand_3), .A1 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_3)) ;
    inv01 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix410 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx409), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_4)) ;
    xnor2 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix412 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx411), .A0 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx413), .A1 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx415)) ;
    xnor2 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix416 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx415), .A0 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothOperand_4), .A1 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_4)) ;
    inv01 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix420 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx419), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_5)) ;
    xnor2 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix422 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx421), .A0 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx423), .A1 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx425)) ;
    xnor2 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix426 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx425), .A0 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothOperand_5), .A1 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_5)) ;
    inv01 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix430 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx429), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_6)) ;
    xnor2 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix432 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx431), .A0 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx433), .A1 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx435)) ;
    xnor2 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix436 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx435), .A0 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothOperand_6), .A1 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_6)) ;
    inv01 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix440 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx439), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_7)) ;
    xnor2 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix442 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx441), .A0 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx443), .A1 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx445)) ;
    xnor2 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix446 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx445), .A0 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothOperand_7), .A1 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_7)) ;
    inv01 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix450 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx449), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_8)) ;
    xnor2 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix452 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx451), .A0 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx453), .A1 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx455)) ;
    xnor2 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix456 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx455), .A0 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothOperand_8), .A1 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_8)) ;
    xor2 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix317 (.Y (
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx316), .A0 (
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx461), .A1 (
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx463)) ;
    xnor2 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix464 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx463), .A0 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothOperand_9), .A1 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_9)) ;
    xor2 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix337 (.Y (
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx336), .A0 (
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx467), .A1 (
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx471)) ;
    inv01 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix470 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx469), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_9)) ;
    xnor2 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix472 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx471), .A0 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothOperand_10), .A1 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_10)) ;
    xor2 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix357 (.Y (
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx356), .A0 (
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx475), .A1 (
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx479)) ;
    inv01 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix478 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx477), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_10)) ;
    xnor2 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix480 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx479), .A0 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothOperand_11), .A1 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_11)) ;
    xor2 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix377 (.Y (
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx376), .A0 (
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx483), .A1 (
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx487)) ;
    inv01 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix486 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx485), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_11)) ;
    xnor2 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix488 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx487), .A0 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothOperand_12), .A1 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_12)) ;
    xor2 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix397 (.Y (
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx396), .A0 (
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx491), .A1 (
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx495)) ;
    inv01 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix494 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx493), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_12)) ;
    xnor2 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix496 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx495), .A0 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothOperand_13), .A1 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_13)) ;
    xor2 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix417 (.Y (
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx416), .A0 (
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx499), .A1 (
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx503)) ;
    inv01 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix502 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx501), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_13)) ;
    xnor2 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix504 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx503), .A0 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothOperand_14), .A1 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_14)) ;
    xor2 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix437 (.Y (
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx436), .A0 (
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx507), .A1 (
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx511)) ;
    inv01 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix510 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx509), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_14)) ;
    xnor2 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix512 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx511), .A0 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothOperand_15), .A1 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_15)) ;
    xnor2 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix457 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx456), .A0 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx515), .A1 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx454)) ;
    inv01 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix518 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx517), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_15)) ;
    xor2 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix455 (.Y (
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx454), .A0 (
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothOperand_16), .A1 (
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_16)) ;
    mux21_ni CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix91 (.Y (
             CALCULATOR_L1SecondOperands_8__0), .A0 (
             CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_1), .A1 (
             CacheWindow_1__3__0), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix99 (.Y (
             CALCULATOR_L1SecondOperands_8__1), .A0 (
             CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_2), .A1 (
             CacheWindow_1__3__1), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix107 (.Y (
             CALCULATOR_L1SecondOperands_8__2), .A0 (
             CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_3), .A1 (
             CacheWindow_1__3__2), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix115 (.Y (
             CALCULATOR_L1SecondOperands_8__3), .A0 (
             CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_4), .A1 (
             CacheWindow_1__3__3), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix123 (.Y (
             CALCULATOR_L1SecondOperands_8__4), .A0 (
             CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_5), .A1 (
             CacheWindow_1__3__4), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix131 (.Y (
             CALCULATOR_L1SecondOperands_8__5), .A0 (
             CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_6), .A1 (
             CacheWindow_1__3__5), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix139 (.Y (
             CALCULATOR_L1SecondOperands_8__6), .A0 (
             CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_7), .A1 (
             CacheWindow_1__3__6), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix147 (.Y (
             CALCULATOR_L1SecondOperands_8__7), .A0 (
             CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_8), .A1 (
             CacheWindow_1__3__7), .S0 (Instr)) ;
    xor2 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix77 (.Y (CALCULATOR_L1Results_8__1), 
         .A0 (CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx529), .A1 (
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx531)) ;
    nand02 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix530 (.Y (
           CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx529), .A0 (
           CALCULATOR_L1SecondOperands_8__0), .A1 (
           CALCULATOR_L1FirstOperands_8__0)) ;
    xnor2 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix532 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx531), .A0 (
          CALCULATOR_L1SecondOperands_8__1), .A1 (
          CALCULATOR_L1FirstOperands_8__1)) ;
    xor2 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix75 (.Y (CALCULATOR_L1Results_8__2), 
         .A0 (CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx534), .A1 (
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx537)) ;
    aoi32 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix535 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx534), .A0 (
          CALCULATOR_L1SecondOperands_8__0), .A1 (
          CALCULATOR_L1FirstOperands_8__0), .A2 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx30), .B0 (
          CALCULATOR_L1FirstOperands_8__1), .B1 (
          CALCULATOR_L1SecondOperands_8__1)) ;
    xnor2 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix538 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx537), .A0 (
          CALCULATOR_L1SecondOperands_8__2), .A1 (
          CALCULATOR_L1FirstOperands_8__2)) ;
    xor2 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix73 (.Y (CALCULATOR_L1Results_8__3), 
         .A0 (CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx540), .A1 (
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx544)) ;
    aoi22 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix541 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx540), .A0 (
          CALCULATOR_L1FirstOperands_8__2), .A1 (
          CALCULATOR_L1SecondOperands_8__2), .B0 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx40), .B1 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx24)) ;
    xnor2 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix545 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx544), .A0 (
          CALCULATOR_L1SecondOperands_8__3), .A1 (
          CALCULATOR_L1FirstOperands_8__3)) ;
    xor2 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix71 (.Y (CALCULATOR_L1Results_8__4), 
         .A0 (CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx547), .A1 (
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx551)) ;
    aoi22 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix548 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx547), .A0 (
          CALCULATOR_L1FirstOperands_8__3), .A1 (
          CALCULATOR_L1SecondOperands_8__3), .B0 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx44), .B1 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx18)) ;
    xnor2 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix552 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx551), .A0 (
          CALCULATOR_L1SecondOperands_8__4), .A1 (
          CALCULATOR_L1FirstOperands_8__4)) ;
    xor2 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix69 (.Y (CALCULATOR_L1Results_8__5), 
         .A0 (CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx554), .A1 (
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx558)) ;
    aoi22 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix555 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx554), .A0 (
          CALCULATOR_L1FirstOperands_8__4), .A1 (
          CALCULATOR_L1SecondOperands_8__4), .B0 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx48), .B1 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx12)) ;
    xnor2 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix559 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx558), .A0 (
          CALCULATOR_L1SecondOperands_8__5), .A1 (
          CALCULATOR_L1FirstOperands_8__5)) ;
    xor2 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix67 (.Y (CALCULATOR_L1Results_8__6), 
         .A0 (CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx561), .A1 (
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx565)) ;
    aoi22 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix562 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx561), .A0 (
          CALCULATOR_L1FirstOperands_8__5), .A1 (
          CALCULATOR_L1SecondOperands_8__5), .B0 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx52), .B1 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx6)) ;
    xnor2 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix566 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx565), .A0 (
          CALCULATOR_L1SecondOperands_8__6), .A1 (
          CALCULATOR_L1FirstOperands_8__6)) ;
    xnor2 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix65 (.Y (CALCULATOR_L1Results_8__7)
          , .A0 (CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx568), .A1 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx62)) ;
    aoi22 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix569 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx568), .A0 (
          CALCULATOR_L1FirstOperands_8__6), .A1 (
          CALCULATOR_L1SecondOperands_8__6), .B0 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx56), .B1 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx0)) ;
    xor2 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix63 (.Y (
         CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx62), .A0 (
         CALCULATOR_L1SecondOperands_8__7), .A1 (CALCULATOR_L1FirstOperands_8__7
         )) ;
    inv01 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix155 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx154), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx383)) ;
    inv01 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix57 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx56), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx561)) ;
    inv01 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix53 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx52), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx554)) ;
    inv01 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix49 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx48), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx547)) ;
    inv01 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix45 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx44), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx540)) ;
    inv01 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix41 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx40), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx534)) ;
    inv01 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix31 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx30), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx531)) ;
    inv01 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix25 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx24), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx537)) ;
    inv01 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix19 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx18), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx544)) ;
    inv01 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix13 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx12), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx551)) ;
    inv01 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix7 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx6), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx558)) ;
    inv01 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix1 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx0), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx565)) ;
    fake_gnd CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix216 (.Y (
             CALCULATOR_L1_1_L2_3_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    aoi21 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix77 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_10), .A0 (
          CacheFilter_1__3__1), .A1 (CacheFilter_1__3__0), .B0 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx4)) ;
    nor02_2x CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix5 (.Y (
             CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx4), .A0 (
             CacheFilter_1__3__0), .A1 (CacheFilter_1__3__1)) ;
    aoi21 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix67 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_11), .A0 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx328), .A1 (
          CacheFilter_1__3__2), .B0 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx8)) ;
    nor03_2x CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix9 (.Y (
             CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx8), .A0 (
             CacheFilter_1__3__2), .A1 (CacheFilter_1__3__0), .A2 (
             CacheFilter_1__3__1)) ;
    xnor2 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix59 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_12), .A0 (
          CacheFilter_1__3__3), .A1 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx8)) ;
    xnor2 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix51 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_13), .A0 (
          CacheFilter_1__3__4), .A1 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx12)) ;
    nor04 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix13 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx12), .A0 (
          CacheFilter_1__3__3), .A1 (CacheFilter_1__3__2), .A2 (
          CacheFilter_1__3__0), .A3 (CacheFilter_1__3__1)) ;
    xnor2 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix43 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_14), .A0 (
          CacheFilter_1__3__5), .A1 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx16)) ;
    nor02ii CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix17 (.Y (
            CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx16), .A0 (
            CacheFilter_1__3__4), .A1 (
            CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx12)) ;
    xnor2 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix35 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_15), .A0 (
          CacheFilter_1__3__6), .A1 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx20)) ;
    nor02ii CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix21 (.Y (
            CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx20), .A0 (
            CacheFilter_1__3__5), .A1 (
            CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx16)) ;
    xnor2 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix27 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_16), .A0 (
          CacheFilter_1__3__7), .A1 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx24)) ;
    nor02ii CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix25 (.Y (
            CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx24), .A0 (
            CacheFilter_1__3__6), .A1 (
            CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx20)) ;
    inv01 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix329 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx328), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx4)) ;
    inv02 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix383 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx384), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_0)) ;
    dff CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_0 (.Q (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_0), .QB (
        \$dummy [435]), .D (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .CLK (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    nor02_2x CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix567 (.Y (
             CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566), .A0 (
             RST), .A1 (
             CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644)) ;
    dff CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_1 (.Q (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_1), .QB (
        \$dummy [436]), .D (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .CLK (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_2 (.Q (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_2), .QB (
        \$dummy [437]), .D (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .CLK (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_3 (.Q (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_3), .QB (
        \$dummy [438]), .D (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .CLK (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_4 (.Q (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_4), .QB (
        \$dummy [439]), .D (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .CLK (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_5 (.Q (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_5), .QB (
        \$dummy [440]), .D (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .CLK (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_6 (.Q (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_6), .QB (
        \$dummy [441]), .D (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .CLK (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_7 (.Q (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_7), .QB (
        \$dummy [442]), .D (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .CLK (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_8 (.Q (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_8), .QB (
        \$dummy [443]), .D (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .CLK (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_9 (.Q (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_9), .QB (
        \$dummy [444]), .D (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .CLK (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_10 (.Q (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_10), .QB (
        \$dummy [445]), .D (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .CLK (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_11 (.Q (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_11), .QB (
        \$dummy [446]), .D (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .CLK (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_12 (.Q (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_12), .QB (
        \$dummy [447]), .D (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .CLK (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_13 (.Q (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_13), .QB (
        \$dummy [448]), .D (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .CLK (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_14 (.Q (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_14), .QB (
        \$dummy [449]), .D (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .CLK (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_15 (.Q (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_15), .QB (
        \$dummy [450]), .D (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .CLK (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_16 (.Q (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_16), .QB (
        \$dummy [451]), .D (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .CLK (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    inv02 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix623 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix625 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix627 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix643 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644), .A (
          nx7699)) ;
    dff CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_0 (.Q (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_0), .QB (
        \$dummy [452]), .D (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .CLK (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    nor02_2x CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix567 (.Y (
             CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566), .A0 (
             RST), .A1 (
             CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644)) ;
    dff CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_1 (.Q (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_1), .QB (
        \$dummy [453]), .D (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .CLK (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_2 (.Q (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_2), .QB (
        \$dummy [454]), .D (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .CLK (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_3 (.Q (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_3), .QB (
        \$dummy [455]), .D (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .CLK (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_4 (.Q (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_4), .QB (
        \$dummy [456]), .D (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .CLK (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_5 (.Q (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_5), .QB (
        \$dummy [457]), .D (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .CLK (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_6 (.Q (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_6), .QB (
        \$dummy [458]), .D (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .CLK (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_7 (.Q (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_7), .QB (
        \$dummy [459]), .D (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .CLK (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_8 (.Q (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_8), .QB (
        \$dummy [460]), .D (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .CLK (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_9 (.Q (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_9), .QB (
        \$dummy [461]), .D (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .CLK (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_10 (.Q (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_10), .QB (
        \$dummy [462]), .D (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .CLK (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_11 (.Q (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_11), .QB (
        \$dummy [463]), .D (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .CLK (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_12 (.Q (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_12), .QB (
        \$dummy [464]), .D (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .CLK (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_13 (.Q (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_13), .QB (
        \$dummy [465]), .D (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .CLK (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_14 (.Q (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_14), .QB (
        \$dummy [466]), .D (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .CLK (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_15 (.Q (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_15), .QB (
        \$dummy [467]), .D (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .CLK (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_16 (.Q (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_16), .QB (
        \$dummy [468]), .D (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .CLK (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    inv02 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix623 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix625 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix627 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix643 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644), .A (
          nx7705)) ;
    dff CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_0 (.Q (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_0), .QB (\$dummy [469]), .D (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .CLK (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    nor02_2x CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix567 (.Y (
             CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566), .A0 (
             RST), .A1 (
             CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    dff CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_1 (.Q (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_1), .QB (\$dummy [470]), .D (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .CLK (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_2 (.Q (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_2), .QB (\$dummy [471]), .D (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .CLK (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_3 (.Q (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_3), .QB (\$dummy [472]), .D (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .CLK (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_4 (.Q (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_4), .QB (\$dummy [473]), .D (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .CLK (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_5 (.Q (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_5), .QB (\$dummy [474]), .D (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .CLK (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_6 (.Q (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_6), .QB (\$dummy [475]), .D (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .CLK (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_7 (.Q (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_7), .QB (\$dummy [476]), .D (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .CLK (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_8 (.Q (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_8), .QB (\$dummy [477]), .D (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .CLK (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_9 (.Q (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_9), .QB (\$dummy [478]), .D (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .CLK (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_10 (.Q (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_10), .QB (\$dummy [479]), .D (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .CLK (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_11 (.Q (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_11), .QB (\$dummy [480]), .D (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .CLK (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_12 (.Q (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_12), .QB (\$dummy [481]), .D (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .CLK (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_13 (.Q (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_13), .QB (\$dummy [482]), .D (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .CLK (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_14 (.Q (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_14), .QB (\$dummy [483]), .D (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .CLK (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_15 (.Q (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_15), .QB (\$dummy [484]), .D (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .CLK (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_16 (.Q (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_16), .QB (\$dummy [485]), .D (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .CLK (
        CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    inv02 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix623 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix625 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix627 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix643 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642)) ;
    xor2 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix83 (.Y (CALCULATOR_L1Results_9__0), 
         .A0 (CALCULATOR_L1SecondOperands_9__0), .A1 (
         CALCULATOR_L1FirstOperands_9__0)) ;
    xnor2 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix380 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx379), .A0 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx381), .A1 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx383)) ;
    nand02 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix382 (.Y (
           CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx381), .A0 (
           CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothOperand_0), .A1 (nx7725)) ;
    xnor2 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix384 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx383), .A0 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothOperand_1), .A1 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_1)) ;
    inv01 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix388 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx387), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_2)) ;
    xnor2 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix390 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx389), .A0 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx391), .A1 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx395)) ;
    aoi32 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix392 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx391), .A0 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothOperand_0), .A1 (nx7725), .A2 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx154), .B0 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_1), .B1 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothOperand_1)) ;
    xnor2 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix396 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx395), .A0 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothOperand_2), .A1 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_2)) ;
    inv01 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix400 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx399), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_3)) ;
    xnor2 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix402 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx401), .A0 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx403), .A1 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx405)) ;
    xnor2 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix406 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx405), .A0 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothOperand_3), .A1 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_3)) ;
    inv01 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix410 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx409), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_4)) ;
    xnor2 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix412 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx411), .A0 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx413), .A1 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx415)) ;
    xnor2 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix416 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx415), .A0 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothOperand_4), .A1 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_4)) ;
    inv01 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix420 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx419), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_5)) ;
    xnor2 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix422 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx421), .A0 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx423), .A1 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx425)) ;
    xnor2 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix426 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx425), .A0 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothOperand_5), .A1 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_5)) ;
    inv01 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix430 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx429), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_6)) ;
    xnor2 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix432 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx431), .A0 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx433), .A1 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx435)) ;
    xnor2 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix436 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx435), .A0 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothOperand_6), .A1 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_6)) ;
    inv01 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix440 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx439), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_7)) ;
    xnor2 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix442 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx441), .A0 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx443), .A1 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx445)) ;
    xnor2 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix446 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx445), .A0 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothOperand_7), .A1 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_7)) ;
    inv01 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix450 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx449), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_8)) ;
    xnor2 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix452 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx451), .A0 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx453), .A1 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx455)) ;
    xnor2 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix456 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx455), .A0 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothOperand_8), .A1 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_8)) ;
    xor2 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix317 (.Y (
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx316), .A0 (
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx461), .A1 (
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx463)) ;
    xnor2 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix464 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx463), .A0 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothOperand_9), .A1 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_9)) ;
    xor2 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix337 (.Y (
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx336), .A0 (
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx467), .A1 (
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx471)) ;
    inv01 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix470 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx469), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_9)) ;
    xnor2 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix472 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx471), .A0 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothOperand_10), .A1 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_10)) ;
    xor2 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix357 (.Y (
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx356), .A0 (
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx475), .A1 (
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx479)) ;
    inv01 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix478 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx477), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_10)) ;
    xnor2 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix480 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx479), .A0 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothOperand_11), .A1 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_11)) ;
    xor2 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix377 (.Y (
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx376), .A0 (
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx483), .A1 (
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx487)) ;
    inv01 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix486 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx485), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_11)) ;
    xnor2 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix488 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx487), .A0 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothOperand_12), .A1 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_12)) ;
    xor2 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix397 (.Y (
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx396), .A0 (
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx491), .A1 (
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx495)) ;
    inv01 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix494 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx493), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_12)) ;
    xnor2 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix496 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx495), .A0 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothOperand_13), .A1 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_13)) ;
    xor2 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix417 (.Y (
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx416), .A0 (
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx499), .A1 (
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx503)) ;
    inv01 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix502 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx501), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_13)) ;
    xnor2 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix504 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx503), .A0 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothOperand_14), .A1 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_14)) ;
    xor2 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix437 (.Y (
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx436), .A0 (
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx507), .A1 (
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx511)) ;
    inv01 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix510 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx509), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_14)) ;
    xnor2 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix512 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx511), .A0 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothOperand_15), .A1 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_15)) ;
    xnor2 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix457 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx456), .A0 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx515), .A1 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx454)) ;
    inv01 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix518 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx517), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_15)) ;
    xor2 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix455 (.Y (
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx454), .A0 (
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothOperand_16), .A1 (
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_16)) ;
    mux21_ni CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix91 (.Y (
             CALCULATOR_L1SecondOperands_9__0), .A0 (
             CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_1), .A1 (
             CacheWindow_1__4__0), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix99 (.Y (
             CALCULATOR_L1SecondOperands_9__1), .A0 (
             CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_2), .A1 (
             CacheWindow_1__4__1), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix107 (.Y (
             CALCULATOR_L1SecondOperands_9__2), .A0 (
             CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_3), .A1 (
             CacheWindow_1__4__2), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix115 (.Y (
             CALCULATOR_L1SecondOperands_9__3), .A0 (
             CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_4), .A1 (
             CacheWindow_1__4__3), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix123 (.Y (
             CALCULATOR_L1SecondOperands_9__4), .A0 (
             CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_5), .A1 (
             CacheWindow_1__4__4), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix131 (.Y (
             CALCULATOR_L1SecondOperands_9__5), .A0 (
             CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_6), .A1 (
             CacheWindow_1__4__5), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix139 (.Y (
             CALCULATOR_L1SecondOperands_9__6), .A0 (
             CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_7), .A1 (
             CacheWindow_1__4__6), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix147 (.Y (
             CALCULATOR_L1SecondOperands_9__7), .A0 (
             CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_8), .A1 (
             CacheWindow_1__4__7), .S0 (Instr)) ;
    xor2 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix77 (.Y (CALCULATOR_L1Results_9__1), 
         .A0 (CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx529), .A1 (
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx531)) ;
    nand02 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix530 (.Y (
           CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx529), .A0 (
           CALCULATOR_L1SecondOperands_9__0), .A1 (
           CALCULATOR_L1FirstOperands_9__0)) ;
    xnor2 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix532 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx531), .A0 (
          CALCULATOR_L1SecondOperands_9__1), .A1 (
          CALCULATOR_L1FirstOperands_9__1)) ;
    xor2 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix75 (.Y (CALCULATOR_L1Results_9__2), 
         .A0 (CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx534), .A1 (
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx537)) ;
    aoi32 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix535 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx534), .A0 (
          CALCULATOR_L1SecondOperands_9__0), .A1 (
          CALCULATOR_L1FirstOperands_9__0), .A2 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx30), .B0 (
          CALCULATOR_L1FirstOperands_9__1), .B1 (
          CALCULATOR_L1SecondOperands_9__1)) ;
    xnor2 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix538 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx537), .A0 (
          CALCULATOR_L1SecondOperands_9__2), .A1 (
          CALCULATOR_L1FirstOperands_9__2)) ;
    xor2 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix73 (.Y (CALCULATOR_L1Results_9__3), 
         .A0 (CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx540), .A1 (
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx544)) ;
    aoi22 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix541 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx540), .A0 (
          CALCULATOR_L1FirstOperands_9__2), .A1 (
          CALCULATOR_L1SecondOperands_9__2), .B0 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx40), .B1 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx24)) ;
    xnor2 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix545 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx544), .A0 (
          CALCULATOR_L1SecondOperands_9__3), .A1 (
          CALCULATOR_L1FirstOperands_9__3)) ;
    xor2 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix71 (.Y (CALCULATOR_L1Results_9__4), 
         .A0 (CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx547), .A1 (
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx551)) ;
    aoi22 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix548 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx547), .A0 (
          CALCULATOR_L1FirstOperands_9__3), .A1 (
          CALCULATOR_L1SecondOperands_9__3), .B0 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx44), .B1 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx18)) ;
    xnor2 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix552 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx551), .A0 (
          CALCULATOR_L1SecondOperands_9__4), .A1 (
          CALCULATOR_L1FirstOperands_9__4)) ;
    xor2 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix69 (.Y (CALCULATOR_L1Results_9__5), 
         .A0 (CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx554), .A1 (
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx558)) ;
    aoi22 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix555 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx554), .A0 (
          CALCULATOR_L1FirstOperands_9__4), .A1 (
          CALCULATOR_L1SecondOperands_9__4), .B0 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx48), .B1 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx12)) ;
    xnor2 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix559 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx558), .A0 (
          CALCULATOR_L1SecondOperands_9__5), .A1 (
          CALCULATOR_L1FirstOperands_9__5)) ;
    xor2 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix67 (.Y (CALCULATOR_L1Results_9__6), 
         .A0 (CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx561), .A1 (
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx565)) ;
    aoi22 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix562 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx561), .A0 (
          CALCULATOR_L1FirstOperands_9__5), .A1 (
          CALCULATOR_L1SecondOperands_9__5), .B0 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx52), .B1 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx6)) ;
    xnor2 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix566 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx565), .A0 (
          CALCULATOR_L1SecondOperands_9__6), .A1 (
          CALCULATOR_L1FirstOperands_9__6)) ;
    xnor2 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix65 (.Y (CALCULATOR_L1Results_9__7)
          , .A0 (CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx568), .A1 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx62)) ;
    aoi22 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix569 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx568), .A0 (
          CALCULATOR_L1FirstOperands_9__6), .A1 (
          CALCULATOR_L1SecondOperands_9__6), .B0 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx56), .B1 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx0)) ;
    xor2 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix63 (.Y (
         CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx62), .A0 (
         CALCULATOR_L1SecondOperands_9__7), .A1 (CALCULATOR_L1FirstOperands_9__7
         )) ;
    inv01 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix155 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx154), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx383)) ;
    inv01 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix57 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx56), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx561)) ;
    inv01 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix53 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx52), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx554)) ;
    inv01 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix49 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx48), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx547)) ;
    inv01 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix45 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx44), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx540)) ;
    inv01 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix41 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx40), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx534)) ;
    inv01 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix31 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx30), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx531)) ;
    inv01 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix25 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx24), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx537)) ;
    inv01 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix19 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx18), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx544)) ;
    inv01 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix13 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx12), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx551)) ;
    inv01 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix7 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx6), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx558)) ;
    inv01 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix1 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx0), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx565)) ;
    fake_gnd CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix216 (.Y (
             CALCULATOR_L1_1_L2_4_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    aoi21 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix77 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_10), .A0 (
          CacheFilter_1__4__1), .A1 (CacheFilter_1__4__0), .B0 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx4)) ;
    nor02_2x CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix5 (.Y (
             CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx4), .A0 (
             CacheFilter_1__4__0), .A1 (CacheFilter_1__4__1)) ;
    aoi21 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix67 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_11), .A0 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx328), .A1 (
          CacheFilter_1__4__2), .B0 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx8)) ;
    nor03_2x CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix9 (.Y (
             CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx8), .A0 (
             CacheFilter_1__4__2), .A1 (CacheFilter_1__4__0), .A2 (
             CacheFilter_1__4__1)) ;
    xnor2 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix59 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_12), .A0 (
          CacheFilter_1__4__3), .A1 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx8)) ;
    xnor2 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix51 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_13), .A0 (
          CacheFilter_1__4__4), .A1 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx12)) ;
    nor04 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix13 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx12), .A0 (
          CacheFilter_1__4__3), .A1 (CacheFilter_1__4__2), .A2 (
          CacheFilter_1__4__0), .A3 (CacheFilter_1__4__1)) ;
    xnor2 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix43 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_14), .A0 (
          CacheFilter_1__4__5), .A1 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx16)) ;
    nor02ii CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix17 (.Y (
            CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx16), .A0 (
            CacheFilter_1__4__4), .A1 (
            CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx12)) ;
    xnor2 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix35 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_15), .A0 (
          CacheFilter_1__4__6), .A1 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx20)) ;
    nor02ii CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix21 (.Y (
            CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx20), .A0 (
            CacheFilter_1__4__5), .A1 (
            CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx16)) ;
    xnor2 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix27 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_16), .A0 (
          CacheFilter_1__4__7), .A1 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx24)) ;
    nor02ii CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix25 (.Y (
            CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx24), .A0 (
            CacheFilter_1__4__6), .A1 (
            CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx20)) ;
    inv01 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix329 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx328), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx4)) ;
    inv02 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix383 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx384), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_0)) ;
    dff CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_0 (.Q (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_0), .QB (
        \$dummy [486]), .D (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .CLK (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    nor02_2x CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix567 (.Y (
             CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566), .A0 (
             RST), .A1 (
             CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644)) ;
    dff CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_1 (.Q (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_1), .QB (
        \$dummy [487]), .D (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .CLK (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_2 (.Q (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_2), .QB (
        \$dummy [488]), .D (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .CLK (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_3 (.Q (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_3), .QB (
        \$dummy [489]), .D (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .CLK (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_4 (.Q (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_4), .QB (
        \$dummy [490]), .D (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .CLK (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_5 (.Q (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_5), .QB (
        \$dummy [491]), .D (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .CLK (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_6 (.Q (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_6), .QB (
        \$dummy [492]), .D (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .CLK (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_7 (.Q (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_7), .QB (
        \$dummy [493]), .D (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .CLK (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_8 (.Q (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_8), .QB (
        \$dummy [494]), .D (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .CLK (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_9 (.Q (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_9), .QB (
        \$dummy [495]), .D (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .CLK (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_10 (.Q (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_10), .QB (
        \$dummy [496]), .D (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .CLK (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_11 (.Q (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_11), .QB (
        \$dummy [497]), .D (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .CLK (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_12 (.Q (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_12), .QB (
        \$dummy [498]), .D (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .CLK (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_13 (.Q (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_13), .QB (
        \$dummy [499]), .D (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .CLK (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_14 (.Q (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_14), .QB (
        \$dummy [500]), .D (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .CLK (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_15 (.Q (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_15), .QB (
        \$dummy [501]), .D (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .CLK (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_16 (.Q (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_16), .QB (
        \$dummy [502]), .D (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .CLK (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    inv02 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix623 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix625 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix627 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix643 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644), .A (
          nx7739)) ;
    dff CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_0 (.Q (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_0), .QB (
        \$dummy [503]), .D (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .CLK (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    nor02_2x CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix567 (.Y (
             CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566), .A0 (
             RST), .A1 (
             CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644)) ;
    dff CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_1 (.Q (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_1), .QB (
        \$dummy [504]), .D (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .CLK (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_2 (.Q (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_2), .QB (
        \$dummy [505]), .D (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .CLK (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_3 (.Q (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_3), .QB (
        \$dummy [506]), .D (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .CLK (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_4 (.Q (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_4), .QB (
        \$dummy [507]), .D (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .CLK (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_5 (.Q (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_5), .QB (
        \$dummy [508]), .D (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .CLK (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_6 (.Q (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_6), .QB (
        \$dummy [509]), .D (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .CLK (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_7 (.Q (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_7), .QB (
        \$dummy [510]), .D (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .CLK (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_8 (.Q (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_8), .QB (
        \$dummy [511]), .D (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .CLK (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_9 (.Q (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_9), .QB (
        \$dummy [512]), .D (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .CLK (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_10 (.Q (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_10), .QB (
        \$dummy [513]), .D (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .CLK (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_11 (.Q (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_11), .QB (
        \$dummy [514]), .D (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .CLK (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_12 (.Q (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_12), .QB (
        \$dummy [515]), .D (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .CLK (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_13 (.Q (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_13), .QB (
        \$dummy [516]), .D (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .CLK (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_14 (.Q (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_14), .QB (
        \$dummy [517]), .D (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .CLK (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_15 (.Q (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_15), .QB (
        \$dummy [518]), .D (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .CLK (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_16 (.Q (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_16), .QB (
        \$dummy [519]), .D (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .CLK (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    inv02 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix623 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix625 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix627 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix643 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644), .A (
          nx7745)) ;
    dff CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_0 (.Q (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_0), .QB (\$dummy [520]), .D (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .CLK (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    nor02_2x CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix567 (.Y (
             CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566), .A0 (
             RST), .A1 (
             CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    dff CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_1 (.Q (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_1), .QB (\$dummy [521]), .D (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .CLK (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_2 (.Q (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_2), .QB (\$dummy [522]), .D (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .CLK (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_3 (.Q (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_3), .QB (\$dummy [523]), .D (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .CLK (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_4 (.Q (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_4), .QB (\$dummy [524]), .D (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .CLK (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_5 (.Q (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_5), .QB (\$dummy [525]), .D (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .CLK (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_6 (.Q (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_6), .QB (\$dummy [526]), .D (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .CLK (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_7 (.Q (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_7), .QB (\$dummy [527]), .D (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .CLK (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_8 (.Q (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_8), .QB (\$dummy [528]), .D (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .CLK (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_9 (.Q (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_9), .QB (\$dummy [529]), .D (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .CLK (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_10 (.Q (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_10), .QB (\$dummy [530]), .D (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .CLK (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_11 (.Q (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_11), .QB (\$dummy [531]), .D (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .CLK (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_12 (.Q (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_12), .QB (\$dummy [532]), .D (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .CLK (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_13 (.Q (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_13), .QB (\$dummy [533]), .D (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .CLK (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_14 (.Q (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_14), .QB (\$dummy [534]), .D (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .CLK (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_15 (.Q (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_15), .QB (\$dummy [535]), .D (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .CLK (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_16 (.Q (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_16), .QB (\$dummy [536]), .D (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .CLK (
        CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    inv02 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix623 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix625 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix627 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix643 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642)) ;
    xor2 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix83 (.Y (CALCULATOR_L1Results_10__0)
         , .A0 (CALCULATOR_L1SecondOperands_10__0), .A1 (
         CALCULATOR_L1FirstOperands_10__0)) ;
    xnor2 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix380 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx379), .A0 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx381), .A1 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx383)) ;
    nand02 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix382 (.Y (
           CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx381), .A0 (
           CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothOperand_0), .A1 (nx7765)) ;
    xnor2 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix384 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx383), .A0 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothOperand_1), .A1 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_1)) ;
    inv01 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix388 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx387), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_2)) ;
    xnor2 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix390 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx389), .A0 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx391), .A1 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx395)) ;
    aoi32 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix392 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx391), .A0 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothOperand_0), .A1 (nx7765), .A2 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx154), .B0 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_1), .B1 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothOperand_1)) ;
    xnor2 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix396 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx395), .A0 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothOperand_2), .A1 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_2)) ;
    inv01 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix400 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx399), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_3)) ;
    xnor2 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix402 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx401), .A0 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx403), .A1 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx405)) ;
    xnor2 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix406 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx405), .A0 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothOperand_3), .A1 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_3)) ;
    inv01 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix410 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx409), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_4)) ;
    xnor2 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix412 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx411), .A0 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx413), .A1 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx415)) ;
    xnor2 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix416 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx415), .A0 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothOperand_4), .A1 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_4)) ;
    inv01 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix420 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx419), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_5)) ;
    xnor2 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix422 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx421), .A0 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx423), .A1 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx425)) ;
    xnor2 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix426 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx425), .A0 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothOperand_5), .A1 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_5)) ;
    inv01 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix430 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx429), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_6)) ;
    xnor2 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix432 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx431), .A0 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx433), .A1 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx435)) ;
    xnor2 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix436 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx435), .A0 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothOperand_6), .A1 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_6)) ;
    inv01 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix440 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx439), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_7)) ;
    xnor2 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix442 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx441), .A0 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx443), .A1 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx445)) ;
    xnor2 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix446 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx445), .A0 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothOperand_7), .A1 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_7)) ;
    inv01 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix450 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx449), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_8)) ;
    xnor2 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix452 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx451), .A0 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx453), .A1 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx455)) ;
    xnor2 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix456 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx455), .A0 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothOperand_8), .A1 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_8)) ;
    xor2 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix317 (.Y (
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx316), .A0 (
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx461), .A1 (
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx463)) ;
    xnor2 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix464 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx463), .A0 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothOperand_9), .A1 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_9)) ;
    xor2 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix337 (.Y (
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx336), .A0 (
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx467), .A1 (
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx471)) ;
    inv01 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix470 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx469), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_9)) ;
    xnor2 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix472 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx471), .A0 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothOperand_10), .A1 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_10)) ;
    xor2 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix357 (.Y (
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx356), .A0 (
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx475), .A1 (
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx479)) ;
    inv01 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix478 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx477), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_10)) ;
    xnor2 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix480 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx479), .A0 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothOperand_11), .A1 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_11)) ;
    xor2 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix377 (.Y (
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx376), .A0 (
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx483), .A1 (
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx487)) ;
    inv01 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix486 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx485), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_11)) ;
    xnor2 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix488 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx487), .A0 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothOperand_12), .A1 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_12)) ;
    xor2 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix397 (.Y (
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx396), .A0 (
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx491), .A1 (
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx495)) ;
    inv01 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix494 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx493), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_12)) ;
    xnor2 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix496 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx495), .A0 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothOperand_13), .A1 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_13)) ;
    xor2 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix417 (.Y (
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx416), .A0 (
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx499), .A1 (
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx503)) ;
    inv01 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix502 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx501), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_13)) ;
    xnor2 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix504 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx503), .A0 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothOperand_14), .A1 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_14)) ;
    xor2 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix437 (.Y (
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx436), .A0 (
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx507), .A1 (
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx511)) ;
    inv01 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix510 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx509), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_14)) ;
    xnor2 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix512 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx511), .A0 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothOperand_15), .A1 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_15)) ;
    xnor2 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix457 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx456), .A0 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx515), .A1 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx454)) ;
    inv01 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix518 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx517), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_15)) ;
    xor2 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix455 (.Y (
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx454), .A0 (
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothOperand_16), .A1 (
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_16)) ;
    mux21_ni CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix91 (.Y (
             CALCULATOR_L1SecondOperands_10__0), .A0 (
             CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_1), .A1 (
             CacheWindow_2__0__0), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix99 (.Y (
             CALCULATOR_L1SecondOperands_10__1), .A0 (
             CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_2), .A1 (
             CacheWindow_2__0__1), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix107 (.Y (
             CALCULATOR_L1SecondOperands_10__2), .A0 (
             CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_3), .A1 (
             CacheWindow_2__0__2), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix115 (.Y (
             CALCULATOR_L1SecondOperands_10__3), .A0 (
             CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_4), .A1 (
             CacheWindow_2__0__3), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix123 (.Y (
             CALCULATOR_L1SecondOperands_10__4), .A0 (
             CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_5), .A1 (
             CacheWindow_2__0__4), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix131 (.Y (
             CALCULATOR_L1SecondOperands_10__5), .A0 (
             CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_6), .A1 (
             CacheWindow_2__0__5), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix139 (.Y (
             CALCULATOR_L1SecondOperands_10__6), .A0 (
             CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_7), .A1 (
             CacheWindow_2__0__6), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix147 (.Y (
             CALCULATOR_L1SecondOperands_10__7), .A0 (
             CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_8), .A1 (
             CacheWindow_2__0__7), .S0 (Instr)) ;
    xor2 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix77 (.Y (CALCULATOR_L1Results_10__1)
         , .A0 (CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx529), .A1 (
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx531)) ;
    nand02 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix530 (.Y (
           CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx529), .A0 (
           CALCULATOR_L1SecondOperands_10__0), .A1 (
           CALCULATOR_L1FirstOperands_10__0)) ;
    xnor2 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix532 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx531), .A0 (
          CALCULATOR_L1SecondOperands_10__1), .A1 (
          CALCULATOR_L1FirstOperands_10__1)) ;
    xor2 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix75 (.Y (CALCULATOR_L1Results_10__2)
         , .A0 (CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx534), .A1 (
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx537)) ;
    aoi32 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix535 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx534), .A0 (
          CALCULATOR_L1SecondOperands_10__0), .A1 (
          CALCULATOR_L1FirstOperands_10__0), .A2 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx30), .B0 (
          CALCULATOR_L1FirstOperands_10__1), .B1 (
          CALCULATOR_L1SecondOperands_10__1)) ;
    xnor2 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix538 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx537), .A0 (
          CALCULATOR_L1SecondOperands_10__2), .A1 (
          CALCULATOR_L1FirstOperands_10__2)) ;
    xor2 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix73 (.Y (CALCULATOR_L1Results_10__3)
         , .A0 (CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx540), .A1 (
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx544)) ;
    aoi22 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix541 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx540), .A0 (
          CALCULATOR_L1FirstOperands_10__2), .A1 (
          CALCULATOR_L1SecondOperands_10__2), .B0 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx40), .B1 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx24)) ;
    xnor2 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix545 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx544), .A0 (
          CALCULATOR_L1SecondOperands_10__3), .A1 (
          CALCULATOR_L1FirstOperands_10__3)) ;
    xor2 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix71 (.Y (CALCULATOR_L1Results_10__4)
         , .A0 (CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx547), .A1 (
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx551)) ;
    aoi22 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix548 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx547), .A0 (
          CALCULATOR_L1FirstOperands_10__3), .A1 (
          CALCULATOR_L1SecondOperands_10__3), .B0 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx44), .B1 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx18)) ;
    xnor2 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix552 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx551), .A0 (
          CALCULATOR_L1SecondOperands_10__4), .A1 (
          CALCULATOR_L1FirstOperands_10__4)) ;
    xor2 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix69 (.Y (CALCULATOR_L1Results_10__5)
         , .A0 (CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx554), .A1 (
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx558)) ;
    aoi22 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix555 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx554), .A0 (
          CALCULATOR_L1FirstOperands_10__4), .A1 (
          CALCULATOR_L1SecondOperands_10__4), .B0 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx48), .B1 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx12)) ;
    xnor2 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix559 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx558), .A0 (
          CALCULATOR_L1SecondOperands_10__5), .A1 (
          CALCULATOR_L1FirstOperands_10__5)) ;
    xor2 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix67 (.Y (CALCULATOR_L1Results_10__6)
         , .A0 (CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx561), .A1 (
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx565)) ;
    aoi22 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix562 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx561), .A0 (
          CALCULATOR_L1FirstOperands_10__5), .A1 (
          CALCULATOR_L1SecondOperands_10__5), .B0 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx52), .B1 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx6)) ;
    xnor2 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix566 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx565), .A0 (
          CALCULATOR_L1SecondOperands_10__6), .A1 (
          CALCULATOR_L1FirstOperands_10__6)) ;
    xnor2 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix65 (.Y (CALCULATOR_L1Results_10__7)
          , .A0 (CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx568), .A1 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx62)) ;
    aoi22 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix569 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx568), .A0 (
          CALCULATOR_L1FirstOperands_10__6), .A1 (
          CALCULATOR_L1SecondOperands_10__6), .B0 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx56), .B1 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx0)) ;
    xor2 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix63 (.Y (
         CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx62), .A0 (
         CALCULATOR_L1SecondOperands_10__7), .A1 (
         CALCULATOR_L1FirstOperands_10__7)) ;
    inv01 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix155 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx154), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx383)) ;
    inv01 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix57 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx56), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx561)) ;
    inv01 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix53 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx52), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx554)) ;
    inv01 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix49 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx48), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx547)) ;
    inv01 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix45 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx44), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx540)) ;
    inv01 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix41 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx40), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx534)) ;
    inv01 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix31 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx30), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx531)) ;
    inv01 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix25 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx24), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx537)) ;
    inv01 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix19 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx18), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx544)) ;
    inv01 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix13 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx12), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx551)) ;
    inv01 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix7 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx6), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx558)) ;
    inv01 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix1 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx0), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx565)) ;
    fake_gnd CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix216 (.Y (
             CALCULATOR_L1_2_L2_0_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    aoi21 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix77 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_10), .A0 (
          CacheFilter_2__0__1), .A1 (CacheFilter_2__0__0), .B0 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx4)) ;
    nor02_2x CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix5 (.Y (
             CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx4), .A0 (
             CacheFilter_2__0__0), .A1 (CacheFilter_2__0__1)) ;
    aoi21 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix67 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_11), .A0 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx328), .A1 (
          CacheFilter_2__0__2), .B0 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx8)) ;
    nor03_2x CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix9 (.Y (
             CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx8), .A0 (
             CacheFilter_2__0__2), .A1 (CacheFilter_2__0__0), .A2 (
             CacheFilter_2__0__1)) ;
    xnor2 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix59 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_12), .A0 (
          CacheFilter_2__0__3), .A1 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx8)) ;
    xnor2 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix51 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_13), .A0 (
          CacheFilter_2__0__4), .A1 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx12)) ;
    nor04 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix13 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx12), .A0 (
          CacheFilter_2__0__3), .A1 (CacheFilter_2__0__2), .A2 (
          CacheFilter_2__0__0), .A3 (CacheFilter_2__0__1)) ;
    xnor2 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix43 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_14), .A0 (
          CacheFilter_2__0__5), .A1 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx16)) ;
    nor02ii CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix17 (.Y (
            CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx16), .A0 (
            CacheFilter_2__0__4), .A1 (
            CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx12)) ;
    xnor2 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix35 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_15), .A0 (
          CacheFilter_2__0__6), .A1 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx20)) ;
    nor02ii CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix21 (.Y (
            CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx20), .A0 (
            CacheFilter_2__0__5), .A1 (
            CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx16)) ;
    xnor2 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix27 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_16), .A0 (
          CacheFilter_2__0__7), .A1 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx24)) ;
    nor02ii CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix25 (.Y (
            CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx24), .A0 (
            CacheFilter_2__0__6), .A1 (
            CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx20)) ;
    inv01 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix329 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx328), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx4)) ;
    inv02 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix383 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx384), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_0)) ;
    dff CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_0 (.Q (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_0), .QB (
        \$dummy [537]), .D (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .CLK (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    nor02_2x CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix567 (.Y (
             CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566), .A0 (
             RST), .A1 (
             CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644)) ;
    dff CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_1 (.Q (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_1), .QB (
        \$dummy [538]), .D (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .CLK (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_2 (.Q (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_2), .QB (
        \$dummy [539]), .D (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .CLK (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_3 (.Q (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_3), .QB (
        \$dummy [540]), .D (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .CLK (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_4 (.Q (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_4), .QB (
        \$dummy [541]), .D (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .CLK (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_5 (.Q (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_5), .QB (
        \$dummy [542]), .D (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .CLK (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_6 (.Q (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_6), .QB (
        \$dummy [543]), .D (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .CLK (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_7 (.Q (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_7), .QB (
        \$dummy [544]), .D (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .CLK (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_8 (.Q (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_8), .QB (
        \$dummy [545]), .D (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .CLK (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_9 (.Q (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_9), .QB (
        \$dummy [546]), .D (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .CLK (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_10 (.Q (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_10), .QB (
        \$dummy [547]), .D (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .CLK (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_11 (.Q (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_11), .QB (
        \$dummy [548]), .D (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .CLK (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_12 (.Q (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_12), .QB (
        \$dummy [549]), .D (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .CLK (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_13 (.Q (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_13), .QB (
        \$dummy [550]), .D (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .CLK (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_14 (.Q (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_14), .QB (
        \$dummy [551]), .D (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .CLK (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_15 (.Q (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_15), .QB (
        \$dummy [552]), .D (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .CLK (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_16 (.Q (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_16), .QB (
        \$dummy [553]), .D (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .CLK (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    inv02 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix623 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix625 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix627 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix643 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644), .A (
          nx7779)) ;
    dff CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_0 (.Q (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_0), .QB (
        \$dummy [554]), .D (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .CLK (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    nor02_2x CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix567 (.Y (
             CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566), .A0 (
             RST), .A1 (
             CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644)) ;
    dff CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_1 (.Q (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_1), .QB (
        \$dummy [555]), .D (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .CLK (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_2 (.Q (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_2), .QB (
        \$dummy [556]), .D (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .CLK (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_3 (.Q (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_3), .QB (
        \$dummy [557]), .D (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .CLK (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_4 (.Q (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_4), .QB (
        \$dummy [558]), .D (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .CLK (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_5 (.Q (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_5), .QB (
        \$dummy [559]), .D (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .CLK (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_6 (.Q (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_6), .QB (
        \$dummy [560]), .D (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .CLK (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_7 (.Q (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_7), .QB (
        \$dummy [561]), .D (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .CLK (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_8 (.Q (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_8), .QB (
        \$dummy [562]), .D (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .CLK (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_9 (.Q (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_9), .QB (
        \$dummy [563]), .D (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .CLK (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_10 (.Q (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_10), .QB (
        \$dummy [564]), .D (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .CLK (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_11 (.Q (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_11), .QB (
        \$dummy [565]), .D (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .CLK (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_12 (.Q (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_12), .QB (
        \$dummy [566]), .D (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .CLK (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_13 (.Q (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_13), .QB (
        \$dummy [567]), .D (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .CLK (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_14 (.Q (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_14), .QB (
        \$dummy [568]), .D (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .CLK (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_15 (.Q (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_15), .QB (
        \$dummy [569]), .D (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .CLK (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_16 (.Q (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_16), .QB (
        \$dummy [570]), .D (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .CLK (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    inv02 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix623 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix625 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix627 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix643 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644), .A (
          nx7785)) ;
    dff CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_0 (.Q (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_0), .QB (\$dummy [571]), .D (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .CLK (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    nor02_2x CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix567 (.Y (
             CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566), .A0 (
             RST), .A1 (
             CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    dff CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_1 (.Q (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_1), .QB (\$dummy [572]), .D (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .CLK (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_2 (.Q (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_2), .QB (\$dummy [573]), .D (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .CLK (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_3 (.Q (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_3), .QB (\$dummy [574]), .D (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .CLK (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_4 (.Q (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_4), .QB (\$dummy [575]), .D (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .CLK (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_5 (.Q (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_5), .QB (\$dummy [576]), .D (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .CLK (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_6 (.Q (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_6), .QB (\$dummy [577]), .D (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .CLK (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_7 (.Q (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_7), .QB (\$dummy [578]), .D (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .CLK (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_8 (.Q (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_8), .QB (\$dummy [579]), .D (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .CLK (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_9 (.Q (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_9), .QB (\$dummy [580]), .D (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .CLK (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_10 (.Q (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_10), .QB (\$dummy [581]), .D (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .CLK (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_11 (.Q (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_11), .QB (\$dummy [582]), .D (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .CLK (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_12 (.Q (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_12), .QB (\$dummy [583]), .D (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .CLK (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_13 (.Q (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_13), .QB (\$dummy [584]), .D (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .CLK (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_14 (.Q (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_14), .QB (\$dummy [585]), .D (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .CLK (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_15 (.Q (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_15), .QB (\$dummy [586]), .D (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .CLK (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_16 (.Q (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_16), .QB (\$dummy [587]), .D (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .CLK (
        CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    inv02 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix623 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix625 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix627 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix643 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642)) ;
    xor2 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix83 (.Y (CALCULATOR_L1Results_11__0)
         , .A0 (CALCULATOR_L1SecondOperands_11__0), .A1 (
         CALCULATOR_L1FirstOperands_11__0)) ;
    xnor2 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix380 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx379), .A0 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx381), .A1 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx383)) ;
    nand02 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix382 (.Y (
           CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx381), .A0 (
           CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothOperand_0), .A1 (nx7805)) ;
    xnor2 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix384 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx383), .A0 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothOperand_1), .A1 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_1)) ;
    inv01 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix388 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx387), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_2)) ;
    xnor2 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix390 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx389), .A0 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx391), .A1 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx395)) ;
    aoi32 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix392 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx391), .A0 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothOperand_0), .A1 (nx7805), .A2 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx154), .B0 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_1), .B1 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothOperand_1)) ;
    xnor2 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix396 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx395), .A0 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothOperand_2), .A1 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_2)) ;
    inv01 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix400 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx399), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_3)) ;
    xnor2 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix402 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx401), .A0 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx403), .A1 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx405)) ;
    xnor2 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix406 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx405), .A0 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothOperand_3), .A1 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_3)) ;
    inv01 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix410 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx409), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_4)) ;
    xnor2 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix412 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx411), .A0 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx413), .A1 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx415)) ;
    xnor2 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix416 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx415), .A0 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothOperand_4), .A1 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_4)) ;
    inv01 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix420 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx419), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_5)) ;
    xnor2 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix422 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx421), .A0 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx423), .A1 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx425)) ;
    xnor2 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix426 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx425), .A0 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothOperand_5), .A1 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_5)) ;
    inv01 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix430 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx429), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_6)) ;
    xnor2 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix432 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx431), .A0 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx433), .A1 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx435)) ;
    xnor2 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix436 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx435), .A0 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothOperand_6), .A1 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_6)) ;
    inv01 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix440 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx439), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_7)) ;
    xnor2 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix442 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx441), .A0 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx443), .A1 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx445)) ;
    xnor2 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix446 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx445), .A0 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothOperand_7), .A1 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_7)) ;
    inv01 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix450 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx449), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_8)) ;
    xnor2 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix452 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx451), .A0 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx453), .A1 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx455)) ;
    xnor2 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix456 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx455), .A0 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothOperand_8), .A1 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_8)) ;
    xor2 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix317 (.Y (
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx316), .A0 (
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx461), .A1 (
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx463)) ;
    xnor2 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix464 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx463), .A0 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothOperand_9), .A1 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_9)) ;
    xor2 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix337 (.Y (
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx336), .A0 (
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx467), .A1 (
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx471)) ;
    inv01 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix470 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx469), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_9)) ;
    xnor2 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix472 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx471), .A0 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothOperand_10), .A1 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_10)) ;
    xor2 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix357 (.Y (
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx356), .A0 (
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx475), .A1 (
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx479)) ;
    inv01 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix478 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx477), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_10)) ;
    xnor2 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix480 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx479), .A0 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothOperand_11), .A1 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_11)) ;
    xor2 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix377 (.Y (
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx376), .A0 (
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx483), .A1 (
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx487)) ;
    inv01 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix486 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx485), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_11)) ;
    xnor2 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix488 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx487), .A0 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothOperand_12), .A1 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_12)) ;
    xor2 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix397 (.Y (
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx396), .A0 (
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx491), .A1 (
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx495)) ;
    inv01 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix494 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx493), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_12)) ;
    xnor2 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix496 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx495), .A0 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothOperand_13), .A1 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_13)) ;
    xor2 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix417 (.Y (
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx416), .A0 (
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx499), .A1 (
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx503)) ;
    inv01 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix502 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx501), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_13)) ;
    xnor2 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix504 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx503), .A0 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothOperand_14), .A1 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_14)) ;
    xor2 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix437 (.Y (
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx436), .A0 (
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx507), .A1 (
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx511)) ;
    inv01 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix510 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx509), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_14)) ;
    xnor2 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix512 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx511), .A0 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothOperand_15), .A1 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_15)) ;
    xnor2 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix457 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx456), .A0 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx515), .A1 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx454)) ;
    inv01 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix518 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx517), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_15)) ;
    xor2 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix455 (.Y (
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx454), .A0 (
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothOperand_16), .A1 (
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_16)) ;
    mux21_ni CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix91 (.Y (
             CALCULATOR_L1SecondOperands_11__0), .A0 (
             CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_1), .A1 (
             CacheWindow_2__1__0), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix99 (.Y (
             CALCULATOR_L1SecondOperands_11__1), .A0 (
             CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_2), .A1 (
             CacheWindow_2__1__1), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix107 (.Y (
             CALCULATOR_L1SecondOperands_11__2), .A0 (
             CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_3), .A1 (
             CacheWindow_2__1__2), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix115 (.Y (
             CALCULATOR_L1SecondOperands_11__3), .A0 (
             CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_4), .A1 (
             CacheWindow_2__1__3), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix123 (.Y (
             CALCULATOR_L1SecondOperands_11__4), .A0 (
             CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_5), .A1 (
             CacheWindow_2__1__4), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix131 (.Y (
             CALCULATOR_L1SecondOperands_11__5), .A0 (
             CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_6), .A1 (
             CacheWindow_2__1__5), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix139 (.Y (
             CALCULATOR_L1SecondOperands_11__6), .A0 (
             CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_7), .A1 (
             CacheWindow_2__1__6), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix147 (.Y (
             CALCULATOR_L1SecondOperands_11__7), .A0 (
             CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_8), .A1 (
             CacheWindow_2__1__7), .S0 (Instr)) ;
    xor2 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix77 (.Y (CALCULATOR_L1Results_11__1)
         , .A0 (CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx529), .A1 (
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx531)) ;
    nand02 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix530 (.Y (
           CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx529), .A0 (
           CALCULATOR_L1SecondOperands_11__0), .A1 (
           CALCULATOR_L1FirstOperands_11__0)) ;
    xnor2 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix532 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx531), .A0 (
          CALCULATOR_L1SecondOperands_11__1), .A1 (
          CALCULATOR_L1FirstOperands_11__1)) ;
    xor2 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix75 (.Y (CALCULATOR_L1Results_11__2)
         , .A0 (CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx534), .A1 (
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx537)) ;
    aoi32 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix535 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx534), .A0 (
          CALCULATOR_L1SecondOperands_11__0), .A1 (
          CALCULATOR_L1FirstOperands_11__0), .A2 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx30), .B0 (
          CALCULATOR_L1FirstOperands_11__1), .B1 (
          CALCULATOR_L1SecondOperands_11__1)) ;
    xnor2 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix538 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx537), .A0 (
          CALCULATOR_L1SecondOperands_11__2), .A1 (
          CALCULATOR_L1FirstOperands_11__2)) ;
    xor2 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix73 (.Y (CALCULATOR_L1Results_11__3)
         , .A0 (CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx540), .A1 (
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx544)) ;
    aoi22 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix541 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx540), .A0 (
          CALCULATOR_L1FirstOperands_11__2), .A1 (
          CALCULATOR_L1SecondOperands_11__2), .B0 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx40), .B1 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx24)) ;
    xnor2 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix545 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx544), .A0 (
          CALCULATOR_L1SecondOperands_11__3), .A1 (
          CALCULATOR_L1FirstOperands_11__3)) ;
    xor2 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix71 (.Y (CALCULATOR_L1Results_11__4)
         , .A0 (CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx547), .A1 (
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx551)) ;
    aoi22 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix548 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx547), .A0 (
          CALCULATOR_L1FirstOperands_11__3), .A1 (
          CALCULATOR_L1SecondOperands_11__3), .B0 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx44), .B1 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx18)) ;
    xnor2 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix552 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx551), .A0 (
          CALCULATOR_L1SecondOperands_11__4), .A1 (
          CALCULATOR_L1FirstOperands_11__4)) ;
    xor2 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix69 (.Y (CALCULATOR_L1Results_11__5)
         , .A0 (CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx554), .A1 (
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx558)) ;
    aoi22 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix555 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx554), .A0 (
          CALCULATOR_L1FirstOperands_11__4), .A1 (
          CALCULATOR_L1SecondOperands_11__4), .B0 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx48), .B1 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx12)) ;
    xnor2 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix559 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx558), .A0 (
          CALCULATOR_L1SecondOperands_11__5), .A1 (
          CALCULATOR_L1FirstOperands_11__5)) ;
    xor2 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix67 (.Y (CALCULATOR_L1Results_11__6)
         , .A0 (CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx561), .A1 (
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx565)) ;
    aoi22 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix562 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx561), .A0 (
          CALCULATOR_L1FirstOperands_11__5), .A1 (
          CALCULATOR_L1SecondOperands_11__5), .B0 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx52), .B1 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx6)) ;
    xnor2 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix566 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx565), .A0 (
          CALCULATOR_L1SecondOperands_11__6), .A1 (
          CALCULATOR_L1FirstOperands_11__6)) ;
    xnor2 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix65 (.Y (CALCULATOR_L1Results_11__7)
          , .A0 (CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx568), .A1 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx62)) ;
    aoi22 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix569 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx568), .A0 (
          CALCULATOR_L1FirstOperands_11__6), .A1 (
          CALCULATOR_L1SecondOperands_11__6), .B0 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx56), .B1 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx0)) ;
    xor2 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix63 (.Y (
         CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx62), .A0 (
         CALCULATOR_L1SecondOperands_11__7), .A1 (
         CALCULATOR_L1FirstOperands_11__7)) ;
    inv01 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix155 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx154), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx383)) ;
    inv01 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix57 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx56), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx561)) ;
    inv01 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix53 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx52), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx554)) ;
    inv01 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix49 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx48), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx547)) ;
    inv01 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix45 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx44), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx540)) ;
    inv01 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix41 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx40), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx534)) ;
    inv01 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix31 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx30), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx531)) ;
    inv01 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix25 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx24), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx537)) ;
    inv01 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix19 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx18), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx544)) ;
    inv01 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix13 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx12), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx551)) ;
    inv01 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix7 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx6), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx558)) ;
    inv01 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix1 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx0), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx565)) ;
    fake_gnd CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix216 (.Y (
             CALCULATOR_L1_2_L2_1_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    aoi21 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix77 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_10), .A0 (
          CacheFilter_2__1__1), .A1 (CacheFilter_2__1__0), .B0 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx4)) ;
    nor02_2x CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix5 (.Y (
             CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx4), .A0 (
             CacheFilter_2__1__0), .A1 (CacheFilter_2__1__1)) ;
    aoi21 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix67 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_11), .A0 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx328), .A1 (
          CacheFilter_2__1__2), .B0 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx8)) ;
    nor03_2x CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix9 (.Y (
             CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx8), .A0 (
             CacheFilter_2__1__2), .A1 (CacheFilter_2__1__0), .A2 (
             CacheFilter_2__1__1)) ;
    xnor2 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix59 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_12), .A0 (
          CacheFilter_2__1__3), .A1 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx8)) ;
    xnor2 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix51 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_13), .A0 (
          CacheFilter_2__1__4), .A1 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx12)) ;
    nor04 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix13 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx12), .A0 (
          CacheFilter_2__1__3), .A1 (CacheFilter_2__1__2), .A2 (
          CacheFilter_2__1__0), .A3 (CacheFilter_2__1__1)) ;
    xnor2 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix43 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_14), .A0 (
          CacheFilter_2__1__5), .A1 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx16)) ;
    nor02ii CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix17 (.Y (
            CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx16), .A0 (
            CacheFilter_2__1__4), .A1 (
            CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx12)) ;
    xnor2 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix35 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_15), .A0 (
          CacheFilter_2__1__6), .A1 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx20)) ;
    nor02ii CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix21 (.Y (
            CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx20), .A0 (
            CacheFilter_2__1__5), .A1 (
            CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx16)) ;
    xnor2 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix27 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_16), .A0 (
          CacheFilter_2__1__7), .A1 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx24)) ;
    nor02ii CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix25 (.Y (
            CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx24), .A0 (
            CacheFilter_2__1__6), .A1 (
            CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx20)) ;
    inv01 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix329 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx328), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx4)) ;
    inv02 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix383 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx384), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_0)) ;
    dff CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_0 (.Q (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_0), .QB (
        \$dummy [588]), .D (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .CLK (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    nor02_2x CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix567 (.Y (
             CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566), .A0 (
             RST), .A1 (
             CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644)) ;
    dff CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_1 (.Q (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_1), .QB (
        \$dummy [589]), .D (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .CLK (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_2 (.Q (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_2), .QB (
        \$dummy [590]), .D (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .CLK (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_3 (.Q (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_3), .QB (
        \$dummy [591]), .D (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .CLK (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_4 (.Q (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_4), .QB (
        \$dummy [592]), .D (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .CLK (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_5 (.Q (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_5), .QB (
        \$dummy [593]), .D (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .CLK (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_6 (.Q (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_6), .QB (
        \$dummy [594]), .D (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .CLK (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_7 (.Q (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_7), .QB (
        \$dummy [595]), .D (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .CLK (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_8 (.Q (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_8), .QB (
        \$dummy [596]), .D (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .CLK (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_9 (.Q (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_9), .QB (
        \$dummy [597]), .D (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .CLK (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_10 (.Q (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_10), .QB (
        \$dummy [598]), .D (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .CLK (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_11 (.Q (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_11), .QB (
        \$dummy [599]), .D (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .CLK (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_12 (.Q (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_12), .QB (
        \$dummy [600]), .D (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .CLK (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_13 (.Q (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_13), .QB (
        \$dummy [601]), .D (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .CLK (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_14 (.Q (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_14), .QB (
        \$dummy [602]), .D (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .CLK (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_15 (.Q (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_15), .QB (
        \$dummy [603]), .D (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .CLK (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_16 (.Q (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_16), .QB (
        \$dummy [604]), .D (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .CLK (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    inv02 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix623 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix625 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix627 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix643 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644), .A (
          nx7819)) ;
    dff CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_0 (.Q (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_0), .QB (
        \$dummy [605]), .D (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .CLK (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    nor02_2x CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix567 (.Y (
             CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566), .A0 (
             RST), .A1 (
             CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644)) ;
    dff CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_1 (.Q (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_1), .QB (
        \$dummy [606]), .D (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .CLK (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_2 (.Q (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_2), .QB (
        \$dummy [607]), .D (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .CLK (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_3 (.Q (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_3), .QB (
        \$dummy [608]), .D (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .CLK (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_4 (.Q (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_4), .QB (
        \$dummy [609]), .D (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .CLK (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_5 (.Q (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_5), .QB (
        \$dummy [610]), .D (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .CLK (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_6 (.Q (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_6), .QB (
        \$dummy [611]), .D (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .CLK (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_7 (.Q (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_7), .QB (
        \$dummy [612]), .D (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .CLK (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_8 (.Q (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_8), .QB (
        \$dummy [613]), .D (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .CLK (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_9 (.Q (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_9), .QB (
        \$dummy [614]), .D (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .CLK (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_10 (.Q (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_10), .QB (
        \$dummy [615]), .D (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .CLK (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_11 (.Q (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_11), .QB (
        \$dummy [616]), .D (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .CLK (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_12 (.Q (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_12), .QB (
        \$dummy [617]), .D (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .CLK (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_13 (.Q (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_13), .QB (
        \$dummy [618]), .D (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .CLK (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_14 (.Q (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_14), .QB (
        \$dummy [619]), .D (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .CLK (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_15 (.Q (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_15), .QB (
        \$dummy [620]), .D (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .CLK (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_16 (.Q (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_16), .QB (
        \$dummy [621]), .D (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .CLK (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    inv02 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix623 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix625 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix627 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix643 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644), .A (
          nx7825)) ;
    dff CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_0 (.Q (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_0), .QB (\$dummy [622]), .D (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .CLK (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    nor02_2x CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix567 (.Y (
             CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566), .A0 (
             RST), .A1 (
             CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    dff CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_1 (.Q (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_1), .QB (\$dummy [623]), .D (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .CLK (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_2 (.Q (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_2), .QB (\$dummy [624]), .D (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .CLK (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_3 (.Q (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_3), .QB (\$dummy [625]), .D (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .CLK (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_4 (.Q (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_4), .QB (\$dummy [626]), .D (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .CLK (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_5 (.Q (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_5), .QB (\$dummy [627]), .D (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .CLK (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_6 (.Q (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_6), .QB (\$dummy [628]), .D (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .CLK (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_7 (.Q (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_7), .QB (\$dummy [629]), .D (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .CLK (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_8 (.Q (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_8), .QB (\$dummy [630]), .D (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .CLK (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_9 (.Q (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_9), .QB (\$dummy [631]), .D (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .CLK (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_10 (.Q (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_10), .QB (\$dummy [632]), .D (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .CLK (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_11 (.Q (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_11), .QB (\$dummy [633]), .D (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .CLK (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_12 (.Q (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_12), .QB (\$dummy [634]), .D (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .CLK (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_13 (.Q (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_13), .QB (\$dummy [635]), .D (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .CLK (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_14 (.Q (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_14), .QB (\$dummy [636]), .D (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .CLK (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_15 (.Q (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_15), .QB (\$dummy [637]), .D (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .CLK (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_16 (.Q (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_16), .QB (\$dummy [638]), .D (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .CLK (
        CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    inv02 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix623 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix625 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix627 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix643 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642)) ;
    xnor2 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix380 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx379), .A0 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx381), .A1 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx383)) ;
    nand02 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix382 (.Y (
           CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx381), .A0 (
           CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothOperand_0), .A1 (nx7845)) ;
    xnor2 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix384 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx383), .A0 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothOperand_1), .A1 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_1)) ;
    inv01 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix388 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx387), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_2)) ;
    xnor2 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix390 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx389), .A0 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx391), .A1 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx395)) ;
    aoi32 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix392 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx391), .A0 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothOperand_0), .A1 (nx7845), .A2 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx154), .B0 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_1), .B1 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothOperand_1)) ;
    xnor2 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix396 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx395), .A0 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothOperand_2), .A1 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_2)) ;
    inv01 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix400 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx399), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_3)) ;
    xnor2 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix402 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx401), .A0 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx403), .A1 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx405)) ;
    xnor2 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix406 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx405), .A0 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothOperand_3), .A1 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_3)) ;
    inv01 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix410 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx409), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_4)) ;
    xnor2 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix412 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx411), .A0 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx413), .A1 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx415)) ;
    xnor2 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix416 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx415), .A0 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothOperand_4), .A1 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_4)) ;
    inv01 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix420 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx419), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_5)) ;
    xnor2 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix422 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx421), .A0 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx423), .A1 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx425)) ;
    xnor2 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix426 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx425), .A0 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothOperand_5), .A1 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_5)) ;
    inv01 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix430 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx429), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_6)) ;
    xnor2 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix432 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx431), .A0 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx433), .A1 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx435)) ;
    xnor2 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix436 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx435), .A0 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothOperand_6), .A1 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_6)) ;
    inv01 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix440 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx439), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_7)) ;
    xnor2 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix442 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx441), .A0 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx443), .A1 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx445)) ;
    xnor2 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix446 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx445), .A0 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothOperand_7), .A1 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_7)) ;
    inv01 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix450 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx449), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_8)) ;
    xnor2 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix452 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx451), .A0 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx453), .A1 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx455)) ;
    xnor2 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix456 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx455), .A0 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothOperand_8), .A1 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_8)) ;
    xor2 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix317 (.Y (
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx316), .A0 (
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx461), .A1 (
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx463)) ;
    xnor2 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix464 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx463), .A0 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothOperand_9), .A1 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_9)) ;
    xor2 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix337 (.Y (
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx336), .A0 (
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx467), .A1 (
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx471)) ;
    inv01 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix470 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx469), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_9)) ;
    xnor2 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix472 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx471), .A0 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothOperand_10), .A1 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_10)) ;
    xor2 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix357 (.Y (
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx356), .A0 (
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx475), .A1 (
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx479)) ;
    inv01 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix478 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx477), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_10)) ;
    xnor2 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix480 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx479), .A0 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothOperand_11), .A1 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_11)) ;
    xor2 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix377 (.Y (
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx376), .A0 (
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx483), .A1 (
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx487)) ;
    inv01 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix486 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx485), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_11)) ;
    xnor2 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix488 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx487), .A0 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothOperand_12), .A1 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_12)) ;
    xor2 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix397 (.Y (
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx396), .A0 (
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx491), .A1 (
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx495)) ;
    inv01 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix494 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx493), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_12)) ;
    xnor2 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix496 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx495), .A0 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothOperand_13), .A1 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_13)) ;
    xor2 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix417 (.Y (
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx416), .A0 (
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx499), .A1 (
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx503)) ;
    inv01 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix502 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx501), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_13)) ;
    xnor2 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix504 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx503), .A0 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothOperand_14), .A1 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_14)) ;
    xor2 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix437 (.Y (
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx436), .A0 (
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx507), .A1 (
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx511)) ;
    inv01 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix510 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx509), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_14)) ;
    xnor2 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix512 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx511), .A0 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothOperand_15), .A1 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_15)) ;
    xnor2 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix457 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx456), .A0 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx515), .A1 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx454)) ;
    inv01 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix518 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx517), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_15)) ;
    xor2 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix455 (.Y (
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx454), .A0 (
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothOperand_16), .A1 (
         CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_16)) ;
    mux21_ni CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix91 (.Y (
             CALCULATOR_L1FirstOperands_11__0), .A0 (
             CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_1), .A1 (
             CacheWindow_2__2__0), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix99 (.Y (
             CALCULATOR_L1FirstOperands_11__1), .A0 (
             CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_2), .A1 (
             CacheWindow_2__2__1), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix107 (.Y (
             CALCULATOR_L1FirstOperands_11__2), .A0 (
             CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_3), .A1 (
             CacheWindow_2__2__2), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix115 (.Y (
             CALCULATOR_L1FirstOperands_11__3), .A0 (
             CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_4), .A1 (
             CacheWindow_2__2__3), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix123 (.Y (
             CALCULATOR_L1FirstOperands_11__4), .A0 (
             CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_5), .A1 (
             CacheWindow_2__2__4), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix131 (.Y (
             CALCULATOR_L1FirstOperands_11__5), .A0 (
             CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_6), .A1 (
             CacheWindow_2__2__5), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix139 (.Y (
             CALCULATOR_L1FirstOperands_11__6), .A0 (
             CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_7), .A1 (
             CacheWindow_2__2__6), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix147 (.Y (
             CALCULATOR_L1FirstOperands_11__7), .A0 (
             CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_8), .A1 (
             CacheWindow_2__2__7), .S0 (Instr)) ;
    inv01 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix155 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx154), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx383)) ;
    fake_gnd CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix216 (.Y (
             CALCULATOR_L1_2_L2_2_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    aoi21 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix77 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_10), .A0 (
          CacheFilter_2__2__1), .A1 (CacheFilter_2__2__0), .B0 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx4)) ;
    nor02_2x CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix5 (.Y (
             CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx4), .A0 (
             CacheFilter_2__2__0), .A1 (CacheFilter_2__2__1)) ;
    aoi21 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix67 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_11), .A0 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx328), .A1 (
          CacheFilter_2__2__2), .B0 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx8)) ;
    nor03_2x CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix9 (.Y (
             CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx8), .A0 (
             CacheFilter_2__2__2), .A1 (CacheFilter_2__2__0), .A2 (
             CacheFilter_2__2__1)) ;
    xnor2 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix59 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_12), .A0 (
          CacheFilter_2__2__3), .A1 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx8)) ;
    xnor2 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix51 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_13), .A0 (
          CacheFilter_2__2__4), .A1 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx12)) ;
    nor04 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix13 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx12), .A0 (
          CacheFilter_2__2__3), .A1 (CacheFilter_2__2__2), .A2 (
          CacheFilter_2__2__0), .A3 (CacheFilter_2__2__1)) ;
    xnor2 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix43 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_14), .A0 (
          CacheFilter_2__2__5), .A1 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx16)) ;
    nor02ii CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix17 (.Y (
            CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx16), .A0 (
            CacheFilter_2__2__4), .A1 (
            CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx12)) ;
    xnor2 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix35 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_15), .A0 (
          CacheFilter_2__2__6), .A1 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx20)) ;
    nor02ii CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix21 (.Y (
            CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx20), .A0 (
            CacheFilter_2__2__5), .A1 (
            CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx16)) ;
    xnor2 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix27 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_16), .A0 (
          CacheFilter_2__2__7), .A1 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx24)) ;
    nor02ii CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix25 (.Y (
            CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx24), .A0 (
            CacheFilter_2__2__6), .A1 (
            CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx20)) ;
    inv01 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix329 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx328), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx4)) ;
    inv02 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix383 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx384), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_0)) ;
    dff CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_0 (.Q (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_0), .QB (
        \$dummy [639]), .D (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .CLK (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    nor02_2x CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix567 (.Y (
             CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566), .A0 (
             RST), .A1 (
             CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644)) ;
    dff CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_1 (.Q (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_1), .QB (
        \$dummy [640]), .D (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .CLK (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_2 (.Q (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_2), .QB (
        \$dummy [641]), .D (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .CLK (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_3 (.Q (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_3), .QB (
        \$dummy [642]), .D (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .CLK (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_4 (.Q (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_4), .QB (
        \$dummy [643]), .D (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .CLK (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_5 (.Q (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_5), .QB (
        \$dummy [644]), .D (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .CLK (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_6 (.Q (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_6), .QB (
        \$dummy [645]), .D (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .CLK (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_7 (.Q (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_7), .QB (
        \$dummy [646]), .D (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .CLK (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_8 (.Q (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_8), .QB (
        \$dummy [647]), .D (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .CLK (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_9 (.Q (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_9), .QB (
        \$dummy [648]), .D (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .CLK (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_10 (.Q (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_10), .QB (
        \$dummy [649]), .D (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .CLK (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_11 (.Q (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_11), .QB (
        \$dummy [650]), .D (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .CLK (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_12 (.Q (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_12), .QB (
        \$dummy [651]), .D (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .CLK (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_13 (.Q (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_13), .QB (
        \$dummy [652]), .D (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .CLK (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_14 (.Q (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_14), .QB (
        \$dummy [653]), .D (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .CLK (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_15 (.Q (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_15), .QB (
        \$dummy [654]), .D (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .CLK (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_16 (.Q (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_16), .QB (
        \$dummy [655]), .D (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .CLK (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    inv02 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix623 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix625 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix627 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix643 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644), .A (
          nx7859)) ;
    dff CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_0 (.Q (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_0), .QB (
        \$dummy [656]), .D (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .CLK (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    nor02_2x CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix567 (.Y (
             CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566), .A0 (
             RST), .A1 (
             CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644)) ;
    dff CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_1 (.Q (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_1), .QB (
        \$dummy [657]), .D (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .CLK (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_2 (.Q (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_2), .QB (
        \$dummy [658]), .D (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .CLK (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_3 (.Q (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_3), .QB (
        \$dummy [659]), .D (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .CLK (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_4 (.Q (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_4), .QB (
        \$dummy [660]), .D (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .CLK (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_5 (.Q (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_5), .QB (
        \$dummy [661]), .D (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .CLK (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_6 (.Q (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_6), .QB (
        \$dummy [662]), .D (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .CLK (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_7 (.Q (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_7), .QB (
        \$dummy [663]), .D (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .CLK (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_8 (.Q (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_8), .QB (
        \$dummy [664]), .D (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .CLK (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_9 (.Q (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_9), .QB (
        \$dummy [665]), .D (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .CLK (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_10 (.Q (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_10), .QB (
        \$dummy [666]), .D (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .CLK (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_11 (.Q (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_11), .QB (
        \$dummy [667]), .D (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .CLK (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_12 (.Q (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_12), .QB (
        \$dummy [668]), .D (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .CLK (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_13 (.Q (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_13), .QB (
        \$dummy [669]), .D (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .CLK (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_14 (.Q (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_14), .QB (
        \$dummy [670]), .D (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .CLK (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_15 (.Q (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_15), .QB (
        \$dummy [671]), .D (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .CLK (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_16 (.Q (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_16), .QB (
        \$dummy [672]), .D (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .CLK (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    inv02 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix623 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix625 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix627 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix643 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644), .A (
          nx7865)) ;
    dff CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_0 (.Q (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_0), .QB (\$dummy [673]), .D (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .CLK (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    nor02_2x CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix567 (.Y (
             CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566), .A0 (
             RST), .A1 (
             CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    dff CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_1 (.Q (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_1), .QB (\$dummy [674]), .D (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .CLK (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_2 (.Q (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_2), .QB (\$dummy [675]), .D (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .CLK (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_3 (.Q (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_3), .QB (\$dummy [676]), .D (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .CLK (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_4 (.Q (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_4), .QB (\$dummy [677]), .D (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .CLK (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_5 (.Q (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_5), .QB (\$dummy [678]), .D (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .CLK (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_6 (.Q (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_6), .QB (\$dummy [679]), .D (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .CLK (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_7 (.Q (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_7), .QB (\$dummy [680]), .D (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .CLK (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_8 (.Q (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_8), .QB (\$dummy [681]), .D (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .CLK (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_9 (.Q (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_9), .QB (\$dummy [682]), .D (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .CLK (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_10 (.Q (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_10), .QB (\$dummy [683]), .D (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .CLK (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_11 (.Q (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_11), .QB (\$dummy [684]), .D (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .CLK (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_12 (.Q (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_12), .QB (\$dummy [685]), .D (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .CLK (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_13 (.Q (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_13), .QB (\$dummy [686]), .D (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .CLK (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_14 (.Q (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_14), .QB (\$dummy [687]), .D (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .CLK (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_15 (.Q (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_15), .QB (\$dummy [688]), .D (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .CLK (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_16 (.Q (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_16), .QB (\$dummy [689]), .D (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .CLK (
        CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    inv02 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix623 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix625 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix627 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix643 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642)) ;
    xor2 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix83 (.Y (CALCULATOR_L2Results_0__0), 
         .A0 (CALCULATOR_L1Results_1__0), .A1 (CALCULATOR_L1Results_0__0)) ;
    xnor2 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix380 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx379), .A0 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx381), .A1 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx383)) ;
    nand02 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix382 (.Y (
           CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx381), .A0 (
           CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothOperand_0), .A1 (nx7885)) ;
    xnor2 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix384 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx383), .A0 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothOperand_1), .A1 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_1)) ;
    inv01 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix388 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx387), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_2)) ;
    xnor2 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix390 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx389), .A0 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx391), .A1 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx395)) ;
    aoi32 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix392 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx391), .A0 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothOperand_0), .A1 (nx7885), .A2 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx154), .B0 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_1), .B1 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothOperand_1)) ;
    xnor2 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix396 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx395), .A0 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothOperand_2), .A1 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_2)) ;
    inv01 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix400 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx399), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_3)) ;
    xnor2 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix402 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx401), .A0 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx403), .A1 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx405)) ;
    xnor2 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix406 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx405), .A0 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothOperand_3), .A1 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_3)) ;
    inv01 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix410 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx409), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_4)) ;
    xnor2 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix412 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx411), .A0 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx413), .A1 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx415)) ;
    xnor2 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix416 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx415), .A0 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothOperand_4), .A1 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_4)) ;
    inv01 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix420 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx419), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_5)) ;
    xnor2 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix422 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx421), .A0 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx423), .A1 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx425)) ;
    xnor2 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix426 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx425), .A0 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothOperand_5), .A1 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_5)) ;
    inv01 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix430 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx429), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_6)) ;
    xnor2 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix432 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx431), .A0 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx433), .A1 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx435)) ;
    xnor2 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix436 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx435), .A0 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothOperand_6), .A1 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_6)) ;
    inv01 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix440 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx439), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_7)) ;
    xnor2 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix442 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx441), .A0 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx443), .A1 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx445)) ;
    xnor2 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix446 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx445), .A0 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothOperand_7), .A1 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_7)) ;
    inv01 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix450 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx449), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_8)) ;
    xnor2 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix452 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx451), .A0 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx453), .A1 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx455)) ;
    xnor2 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix456 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx455), .A0 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothOperand_8), .A1 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_8)) ;
    xor2 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix317 (.Y (
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx316), .A0 (
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx461), .A1 (
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx463)) ;
    xnor2 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix464 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx463), .A0 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothOperand_9), .A1 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_9)) ;
    xor2 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix337 (.Y (
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx336), .A0 (
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx467), .A1 (
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx471)) ;
    inv01 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix470 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx469), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_9)) ;
    xnor2 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix472 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx471), .A0 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothOperand_10), .A1 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_10)) ;
    xor2 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix357 (.Y (
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx356), .A0 (
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx475), .A1 (
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx479)) ;
    inv01 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix478 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx477), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_10)) ;
    xnor2 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix480 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx479), .A0 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothOperand_11), .A1 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_11)) ;
    xor2 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix377 (.Y (
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx376), .A0 (
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx483), .A1 (
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx487)) ;
    inv01 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix486 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx485), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_11)) ;
    xnor2 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix488 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx487), .A0 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothOperand_12), .A1 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_12)) ;
    xor2 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix397 (.Y (
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx396), .A0 (
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx491), .A1 (
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx495)) ;
    inv01 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix494 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx493), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_12)) ;
    xnor2 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix496 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx495), .A0 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothOperand_13), .A1 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_13)) ;
    xor2 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix417 (.Y (
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx416), .A0 (
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx499), .A1 (
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx503)) ;
    inv01 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix502 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx501), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_13)) ;
    xnor2 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix504 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx503), .A0 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothOperand_14), .A1 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_14)) ;
    xor2 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix437 (.Y (
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx436), .A0 (
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx507), .A1 (
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx511)) ;
    inv01 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix510 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx509), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_14)) ;
    xnor2 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix512 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx511), .A0 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothOperand_15), .A1 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_15)) ;
    xnor2 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix457 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx456), .A0 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx515), .A1 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx454)) ;
    inv01 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix518 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx517), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_15)) ;
    xor2 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix455 (.Y (
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx454), .A0 (
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothOperand_16), .A1 (
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_16)) ;
    mux21_ni CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix91 (.Y (
             CALCULATOR_L1FirstOperands_0__0), .A0 (
             CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_1), .A1 (
             CacheWindow_2__3__0), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix99 (.Y (
             CALCULATOR_L1FirstOperands_0__1), .A0 (
             CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_2), .A1 (
             CacheWindow_2__3__1), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix107 (.Y (
             CALCULATOR_L1FirstOperands_0__2), .A0 (
             CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_3), .A1 (
             CacheWindow_2__3__2), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix115 (.Y (
             CALCULATOR_L1FirstOperands_0__3), .A0 (
             CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_4), .A1 (
             CacheWindow_2__3__3), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix123 (.Y (
             CALCULATOR_L1FirstOperands_0__4), .A0 (
             CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_5), .A1 (
             CacheWindow_2__3__4), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix131 (.Y (
             CALCULATOR_L1FirstOperands_0__5), .A0 (
             CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_6), .A1 (
             CacheWindow_2__3__5), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix139 (.Y (
             CALCULATOR_L1FirstOperands_0__6), .A0 (
             CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_7), .A1 (
             CacheWindow_2__3__6), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix147 (.Y (
             CALCULATOR_L1FirstOperands_0__7), .A0 (
             CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_8), .A1 (
             CacheWindow_2__3__7), .S0 (Instr)) ;
    xor2 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix77 (.Y (CALCULATOR_L2Results_0__1), 
         .A0 (CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx529), .A1 (
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx531)) ;
    nand02 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix530 (.Y (
           CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx529), .A0 (
           CALCULATOR_L1Results_1__0), .A1 (CALCULATOR_L1Results_0__0)) ;
    xnor2 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix532 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx531), .A0 (
          CALCULATOR_L1Results_1__1), .A1 (CALCULATOR_L1Results_0__1)) ;
    xor2 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix75 (.Y (CALCULATOR_L2Results_0__2), 
         .A0 (CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx534), .A1 (
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx537)) ;
    aoi32 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix535 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx534), .A0 (
          CALCULATOR_L1Results_1__0), .A1 (CALCULATOR_L1Results_0__0), .A2 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx30), .B0 (CALCULATOR_L1Results_0__1
          ), .B1 (CALCULATOR_L1Results_1__1)) ;
    xnor2 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix538 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx537), .A0 (
          CALCULATOR_L1Results_1__2), .A1 (CALCULATOR_L1Results_0__2)) ;
    xor2 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix73 (.Y (CALCULATOR_L2Results_0__3), 
         .A0 (CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx540), .A1 (
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx544)) ;
    aoi22 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix541 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx540), .A0 (
          CALCULATOR_L1Results_0__2), .A1 (CALCULATOR_L1Results_1__2), .B0 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx40), .B1 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx24)) ;
    xnor2 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix545 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx544), .A0 (
          CALCULATOR_L1Results_1__3), .A1 (CALCULATOR_L1Results_0__3)) ;
    xor2 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix71 (.Y (CALCULATOR_L2Results_0__4), 
         .A0 (CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx547), .A1 (
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx551)) ;
    aoi22 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix548 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx547), .A0 (
          CALCULATOR_L1Results_0__3), .A1 (CALCULATOR_L1Results_1__3), .B0 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx44), .B1 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx18)) ;
    xnor2 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix552 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx551), .A0 (
          CALCULATOR_L1Results_1__4), .A1 (CALCULATOR_L1Results_0__4)) ;
    xor2 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix69 (.Y (CALCULATOR_L2Results_0__5), 
         .A0 (CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx554), .A1 (
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx558)) ;
    aoi22 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix555 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx554), .A0 (
          CALCULATOR_L1Results_0__4), .A1 (CALCULATOR_L1Results_1__4), .B0 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx48), .B1 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx12)) ;
    xnor2 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix559 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx558), .A0 (
          CALCULATOR_L1Results_1__5), .A1 (CALCULATOR_L1Results_0__5)) ;
    xor2 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix67 (.Y (CALCULATOR_L2Results_0__6), 
         .A0 (CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx561), .A1 (
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx565)) ;
    aoi22 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix562 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx561), .A0 (
          CALCULATOR_L1Results_0__5), .A1 (CALCULATOR_L1Results_1__5), .B0 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx52), .B1 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx6)) ;
    xnor2 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix566 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx565), .A0 (
          CALCULATOR_L1Results_1__6), .A1 (CALCULATOR_L1Results_0__6)) ;
    xnor2 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix65 (.Y (CALCULATOR_L2Results_0__7)
          , .A0 (CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx568), .A1 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx62)) ;
    aoi22 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix569 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx568), .A0 (
          CALCULATOR_L1Results_0__6), .A1 (CALCULATOR_L1Results_1__6), .B0 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx56), .B1 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx0)) ;
    xor2 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix63 (.Y (
         CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx62), .A0 (CALCULATOR_L1Results_1__7)
         , .A1 (CALCULATOR_L1Results_0__7)) ;
    inv01 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix155 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx154), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx383)) ;
    inv01 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix57 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx56), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx561)) ;
    inv01 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix53 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx52), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx554)) ;
    inv01 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix49 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx48), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx547)) ;
    inv01 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix45 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx44), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx540)) ;
    inv01 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix41 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx40), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx534)) ;
    inv01 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix31 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx30), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx531)) ;
    inv01 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix25 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx24), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx537)) ;
    inv01 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix19 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx18), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx544)) ;
    inv01 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix13 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx12), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx551)) ;
    inv01 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix7 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx6), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx558)) ;
    inv01 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix1 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx0), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx565)) ;
    fake_gnd CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix216 (.Y (
             CALCULATOR_L1_2_L2_3_G2_MINI_ALU_WindowCellShiftedLeft_16)) ;
    aoi21 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix77 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_10), .A0 (
          CacheFilter_2__3__1), .A1 (CacheFilter_2__3__0), .B0 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx4)) ;
    nor02_2x CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix5 (.Y (
             CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx4), .A0 (
             CacheFilter_2__3__0), .A1 (CacheFilter_2__3__1)) ;
    aoi21 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix67 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_11), .A0 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx328), .A1 (
          CacheFilter_2__3__2), .B0 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx8)) ;
    nor03_2x CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix9 (.Y (
             CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx8), .A0 (
             CacheFilter_2__3__2), .A1 (CacheFilter_2__3__0), .A2 (
             CacheFilter_2__3__1)) ;
    xnor2 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix59 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_12), .A0 (
          CacheFilter_2__3__3), .A1 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx8)) ;
    xnor2 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix51 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_13), .A0 (
          CacheFilter_2__3__4), .A1 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx12)) ;
    nor04 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix13 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx12), .A0 (
          CacheFilter_2__3__3), .A1 (CacheFilter_2__3__2), .A2 (
          CacheFilter_2__3__0), .A3 (CacheFilter_2__3__1)) ;
    xnor2 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix43 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_14), .A0 (
          CacheFilter_2__3__5), .A1 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx16)) ;
    nor02ii CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix17 (.Y (
            CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx16), .A0 (
            CacheFilter_2__3__4), .A1 (
            CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx12)) ;
    xnor2 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix35 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_15), .A0 (
          CacheFilter_2__3__6), .A1 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx20)) ;
    nor02ii CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix21 (.Y (
            CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx20), .A0 (
            CacheFilter_2__3__5), .A1 (
            CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx16)) ;
    xnor2 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix27 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_16), .A0 (
          CacheFilter_2__3__7), .A1 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx24)) ;
    nor02ii CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix25 (.Y (
            CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx24), .A0 (
            CacheFilter_2__3__6), .A1 (
            CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx20)) ;
    inv01 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix329 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx328), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx4)) ;
    inv02 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix383 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx384), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_0)) ;
    dff CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_0 (.Q (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_0), .QB (
        \$dummy [690]), .D (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .CLK (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    nor02_2x CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix567 (.Y (
             CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566), .A0 (
             RST), .A1 (
             CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644)) ;
    dff CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_1 (.Q (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_1), .QB (
        \$dummy [691]), .D (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .CLK (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_2 (.Q (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_2), .QB (
        \$dummy [692]), .D (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .CLK (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_3 (.Q (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_3), .QB (
        \$dummy [693]), .D (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .CLK (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_4 (.Q (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_4), .QB (
        \$dummy [694]), .D (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .CLK (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_5 (.Q (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_5), .QB (
        \$dummy [695]), .D (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .CLK (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_6 (.Q (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_6), .QB (
        \$dummy [696]), .D (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .CLK (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_7 (.Q (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_7), .QB (
        \$dummy [697]), .D (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .CLK (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_8 (.Q (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_8), .QB (
        \$dummy [698]), .D (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .CLK (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_9 (.Q (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_9), .QB (
        \$dummy [699]), .D (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .CLK (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_10 (.Q (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_10), .QB (
        \$dummy [700]), .D (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .CLK (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_11 (.Q (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_11), .QB (
        \$dummy [701]), .D (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .CLK (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_12 (.Q (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_12), .QB (
        \$dummy [702]), .D (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .CLK (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_13 (.Q (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_13), .QB (
        \$dummy [703]), .D (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .CLK (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_14 (.Q (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_14), .QB (
        \$dummy [704]), .D (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .CLK (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_15 (.Q (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_15), .QB (
        \$dummy [705]), .D (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .CLK (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_16 (.Q (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_16), .QB (
        \$dummy [706]), .D (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .CLK (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    inv02 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix623 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix625 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix627 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix643 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644), .A (
          nx7899)) ;
    dff CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_0 (.Q (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_0), .QB (
        \$dummy [707]), .D (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .CLK (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    nor02_2x CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix567 (.Y (
             CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566), .A0 (
             RST), .A1 (
             CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644)) ;
    dff CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_1 (.Q (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_1), .QB (
        \$dummy [708]), .D (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .CLK (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_2 (.Q (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_2), .QB (
        \$dummy [709]), .D (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .CLK (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_3 (.Q (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_3), .QB (
        \$dummy [710]), .D (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .CLK (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_4 (.Q (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_4), .QB (
        \$dummy [711]), .D (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .CLK (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_5 (.Q (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_5), .QB (
        \$dummy [712]), .D (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .CLK (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_6 (.Q (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_6), .QB (
        \$dummy [713]), .D (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .CLK (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_7 (.Q (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_7), .QB (
        \$dummy [714]), .D (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .CLK (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_8 (.Q (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_8), .QB (
        \$dummy [715]), .D (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .CLK (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_9 (.Q (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_9), .QB (
        \$dummy [716]), .D (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .CLK (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_10 (.Q (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_10), .QB (
        \$dummy [717]), .D (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .CLK (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_11 (.Q (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_11), .QB (
        \$dummy [718]), .D (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .CLK (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_12 (.Q (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_12), .QB (
        \$dummy [719]), .D (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .CLK (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_13 (.Q (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_13), .QB (
        \$dummy [720]), .D (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .CLK (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_14 (.Q (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_14), .QB (
        \$dummy [721]), .D (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .CLK (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_15 (.Q (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_15), .QB (
        \$dummy [722]), .D (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .CLK (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_16 (.Q (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_16), .QB (
        \$dummy [723]), .D (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .CLK (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    inv02 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix623 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix625 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix627 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix643 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644), .A (
          nx7905)) ;
    dff CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_0 (.Q (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_0), .QB (\$dummy [724]), .D (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .CLK (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    nor02_2x CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix567 (.Y (
             CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566), .A0 (
             RST), .A1 (
             CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    dff CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_1 (.Q (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_1), .QB (\$dummy [725]), .D (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .CLK (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_2 (.Q (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_2), .QB (\$dummy [726]), .D (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .CLK (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_3 (.Q (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_3), .QB (\$dummy [727]), .D (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .CLK (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_4 (.Q (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_4), .QB (\$dummy [728]), .D (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .CLK (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_5 (.Q (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_5), .QB (\$dummy [729]), .D (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .CLK (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_6 (.Q (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_6), .QB (\$dummy [730]), .D (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .CLK (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_7 (.Q (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_7), .QB (\$dummy [731]), .D (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .CLK (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_8 (.Q (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_8), .QB (\$dummy [732]), .D (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .CLK (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_9 (.Q (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_9), .QB (\$dummy [733]), .D (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .CLK (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_10 (.Q (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_10), .QB (\$dummy [734]), .D (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .CLK (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_11 (.Q (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_11), .QB (\$dummy [735]), .D (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .CLK (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_12 (.Q (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_12), .QB (\$dummy [736]), .D (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .CLK (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_13 (.Q (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_13), .QB (\$dummy [737]), .D (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .CLK (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_14 (.Q (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_14), .QB (\$dummy [738]), .D (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .CLK (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_15 (.Q (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_15), .QB (\$dummy [739]), .D (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .CLK (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_16 (.Q (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_16), .QB (\$dummy [740]), .D (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .CLK (
        CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    inv02 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix623 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix625 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix627 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix643 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642)) ;
    xor2 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix83 (.Y (CALCULATOR_L2Results_1__0), 
         .A0 (CALCULATOR_L1Results_3__0), .A1 (CALCULATOR_L1Results_2__0)) ;
    xnor2 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix380 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx379), .A0 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx381), .A1 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx383)) ;
    nand02 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix382 (.Y (
           CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx381), .A0 (
           CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothOperand_0), .A1 (nx7925)) ;
    xnor2 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix384 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx383), .A0 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothOperand_1), .A1 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_1)) ;
    inv01 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix388 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx387), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_2)) ;
    xnor2 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix390 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx389), .A0 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx391), .A1 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx395)) ;
    aoi32 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix392 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx391), .A0 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothOperand_0), .A1 (nx7925), .A2 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx154), .B0 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_1), .B1 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothOperand_1)) ;
    xnor2 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix396 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx395), .A0 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothOperand_2), .A1 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_2)) ;
    inv01 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix400 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx399), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_3)) ;
    xnor2 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix402 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx401), .A0 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx403), .A1 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx405)) ;
    xnor2 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix406 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx405), .A0 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothOperand_3), .A1 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_3)) ;
    inv01 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix410 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx409), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_4)) ;
    xnor2 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix412 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx411), .A0 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx413), .A1 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx415)) ;
    xnor2 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix416 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx415), .A0 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothOperand_4), .A1 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_4)) ;
    inv01 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix420 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx419), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_5)) ;
    xnor2 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix422 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx421), .A0 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx423), .A1 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx425)) ;
    xnor2 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix426 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx425), .A0 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothOperand_5), .A1 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_5)) ;
    inv01 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix430 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx429), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_6)) ;
    xnor2 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix432 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx431), .A0 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx433), .A1 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx435)) ;
    xnor2 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix436 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx435), .A0 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothOperand_6), .A1 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_6)) ;
    inv01 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix440 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx439), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_7)) ;
    xnor2 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix442 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx441), .A0 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx443), .A1 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx445)) ;
    xnor2 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix446 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx445), .A0 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothOperand_7), .A1 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_7)) ;
    inv01 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix450 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx449), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_8)) ;
    xnor2 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix452 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx451), .A0 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx453), .A1 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx455)) ;
    xnor2 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix456 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx455), .A0 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothOperand_8), .A1 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_8)) ;
    xor2 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix317 (.Y (
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx316), .A0 (
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx461), .A1 (
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx463)) ;
    xnor2 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix464 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx463), .A0 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothOperand_9), .A1 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_9)) ;
    xor2 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix337 (.Y (
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx336), .A0 (
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx467), .A1 (
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx471)) ;
    inv01 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix470 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx469), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_9)) ;
    xnor2 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix472 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx471), .A0 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothOperand_10), .A1 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_10)) ;
    xor2 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix357 (.Y (
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx356), .A0 (
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx475), .A1 (
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx479)) ;
    inv01 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix478 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx477), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_10)) ;
    xnor2 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix480 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx479), .A0 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothOperand_11), .A1 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_11)) ;
    xor2 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix377 (.Y (
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx376), .A0 (
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx483), .A1 (
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx487)) ;
    inv01 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix486 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx485), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_11)) ;
    xnor2 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix488 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx487), .A0 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothOperand_12), .A1 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_12)) ;
    xor2 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix397 (.Y (
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx396), .A0 (
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx491), .A1 (
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx495)) ;
    inv01 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix494 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx493), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_12)) ;
    xnor2 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix496 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx495), .A0 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothOperand_13), .A1 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_13)) ;
    xor2 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix417 (.Y (
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx416), .A0 (
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx499), .A1 (
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx503)) ;
    inv01 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix502 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx501), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_13)) ;
    xnor2 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix504 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx503), .A0 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothOperand_14), .A1 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_14)) ;
    xor2 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix437 (.Y (
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx436), .A0 (
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx507), .A1 (
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx511)) ;
    inv01 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix510 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx509), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_14)) ;
    xnor2 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix512 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx511), .A0 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothOperand_15), .A1 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_15)) ;
    xnor2 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix457 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx456), .A0 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx515), .A1 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx454)) ;
    inv01 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix518 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx517), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_15)) ;
    xor2 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix455 (.Y (
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx454), .A0 (
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothOperand_16), .A1 (
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_16)) ;
    mux21_ni CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix91 (.Y (
             CALCULATOR_L1FirstOperands_2__0), .A0 (
             CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_1), .A1 (
             CacheWindow_2__4__0), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix99 (.Y (
             CALCULATOR_L1FirstOperands_2__1), .A0 (
             CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_2), .A1 (
             CacheWindow_2__4__1), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix107 (.Y (
             CALCULATOR_L1FirstOperands_2__2), .A0 (
             CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_3), .A1 (
             CacheWindow_2__4__2), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix115 (.Y (
             CALCULATOR_L1FirstOperands_2__3), .A0 (
             CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_4), .A1 (
             CacheWindow_2__4__3), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix123 (.Y (
             CALCULATOR_L1FirstOperands_2__4), .A0 (
             CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_5), .A1 (
             CacheWindow_2__4__4), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix131 (.Y (
             CALCULATOR_L1FirstOperands_2__5), .A0 (
             CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_6), .A1 (
             CacheWindow_2__4__5), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix139 (.Y (
             CALCULATOR_L1FirstOperands_2__6), .A0 (
             CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_7), .A1 (
             CacheWindow_2__4__6), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix147 (.Y (
             CALCULATOR_L1FirstOperands_2__7), .A0 (
             CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_8), .A1 (
             CacheWindow_2__4__7), .S0 (Instr)) ;
    xor2 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix77 (.Y (CALCULATOR_L2Results_1__1), 
         .A0 (CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx529), .A1 (
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx531)) ;
    nand02 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix530 (.Y (
           CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx529), .A0 (
           CALCULATOR_L1Results_3__0), .A1 (CALCULATOR_L1Results_2__0)) ;
    xnor2 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix532 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx531), .A0 (
          CALCULATOR_L1Results_3__1), .A1 (CALCULATOR_L1Results_2__1)) ;
    xor2 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix75 (.Y (CALCULATOR_L2Results_1__2), 
         .A0 (CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx534), .A1 (
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx537)) ;
    aoi32 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix535 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx534), .A0 (
          CALCULATOR_L1Results_3__0), .A1 (CALCULATOR_L1Results_2__0), .A2 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx30), .B0 (CALCULATOR_L1Results_2__1
          ), .B1 (CALCULATOR_L1Results_3__1)) ;
    xnor2 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix538 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx537), .A0 (
          CALCULATOR_L1Results_3__2), .A1 (CALCULATOR_L1Results_2__2)) ;
    xor2 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix73 (.Y (CALCULATOR_L2Results_1__3), 
         .A0 (CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx540), .A1 (
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx544)) ;
    aoi22 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix541 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx540), .A0 (
          CALCULATOR_L1Results_2__2), .A1 (CALCULATOR_L1Results_3__2), .B0 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx40), .B1 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx24)) ;
    xnor2 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix545 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx544), .A0 (
          CALCULATOR_L1Results_3__3), .A1 (CALCULATOR_L1Results_2__3)) ;
    xor2 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix71 (.Y (CALCULATOR_L2Results_1__4), 
         .A0 (CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx547), .A1 (
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx551)) ;
    aoi22 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix548 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx547), .A0 (
          CALCULATOR_L1Results_2__3), .A1 (CALCULATOR_L1Results_3__3), .B0 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx44), .B1 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx18)) ;
    xnor2 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix552 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx551), .A0 (
          CALCULATOR_L1Results_3__4), .A1 (CALCULATOR_L1Results_2__4)) ;
    xor2 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix69 (.Y (CALCULATOR_L2Results_1__5), 
         .A0 (CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx554), .A1 (
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx558)) ;
    aoi22 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix555 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx554), .A0 (
          CALCULATOR_L1Results_2__4), .A1 (CALCULATOR_L1Results_3__4), .B0 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx48), .B1 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx12)) ;
    xnor2 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix559 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx558), .A0 (
          CALCULATOR_L1Results_3__5), .A1 (CALCULATOR_L1Results_2__5)) ;
    xor2 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix67 (.Y (CALCULATOR_L2Results_1__6), 
         .A0 (CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx561), .A1 (
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx565)) ;
    aoi22 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix562 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx561), .A0 (
          CALCULATOR_L1Results_2__5), .A1 (CALCULATOR_L1Results_3__5), .B0 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx52), .B1 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx6)) ;
    xnor2 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix566 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx565), .A0 (
          CALCULATOR_L1Results_3__6), .A1 (CALCULATOR_L1Results_2__6)) ;
    xnor2 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix65 (.Y (CALCULATOR_L2Results_1__7)
          , .A0 (CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx568), .A1 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx62)) ;
    aoi22 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix569 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx568), .A0 (
          CALCULATOR_L1Results_2__6), .A1 (CALCULATOR_L1Results_3__6), .B0 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx56), .B1 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx0)) ;
    xor2 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix63 (.Y (
         CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx62), .A0 (CALCULATOR_L1Results_3__7)
         , .A1 (CALCULATOR_L1Results_2__7)) ;
    inv01 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix155 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx154), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx383)) ;
    inv01 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix57 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx56), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx561)) ;
    inv01 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix53 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx52), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx554)) ;
    inv01 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix49 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx48), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx547)) ;
    inv01 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix45 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx44), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx540)) ;
    inv01 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix41 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx40), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx534)) ;
    inv01 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix31 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx30), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx531)) ;
    inv01 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix25 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx24), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx537)) ;
    inv01 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix19 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx18), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx544)) ;
    inv01 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix13 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx12), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx551)) ;
    inv01 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix7 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx6), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx558)) ;
    inv01 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix1 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx0), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx565)) ;
    fake_gnd CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix216 (.Y (
             CALCULATOR_L1_2_L2_4_G2_MINI_ALU_WindowCellShiftedLeft_16)) ;
    aoi21 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix77 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_10), .A0 (
          CacheFilter_2__4__1), .A1 (CacheFilter_2__4__0), .B0 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_nx4)) ;
    nor02_2x CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix5 (.Y (
             CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_nx4), .A0 (
             CacheFilter_2__4__0), .A1 (CacheFilter_2__4__1)) ;
    aoi21 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix67 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_11), .A0 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_nx328), .A1 (
          CacheFilter_2__4__2), .B0 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_nx8)) ;
    nor03_2x CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix9 (.Y (
             CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_nx8), .A0 (
             CacheFilter_2__4__2), .A1 (CacheFilter_2__4__0), .A2 (
             CacheFilter_2__4__1)) ;
    xnor2 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix59 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_12), .A0 (
          CacheFilter_2__4__3), .A1 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_nx8)) ;
    xnor2 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix51 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_13), .A0 (
          CacheFilter_2__4__4), .A1 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_nx12)) ;
    nor04 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix13 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_nx12), .A0 (
          CacheFilter_2__4__3), .A1 (CacheFilter_2__4__2), .A2 (
          CacheFilter_2__4__0), .A3 (CacheFilter_2__4__1)) ;
    xnor2 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix43 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_14), .A0 (
          CacheFilter_2__4__5), .A1 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_nx16)) ;
    nor02ii CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix17 (.Y (
            CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_nx16), .A0 (
            CacheFilter_2__4__4), .A1 (
            CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_nx12)) ;
    xnor2 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix35 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_15), .A0 (
          CacheFilter_2__4__6), .A1 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_nx20)) ;
    nor02ii CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix21 (.Y (
            CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_nx20), .A0 (
            CacheFilter_2__4__5), .A1 (
            CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_nx16)) ;
    xnor2 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix27 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_16), .A0 (
          CacheFilter_2__4__7), .A1 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_nx24)) ;
    nor02ii CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix25 (.Y (
            CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_nx24), .A0 (
            CacheFilter_2__4__6), .A1 (
            CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_nx20)) ;
    inv01 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix329 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_nx328), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_nx4)) ;
    inv02 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix383 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_nx384), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_0)) ;
    dff CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_0 (.Q (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_0), .QB (
        \$dummy [741]), .D (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .CLK (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    nor02_2x CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix567 (.Y (
             CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566), .A0 (
             RST), .A1 (
             CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644)) ;
    dff CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_1 (.Q (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_1), .QB (
        \$dummy [742]), .D (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .CLK (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_2 (.Q (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_2), .QB (
        \$dummy [743]), .D (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .CLK (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_3 (.Q (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_3), .QB (
        \$dummy [744]), .D (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .CLK (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_4 (.Q (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_4), .QB (
        \$dummy [745]), .D (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .CLK (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_5 (.Q (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_5), .QB (
        \$dummy [746]), .D (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .CLK (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_6 (.Q (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_6), .QB (
        \$dummy [747]), .D (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .CLK (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_7 (.Q (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_7), .QB (
        \$dummy [748]), .D (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .CLK (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_8 (.Q (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_8), .QB (
        \$dummy [749]), .D (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .CLK (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_9 (.Q (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_9), .QB (
        \$dummy [750]), .D (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .CLK (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_10 (.Q (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_10), .QB (
        \$dummy [751]), .D (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .CLK (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_11 (.Q (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_11), .QB (
        \$dummy [752]), .D (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .CLK (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_12 (.Q (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_12), .QB (
        \$dummy [753]), .D (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .CLK (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_13 (.Q (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_13), .QB (
        \$dummy [754]), .D (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .CLK (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_14 (.Q (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_14), .QB (
        \$dummy [755]), .D (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .CLK (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_15 (.Q (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_15), .QB (
        \$dummy [756]), .D (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .CLK (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_16 (.Q (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_16), .QB (
        \$dummy [757]), .D (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .CLK (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    inv02 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix623 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix625 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix627 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix643 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644), .A (
          nx7939)) ;
    dff CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_0 (.Q (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_0), .QB (
        \$dummy [758]), .D (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .CLK (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    nor02_2x CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix567 (.Y (
             CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566), .A0 (
             RST), .A1 (
             CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644)) ;
    dff CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_1 (.Q (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_1), .QB (
        \$dummy [759]), .D (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .CLK (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_2 (.Q (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_2), .QB (
        \$dummy [760]), .D (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .CLK (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_3 (.Q (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_3), .QB (
        \$dummy [761]), .D (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .CLK (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_4 (.Q (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_4), .QB (
        \$dummy [762]), .D (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .CLK (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_5 (.Q (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_5), .QB (
        \$dummy [763]), .D (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .CLK (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_6 (.Q (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_6), .QB (
        \$dummy [764]), .D (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .CLK (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_7 (.Q (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_7), .QB (
        \$dummy [765]), .D (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .CLK (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_8 (.Q (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_8), .QB (
        \$dummy [766]), .D (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .CLK (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_9 (.Q (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_9), .QB (
        \$dummy [767]), .D (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .CLK (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_10 (.Q (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_10), .QB (
        \$dummy [768]), .D (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .CLK (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_11 (.Q (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_11), .QB (
        \$dummy [769]), .D (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .CLK (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_12 (.Q (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_12), .QB (
        \$dummy [770]), .D (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .CLK (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_13 (.Q (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_13), .QB (
        \$dummy [771]), .D (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .CLK (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_14 (.Q (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_14), .QB (
        \$dummy [772]), .D (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .CLK (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_15 (.Q (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_15), .QB (
        \$dummy [773]), .D (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .CLK (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_16 (.Q (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_16), .QB (
        \$dummy [774]), .D (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .CLK (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    inv02 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix623 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix625 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix627 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix643 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644), .A (
          nx7945)) ;
    dff CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_0 (.Q (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_0), .QB (\$dummy [775]), .D (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .CLK (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    nor02_2x CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix567 (.Y (
             CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566), .A0 (
             RST), .A1 (
             CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    dff CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_1 (.Q (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_1), .QB (\$dummy [776]), .D (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .CLK (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_2 (.Q (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_2), .QB (\$dummy [777]), .D (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .CLK (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_3 (.Q (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_3), .QB (\$dummy [778]), .D (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .CLK (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_4 (.Q (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_4), .QB (\$dummy [779]), .D (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .CLK (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_5 (.Q (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_5), .QB (\$dummy [780]), .D (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .CLK (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_6 (.Q (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_6), .QB (\$dummy [781]), .D (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .CLK (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_7 (.Q (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_7), .QB (\$dummy [782]), .D (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .CLK (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_8 (.Q (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_8), .QB (\$dummy [783]), .D (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .CLK (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_9 (.Q (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_9), .QB (\$dummy [784]), .D (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .CLK (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_10 (.Q (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_10), .QB (\$dummy [785]), .D (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .CLK (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_11 (.Q (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_11), .QB (\$dummy [786]), .D (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .CLK (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_12 (.Q (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_12), .QB (\$dummy [787]), .D (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .CLK (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_13 (.Q (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_13), .QB (\$dummy [788]), .D (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .CLK (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_14 (.Q (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_14), .QB (\$dummy [789]), .D (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .CLK (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_15 (.Q (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_15), .QB (\$dummy [790]), .D (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .CLK (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_16 (.Q (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_16), .QB (\$dummy [791]), .D (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .CLK (
        CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    inv02 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix623 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix625 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix627 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix643 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642)) ;
    xor2 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix83 (.Y (CALCULATOR_L2Results_2__0), 
         .A0 (CALCULATOR_L1Results_5__0), .A1 (CALCULATOR_L1Results_4__0)) ;
    xnor2 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix380 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx379), .A0 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx381), .A1 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx383)) ;
    nand02 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix382 (.Y (
           CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx381), .A0 (
           CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothOperand_0), .A1 (nx7965)) ;
    xnor2 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix384 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx383), .A0 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothOperand_1), .A1 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_1)) ;
    inv01 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix388 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx387), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_2)) ;
    xnor2 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix390 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx389), .A0 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx391), .A1 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx395)) ;
    aoi32 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix392 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx391), .A0 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothOperand_0), .A1 (nx7965), .A2 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx154), .B0 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_1), .B1 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothOperand_1)) ;
    xnor2 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix396 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx395), .A0 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothOperand_2), .A1 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_2)) ;
    inv01 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix400 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx399), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_3)) ;
    xnor2 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix402 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx401), .A0 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx403), .A1 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx405)) ;
    xnor2 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix406 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx405), .A0 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothOperand_3), .A1 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_3)) ;
    inv01 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix410 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx409), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_4)) ;
    xnor2 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix412 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx411), .A0 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx413), .A1 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx415)) ;
    xnor2 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix416 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx415), .A0 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothOperand_4), .A1 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_4)) ;
    inv01 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix420 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx419), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_5)) ;
    xnor2 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix422 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx421), .A0 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx423), .A1 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx425)) ;
    xnor2 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix426 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx425), .A0 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothOperand_5), .A1 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_5)) ;
    inv01 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix430 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx429), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_6)) ;
    xnor2 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix432 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx431), .A0 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx433), .A1 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx435)) ;
    xnor2 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix436 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx435), .A0 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothOperand_6), .A1 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_6)) ;
    inv01 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix440 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx439), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_7)) ;
    xnor2 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix442 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx441), .A0 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx443), .A1 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx445)) ;
    xnor2 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix446 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx445), .A0 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothOperand_7), .A1 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_7)) ;
    inv01 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix450 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx449), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_8)) ;
    xnor2 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix452 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx451), .A0 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx453), .A1 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx455)) ;
    xnor2 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix456 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx455), .A0 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothOperand_8), .A1 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_8)) ;
    xor2 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix317 (.Y (
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx316), .A0 (
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx461), .A1 (
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx463)) ;
    xnor2 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix464 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx463), .A0 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothOperand_9), .A1 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_9)) ;
    xor2 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix337 (.Y (
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx336), .A0 (
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx467), .A1 (
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx471)) ;
    inv01 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix470 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx469), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_9)) ;
    xnor2 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix472 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx471), .A0 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothOperand_10), .A1 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_10)) ;
    xor2 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix357 (.Y (
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx356), .A0 (
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx475), .A1 (
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx479)) ;
    inv01 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix478 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx477), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_10)) ;
    xnor2 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix480 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx479), .A0 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothOperand_11), .A1 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_11)) ;
    xor2 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix377 (.Y (
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx376), .A0 (
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx483), .A1 (
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx487)) ;
    inv01 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix486 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx485), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_11)) ;
    xnor2 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix488 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx487), .A0 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothOperand_12), .A1 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_12)) ;
    xor2 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix397 (.Y (
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx396), .A0 (
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx491), .A1 (
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx495)) ;
    inv01 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix494 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx493), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_12)) ;
    xnor2 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix496 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx495), .A0 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothOperand_13), .A1 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_13)) ;
    xor2 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix417 (.Y (
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx416), .A0 (
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx499), .A1 (
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx503)) ;
    inv01 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix502 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx501), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_13)) ;
    xnor2 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix504 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx503), .A0 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothOperand_14), .A1 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_14)) ;
    xor2 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix437 (.Y (
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx436), .A0 (
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx507), .A1 (
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx511)) ;
    inv01 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix510 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx509), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_14)) ;
    xnor2 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix512 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx511), .A0 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothOperand_15), .A1 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_15)) ;
    xnor2 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix457 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx456), .A0 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx515), .A1 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx454)) ;
    inv01 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix518 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx517), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_15)) ;
    xor2 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix455 (.Y (
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx454), .A0 (
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothOperand_16), .A1 (
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_16)) ;
    mux21_ni CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix91 (.Y (
             CALCULATOR_L1FirstOperands_4__0), .A0 (
             CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_1), .A1 (
             CacheWindow_3__0__0), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix99 (.Y (
             CALCULATOR_L1FirstOperands_4__1), .A0 (
             CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_2), .A1 (
             CacheWindow_3__0__1), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix107 (.Y (
             CALCULATOR_L1FirstOperands_4__2), .A0 (
             CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_3), .A1 (
             CacheWindow_3__0__2), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix115 (.Y (
             CALCULATOR_L1FirstOperands_4__3), .A0 (
             CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_4), .A1 (
             CacheWindow_3__0__3), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix123 (.Y (
             CALCULATOR_L1FirstOperands_4__4), .A0 (
             CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_5), .A1 (
             CacheWindow_3__0__4), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix131 (.Y (
             CALCULATOR_L1FirstOperands_4__5), .A0 (
             CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_6), .A1 (
             CacheWindow_3__0__5), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix139 (.Y (
             CALCULATOR_L1FirstOperands_4__6), .A0 (
             CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_7), .A1 (
             CacheWindow_3__0__6), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix147 (.Y (
             CALCULATOR_L1FirstOperands_4__7), .A0 (
             CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_8), .A1 (
             CacheWindow_3__0__7), .S0 (Instr)) ;
    xor2 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix77 (.Y (CALCULATOR_L2Results_2__1), 
         .A0 (CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx529), .A1 (
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx531)) ;
    nand02 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix530 (.Y (
           CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx529), .A0 (
           CALCULATOR_L1Results_5__0), .A1 (CALCULATOR_L1Results_4__0)) ;
    xnor2 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix532 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx531), .A0 (
          CALCULATOR_L1Results_5__1), .A1 (CALCULATOR_L1Results_4__1)) ;
    xor2 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix75 (.Y (CALCULATOR_L2Results_2__2), 
         .A0 (CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx534), .A1 (
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx537)) ;
    aoi32 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix535 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx534), .A0 (
          CALCULATOR_L1Results_5__0), .A1 (CALCULATOR_L1Results_4__0), .A2 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx30), .B0 (CALCULATOR_L1Results_4__1
          ), .B1 (CALCULATOR_L1Results_5__1)) ;
    xnor2 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix538 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx537), .A0 (
          CALCULATOR_L1Results_5__2), .A1 (CALCULATOR_L1Results_4__2)) ;
    xor2 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix73 (.Y (CALCULATOR_L2Results_2__3), 
         .A0 (CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx540), .A1 (
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx544)) ;
    aoi22 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix541 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx540), .A0 (
          CALCULATOR_L1Results_4__2), .A1 (CALCULATOR_L1Results_5__2), .B0 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx40), .B1 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx24)) ;
    xnor2 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix545 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx544), .A0 (
          CALCULATOR_L1Results_5__3), .A1 (CALCULATOR_L1Results_4__3)) ;
    xor2 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix71 (.Y (CALCULATOR_L2Results_2__4), 
         .A0 (CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx547), .A1 (
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx551)) ;
    aoi22 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix548 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx547), .A0 (
          CALCULATOR_L1Results_4__3), .A1 (CALCULATOR_L1Results_5__3), .B0 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx44), .B1 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx18)) ;
    xnor2 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix552 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx551), .A0 (
          CALCULATOR_L1Results_5__4), .A1 (CALCULATOR_L1Results_4__4)) ;
    xor2 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix69 (.Y (CALCULATOR_L2Results_2__5), 
         .A0 (CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx554), .A1 (
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx558)) ;
    aoi22 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix555 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx554), .A0 (
          CALCULATOR_L1Results_4__4), .A1 (CALCULATOR_L1Results_5__4), .B0 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx48), .B1 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx12)) ;
    xnor2 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix559 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx558), .A0 (
          CALCULATOR_L1Results_5__5), .A1 (CALCULATOR_L1Results_4__5)) ;
    xor2 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix67 (.Y (CALCULATOR_L2Results_2__6), 
         .A0 (CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx561), .A1 (
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx565)) ;
    aoi22 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix562 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx561), .A0 (
          CALCULATOR_L1Results_4__5), .A1 (CALCULATOR_L1Results_5__5), .B0 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx52), .B1 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx6)) ;
    xnor2 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix566 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx565), .A0 (
          CALCULATOR_L1Results_5__6), .A1 (CALCULATOR_L1Results_4__6)) ;
    xnor2 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix65 (.Y (CALCULATOR_L2Results_2__7)
          , .A0 (CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx568), .A1 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx62)) ;
    aoi22 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix569 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx568), .A0 (
          CALCULATOR_L1Results_4__6), .A1 (CALCULATOR_L1Results_5__6), .B0 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx56), .B1 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx0)) ;
    xor2 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix63 (.Y (
         CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx62), .A0 (CALCULATOR_L1Results_5__7)
         , .A1 (CALCULATOR_L1Results_4__7)) ;
    inv01 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix155 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx154), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx383)) ;
    inv01 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix57 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx56), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx561)) ;
    inv01 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix53 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx52), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx554)) ;
    inv01 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix49 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx48), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx547)) ;
    inv01 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix45 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx44), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx540)) ;
    inv01 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix41 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx40), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx534)) ;
    inv01 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix31 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx30), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx531)) ;
    inv01 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix25 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx24), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx537)) ;
    inv01 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix19 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx18), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx544)) ;
    inv01 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix13 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx12), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx551)) ;
    inv01 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix7 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx6), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx558)) ;
    inv01 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix1 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx0), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx565)) ;
    fake_gnd CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix216 (.Y (
             CALCULATOR_L1_3_L2_0_G2_MINI_ALU_WindowCellShiftedLeft_16)) ;
    aoi21 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix77 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_10), .A0 (
          CacheFilter_3__0__1), .A1 (CacheFilter_3__0__0), .B0 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_nx4)) ;
    nor02_2x CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix5 (.Y (
             CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_nx4), .A0 (
             CacheFilter_3__0__0), .A1 (CacheFilter_3__0__1)) ;
    aoi21 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix67 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_11), .A0 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_nx328), .A1 (
          CacheFilter_3__0__2), .B0 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_nx8)) ;
    nor03_2x CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix9 (.Y (
             CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_nx8), .A0 (
             CacheFilter_3__0__2), .A1 (CacheFilter_3__0__0), .A2 (
             CacheFilter_3__0__1)) ;
    xnor2 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix59 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_12), .A0 (
          CacheFilter_3__0__3), .A1 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_nx8)) ;
    xnor2 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix51 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_13), .A0 (
          CacheFilter_3__0__4), .A1 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_nx12)) ;
    nor04 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix13 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_nx12), .A0 (
          CacheFilter_3__0__3), .A1 (CacheFilter_3__0__2), .A2 (
          CacheFilter_3__0__0), .A3 (CacheFilter_3__0__1)) ;
    xnor2 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix43 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_14), .A0 (
          CacheFilter_3__0__5), .A1 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_nx16)) ;
    nor02ii CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix17 (.Y (
            CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_nx16), .A0 (
            CacheFilter_3__0__4), .A1 (
            CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_nx12)) ;
    xnor2 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix35 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_15), .A0 (
          CacheFilter_3__0__6), .A1 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_nx20)) ;
    nor02ii CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix21 (.Y (
            CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_nx20), .A0 (
            CacheFilter_3__0__5), .A1 (
            CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_nx16)) ;
    xnor2 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix27 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_16), .A0 (
          CacheFilter_3__0__7), .A1 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_nx24)) ;
    nor02ii CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix25 (.Y (
            CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_nx24), .A0 (
            CacheFilter_3__0__6), .A1 (
            CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_nx20)) ;
    inv01 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix329 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_nx328), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_nx4)) ;
    inv02 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix383 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_nx384), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_0)) ;
    dff CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_0 (.Q (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_0), .QB (
        \$dummy [792]), .D (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .CLK (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    nor02_2x CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix567 (.Y (
             CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566), .A0 (
             RST), .A1 (
             CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644)) ;
    dff CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_1 (.Q (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_1), .QB (
        \$dummy [793]), .D (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .CLK (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_2 (.Q (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_2), .QB (
        \$dummy [794]), .D (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .CLK (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_3 (.Q (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_3), .QB (
        \$dummy [795]), .D (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .CLK (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_4 (.Q (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_4), .QB (
        \$dummy [796]), .D (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .CLK (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_5 (.Q (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_5), .QB (
        \$dummy [797]), .D (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .CLK (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_6 (.Q (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_6), .QB (
        \$dummy [798]), .D (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .CLK (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_7 (.Q (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_7), .QB (
        \$dummy [799]), .D (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .CLK (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_8 (.Q (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_8), .QB (
        \$dummy [800]), .D (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .CLK (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_9 (.Q (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_9), .QB (
        \$dummy [801]), .D (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .CLK (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_10 (.Q (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_10), .QB (
        \$dummy [802]), .D (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .CLK (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_11 (.Q (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_11), .QB (
        \$dummy [803]), .D (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .CLK (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_12 (.Q (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_12), .QB (
        \$dummy [804]), .D (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .CLK (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_13 (.Q (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_13), .QB (
        \$dummy [805]), .D (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .CLK (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_14 (.Q (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_14), .QB (
        \$dummy [806]), .D (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .CLK (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_15 (.Q (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_15), .QB (
        \$dummy [807]), .D (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .CLK (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_16 (.Q (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_16), .QB (
        \$dummy [808]), .D (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .CLK (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    inv02 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix623 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix625 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix627 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix643 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644), .A (
          nx7979)) ;
    dff CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_0 (.Q (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_0), .QB (
        \$dummy [809]), .D (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .CLK (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    nor02_2x CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix567 (.Y (
             CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566), .A0 (
             RST), .A1 (
             CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644)) ;
    dff CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_1 (.Q (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_1), .QB (
        \$dummy [810]), .D (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .CLK (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_2 (.Q (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_2), .QB (
        \$dummy [811]), .D (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .CLK (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_3 (.Q (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_3), .QB (
        \$dummy [812]), .D (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .CLK (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_4 (.Q (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_4), .QB (
        \$dummy [813]), .D (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .CLK (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_5 (.Q (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_5), .QB (
        \$dummy [814]), .D (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .CLK (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_6 (.Q (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_6), .QB (
        \$dummy [815]), .D (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .CLK (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_7 (.Q (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_7), .QB (
        \$dummy [816]), .D (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .CLK (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_8 (.Q (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_8), .QB (
        \$dummy [817]), .D (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .CLK (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_9 (.Q (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_9), .QB (
        \$dummy [818]), .D (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .CLK (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_10 (.Q (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_10), .QB (
        \$dummy [819]), .D (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .CLK (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_11 (.Q (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_11), .QB (
        \$dummy [820]), .D (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .CLK (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_12 (.Q (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_12), .QB (
        \$dummy [821]), .D (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .CLK (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_13 (.Q (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_13), .QB (
        \$dummy [822]), .D (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .CLK (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_14 (.Q (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_14), .QB (
        \$dummy [823]), .D (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .CLK (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_15 (.Q (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_15), .QB (
        \$dummy [824]), .D (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .CLK (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_16 (.Q (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_16), .QB (
        \$dummy [825]), .D (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .CLK (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    inv02 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix623 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix625 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix627 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix643 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644), .A (
          nx7985)) ;
    dff CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_0 (.Q (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_0), .QB (\$dummy [826]), .D (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .CLK (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    nor02_2x CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix567 (.Y (
             CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566), .A0 (
             RST), .A1 (
             CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    dff CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_1 (.Q (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_1), .QB (\$dummy [827]), .D (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .CLK (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_2 (.Q (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_2), .QB (\$dummy [828]), .D (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .CLK (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_3 (.Q (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_3), .QB (\$dummy [829]), .D (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .CLK (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_4 (.Q (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_4), .QB (\$dummy [830]), .D (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .CLK (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_5 (.Q (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_5), .QB (\$dummy [831]), .D (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .CLK (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_6 (.Q (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_6), .QB (\$dummy [832]), .D (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .CLK (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_7 (.Q (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_7), .QB (\$dummy [833]), .D (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .CLK (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_8 (.Q (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_8), .QB (\$dummy [834]), .D (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .CLK (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_9 (.Q (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_9), .QB (\$dummy [835]), .D (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .CLK (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_10 (.Q (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_10), .QB (\$dummy [836]), .D (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .CLK (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_11 (.Q (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_11), .QB (\$dummy [837]), .D (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .CLK (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_12 (.Q (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_12), .QB (\$dummy [838]), .D (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .CLK (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_13 (.Q (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_13), .QB (\$dummy [839]), .D (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .CLK (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_14 (.Q (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_14), .QB (\$dummy [840]), .D (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .CLK (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_15 (.Q (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_15), .QB (\$dummy [841]), .D (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .CLK (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_16 (.Q (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_16), .QB (\$dummy [842]), .D (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .CLK (
        CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    inv02 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix623 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix625 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix627 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix643 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642)) ;
    xor2 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix83 (.Y (CALCULATOR_L2Results_3__0), 
         .A0 (CALCULATOR_L1Results_7__0), .A1 (CALCULATOR_L1Results_6__0)) ;
    xnor2 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix380 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx379), .A0 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx381), .A1 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx383)) ;
    nand02 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix382 (.Y (
           CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx381), .A0 (
           CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothOperand_0), .A1 (nx8005)) ;
    xnor2 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix384 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx383), .A0 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothOperand_1), .A1 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_1)) ;
    inv01 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix388 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx387), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_2)) ;
    xnor2 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix390 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx389), .A0 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx391), .A1 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx395)) ;
    aoi32 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix392 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx391), .A0 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothOperand_0), .A1 (nx8005), .A2 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx154), .B0 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_1), .B1 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothOperand_1)) ;
    xnor2 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix396 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx395), .A0 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothOperand_2), .A1 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_2)) ;
    inv01 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix400 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx399), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_3)) ;
    xnor2 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix402 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx401), .A0 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx403), .A1 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx405)) ;
    xnor2 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix406 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx405), .A0 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothOperand_3), .A1 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_3)) ;
    inv01 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix410 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx409), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_4)) ;
    xnor2 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix412 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx411), .A0 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx413), .A1 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx415)) ;
    xnor2 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix416 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx415), .A0 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothOperand_4), .A1 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_4)) ;
    inv01 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix420 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx419), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_5)) ;
    xnor2 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix422 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx421), .A0 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx423), .A1 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx425)) ;
    xnor2 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix426 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx425), .A0 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothOperand_5), .A1 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_5)) ;
    inv01 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix430 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx429), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_6)) ;
    xnor2 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix432 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx431), .A0 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx433), .A1 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx435)) ;
    xnor2 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix436 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx435), .A0 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothOperand_6), .A1 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_6)) ;
    inv01 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix440 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx439), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_7)) ;
    xnor2 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix442 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx441), .A0 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx443), .A1 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx445)) ;
    xnor2 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix446 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx445), .A0 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothOperand_7), .A1 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_7)) ;
    inv01 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix450 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx449), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_8)) ;
    xnor2 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix452 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx451), .A0 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx453), .A1 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx455)) ;
    xnor2 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix456 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx455), .A0 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothOperand_8), .A1 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_8)) ;
    xor2 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix317 (.Y (
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx316), .A0 (
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx461), .A1 (
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx463)) ;
    xnor2 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix464 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx463), .A0 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothOperand_9), .A1 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_9)) ;
    xor2 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix337 (.Y (
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx336), .A0 (
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx467), .A1 (
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx471)) ;
    inv01 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix470 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx469), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_9)) ;
    xnor2 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix472 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx471), .A0 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothOperand_10), .A1 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_10)) ;
    xor2 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix357 (.Y (
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx356), .A0 (
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx475), .A1 (
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx479)) ;
    inv01 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix478 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx477), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_10)) ;
    xnor2 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix480 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx479), .A0 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothOperand_11), .A1 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_11)) ;
    xor2 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix377 (.Y (
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx376), .A0 (
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx483), .A1 (
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx487)) ;
    inv01 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix486 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx485), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_11)) ;
    xnor2 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix488 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx487), .A0 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothOperand_12), .A1 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_12)) ;
    xor2 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix397 (.Y (
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx396), .A0 (
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx491), .A1 (
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx495)) ;
    inv01 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix494 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx493), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_12)) ;
    xnor2 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix496 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx495), .A0 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothOperand_13), .A1 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_13)) ;
    xor2 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix417 (.Y (
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx416), .A0 (
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx499), .A1 (
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx503)) ;
    inv01 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix502 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx501), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_13)) ;
    xnor2 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix504 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx503), .A0 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothOperand_14), .A1 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_14)) ;
    xor2 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix437 (.Y (
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx436), .A0 (
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx507), .A1 (
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx511)) ;
    inv01 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix510 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx509), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_14)) ;
    xnor2 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix512 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx511), .A0 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothOperand_15), .A1 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_15)) ;
    xnor2 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix457 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx456), .A0 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx515), .A1 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx454)) ;
    inv01 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix518 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx517), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_15)) ;
    xor2 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix455 (.Y (
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx454), .A0 (
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothOperand_16), .A1 (
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_16)) ;
    mux21_ni CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix91 (.Y (
             CALCULATOR_L1FirstOperands_6__0), .A0 (
             CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_1), .A1 (
             CacheWindow_3__1__0), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix99 (.Y (
             CALCULATOR_L1FirstOperands_6__1), .A0 (
             CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_2), .A1 (
             CacheWindow_3__1__1), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix107 (.Y (
             CALCULATOR_L1FirstOperands_6__2), .A0 (
             CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_3), .A1 (
             CacheWindow_3__1__2), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix115 (.Y (
             CALCULATOR_L1FirstOperands_6__3), .A0 (
             CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_4), .A1 (
             CacheWindow_3__1__3), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix123 (.Y (
             CALCULATOR_L1FirstOperands_6__4), .A0 (
             CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_5), .A1 (
             CacheWindow_3__1__4), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix131 (.Y (
             CALCULATOR_L1FirstOperands_6__5), .A0 (
             CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_6), .A1 (
             CacheWindow_3__1__5), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix139 (.Y (
             CALCULATOR_L1FirstOperands_6__6), .A0 (
             CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_7), .A1 (
             CacheWindow_3__1__6), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix147 (.Y (
             CALCULATOR_L1FirstOperands_6__7), .A0 (
             CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_8), .A1 (
             CacheWindow_3__1__7), .S0 (Instr)) ;
    xor2 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix77 (.Y (CALCULATOR_L2Results_3__1), 
         .A0 (CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx529), .A1 (
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx531)) ;
    nand02 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix530 (.Y (
           CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx529), .A0 (
           CALCULATOR_L1Results_7__0), .A1 (CALCULATOR_L1Results_6__0)) ;
    xnor2 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix532 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx531), .A0 (
          CALCULATOR_L1Results_7__1), .A1 (CALCULATOR_L1Results_6__1)) ;
    xor2 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix75 (.Y (CALCULATOR_L2Results_3__2), 
         .A0 (CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx534), .A1 (
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx537)) ;
    aoi32 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix535 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx534), .A0 (
          CALCULATOR_L1Results_7__0), .A1 (CALCULATOR_L1Results_6__0), .A2 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx30), .B0 (CALCULATOR_L1Results_6__1
          ), .B1 (CALCULATOR_L1Results_7__1)) ;
    xnor2 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix538 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx537), .A0 (
          CALCULATOR_L1Results_7__2), .A1 (CALCULATOR_L1Results_6__2)) ;
    xor2 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix73 (.Y (CALCULATOR_L2Results_3__3), 
         .A0 (CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx540), .A1 (
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx544)) ;
    aoi22 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix541 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx540), .A0 (
          CALCULATOR_L1Results_6__2), .A1 (CALCULATOR_L1Results_7__2), .B0 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx40), .B1 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx24)) ;
    xnor2 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix545 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx544), .A0 (
          CALCULATOR_L1Results_7__3), .A1 (CALCULATOR_L1Results_6__3)) ;
    xor2 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix71 (.Y (CALCULATOR_L2Results_3__4), 
         .A0 (CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx547), .A1 (
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx551)) ;
    aoi22 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix548 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx547), .A0 (
          CALCULATOR_L1Results_6__3), .A1 (CALCULATOR_L1Results_7__3), .B0 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx44), .B1 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx18)) ;
    xnor2 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix552 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx551), .A0 (
          CALCULATOR_L1Results_7__4), .A1 (CALCULATOR_L1Results_6__4)) ;
    xor2 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix69 (.Y (CALCULATOR_L2Results_3__5), 
         .A0 (CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx554), .A1 (
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx558)) ;
    aoi22 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix555 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx554), .A0 (
          CALCULATOR_L1Results_6__4), .A1 (CALCULATOR_L1Results_7__4), .B0 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx48), .B1 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx12)) ;
    xnor2 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix559 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx558), .A0 (
          CALCULATOR_L1Results_7__5), .A1 (CALCULATOR_L1Results_6__5)) ;
    xor2 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix67 (.Y (CALCULATOR_L2Results_3__6), 
         .A0 (CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx561), .A1 (
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx565)) ;
    aoi22 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix562 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx561), .A0 (
          CALCULATOR_L1Results_6__5), .A1 (CALCULATOR_L1Results_7__5), .B0 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx52), .B1 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx6)) ;
    xnor2 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix566 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx565), .A0 (
          CALCULATOR_L1Results_7__6), .A1 (CALCULATOR_L1Results_6__6)) ;
    xnor2 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix65 (.Y (CALCULATOR_L2Results_3__7)
          , .A0 (CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx568), .A1 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx62)) ;
    aoi22 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix569 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx568), .A0 (
          CALCULATOR_L1Results_6__6), .A1 (CALCULATOR_L1Results_7__6), .B0 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx56), .B1 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx0)) ;
    xor2 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix63 (.Y (
         CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx62), .A0 (CALCULATOR_L1Results_7__7)
         , .A1 (CALCULATOR_L1Results_6__7)) ;
    inv01 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix155 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx154), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx383)) ;
    inv01 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix57 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx56), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx561)) ;
    inv01 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix53 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx52), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx554)) ;
    inv01 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix49 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx48), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx547)) ;
    inv01 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix45 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx44), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx540)) ;
    inv01 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix41 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx40), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx534)) ;
    inv01 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix31 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx30), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx531)) ;
    inv01 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix25 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx24), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx537)) ;
    inv01 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix19 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx18), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx544)) ;
    inv01 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix13 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx12), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx551)) ;
    inv01 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix7 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx6), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx558)) ;
    inv01 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix1 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx0), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx565)) ;
    fake_gnd CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix216 (.Y (
             CALCULATOR_L1_3_L2_1_G2_MINI_ALU_WindowCellShiftedLeft_16)) ;
    aoi21 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix77 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_10), .A0 (
          CacheFilter_3__1__1), .A1 (CacheFilter_3__1__0), .B0 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_nx4)) ;
    nor02_2x CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix5 (.Y (
             CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_nx4), .A0 (
             CacheFilter_3__1__0), .A1 (CacheFilter_3__1__1)) ;
    aoi21 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix67 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_11), .A0 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_nx328), .A1 (
          CacheFilter_3__1__2), .B0 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_nx8)) ;
    nor03_2x CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix9 (.Y (
             CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_nx8), .A0 (
             CacheFilter_3__1__2), .A1 (CacheFilter_3__1__0), .A2 (
             CacheFilter_3__1__1)) ;
    xnor2 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix59 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_12), .A0 (
          CacheFilter_3__1__3), .A1 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_nx8)) ;
    xnor2 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix51 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_13), .A0 (
          CacheFilter_3__1__4), .A1 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_nx12)) ;
    nor04 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix13 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_nx12), .A0 (
          CacheFilter_3__1__3), .A1 (CacheFilter_3__1__2), .A2 (
          CacheFilter_3__1__0), .A3 (CacheFilter_3__1__1)) ;
    xnor2 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix43 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_14), .A0 (
          CacheFilter_3__1__5), .A1 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_nx16)) ;
    nor02ii CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix17 (.Y (
            CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_nx16), .A0 (
            CacheFilter_3__1__4), .A1 (
            CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_nx12)) ;
    xnor2 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix35 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_15), .A0 (
          CacheFilter_3__1__6), .A1 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_nx20)) ;
    nor02ii CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix21 (.Y (
            CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_nx20), .A0 (
            CacheFilter_3__1__5), .A1 (
            CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_nx16)) ;
    xnor2 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix27 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_16), .A0 (
          CacheFilter_3__1__7), .A1 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_nx24)) ;
    nor02ii CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix25 (.Y (
            CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_nx24), .A0 (
            CacheFilter_3__1__6), .A1 (
            CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_nx20)) ;
    inv01 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix329 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_nx328), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_nx4)) ;
    inv02 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix383 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_nx384), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_0)) ;
    dff CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_0 (.Q (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_0), .QB (
        \$dummy [843]), .D (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .CLK (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    nor02_2x CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix567 (.Y (
             CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566), .A0 (
             RST), .A1 (
             CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644)) ;
    dff CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_1 (.Q (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_1), .QB (
        \$dummy [844]), .D (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .CLK (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_2 (.Q (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_2), .QB (
        \$dummy [845]), .D (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .CLK (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_3 (.Q (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_3), .QB (
        \$dummy [846]), .D (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .CLK (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_4 (.Q (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_4), .QB (
        \$dummy [847]), .D (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .CLK (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_5 (.Q (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_5), .QB (
        \$dummy [848]), .D (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .CLK (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_6 (.Q (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_6), .QB (
        \$dummy [849]), .D (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .CLK (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_7 (.Q (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_7), .QB (
        \$dummy [850]), .D (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .CLK (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_8 (.Q (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_8), .QB (
        \$dummy [851]), .D (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .CLK (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_9 (.Q (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_9), .QB (
        \$dummy [852]), .D (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .CLK (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_10 (.Q (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_10), .QB (
        \$dummy [853]), .D (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .CLK (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_11 (.Q (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_11), .QB (
        \$dummy [854]), .D (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .CLK (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_12 (.Q (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_12), .QB (
        \$dummy [855]), .D (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .CLK (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_13 (.Q (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_13), .QB (
        \$dummy [856]), .D (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .CLK (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_14 (.Q (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_14), .QB (
        \$dummy [857]), .D (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .CLK (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_15 (.Q (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_15), .QB (
        \$dummy [858]), .D (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .CLK (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_16 (.Q (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_16), .QB (
        \$dummy [859]), .D (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .CLK (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    inv02 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix623 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix625 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix627 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix643 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644), .A (
          nx8019)) ;
    dff CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_0 (.Q (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_0), .QB (
        \$dummy [860]), .D (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .CLK (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    nor02_2x CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix567 (.Y (
             CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566), .A0 (
             RST), .A1 (
             CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644)) ;
    dff CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_1 (.Q (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_1), .QB (
        \$dummy [861]), .D (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .CLK (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_2 (.Q (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_2), .QB (
        \$dummy [862]), .D (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .CLK (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_3 (.Q (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_3), .QB (
        \$dummy [863]), .D (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .CLK (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_4 (.Q (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_4), .QB (
        \$dummy [864]), .D (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .CLK (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_5 (.Q (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_5), .QB (
        \$dummy [865]), .D (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .CLK (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_6 (.Q (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_6), .QB (
        \$dummy [866]), .D (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .CLK (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_7 (.Q (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_7), .QB (
        \$dummy [867]), .D (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .CLK (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_8 (.Q (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_8), .QB (
        \$dummy [868]), .D (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .CLK (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_9 (.Q (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_9), .QB (
        \$dummy [869]), .D (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .CLK (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_10 (.Q (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_10), .QB (
        \$dummy [870]), .D (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .CLK (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_11 (.Q (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_11), .QB (
        \$dummy [871]), .D (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .CLK (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_12 (.Q (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_12), .QB (
        \$dummy [872]), .D (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .CLK (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_13 (.Q (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_13), .QB (
        \$dummy [873]), .D (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .CLK (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_14 (.Q (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_14), .QB (
        \$dummy [874]), .D (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .CLK (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_15 (.Q (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_15), .QB (
        \$dummy [875]), .D (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .CLK (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_16 (.Q (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_16), .QB (
        \$dummy [876]), .D (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .CLK (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    inv02 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix623 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix625 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix627 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix643 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644), .A (
          nx8025)) ;
    dff CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_0 (.Q (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_0), .QB (\$dummy [877]), .D (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .CLK (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    nor02_2x CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix567 (.Y (
             CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566), .A0 (
             RST), .A1 (
             CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    dff CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_1 (.Q (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_1), .QB (\$dummy [878]), .D (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .CLK (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_2 (.Q (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_2), .QB (\$dummy [879]), .D (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .CLK (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_3 (.Q (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_3), .QB (\$dummy [880]), .D (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .CLK (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_4 (.Q (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_4), .QB (\$dummy [881]), .D (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .CLK (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_5 (.Q (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_5), .QB (\$dummy [882]), .D (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .CLK (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_6 (.Q (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_6), .QB (\$dummy [883]), .D (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .CLK (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_7 (.Q (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_7), .QB (\$dummy [884]), .D (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .CLK (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_8 (.Q (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_8), .QB (\$dummy [885]), .D (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .CLK (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_9 (.Q (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_9), .QB (\$dummy [886]), .D (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .CLK (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_10 (.Q (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_10), .QB (\$dummy [887]), .D (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .CLK (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_11 (.Q (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_11), .QB (\$dummy [888]), .D (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .CLK (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_12 (.Q (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_12), .QB (\$dummy [889]), .D (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .CLK (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_13 (.Q (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_13), .QB (\$dummy [890]), .D (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .CLK (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_14 (.Q (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_14), .QB (\$dummy [891]), .D (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .CLK (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_15 (.Q (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_15), .QB (\$dummy [892]), .D (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .CLK (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_16 (.Q (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_16), .QB (\$dummy [893]), .D (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .CLK (
        CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    inv02 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix623 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix625 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix627 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix643 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642)) ;
    xor2 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix83 (.Y (CALCULATOR_L2Results_4__0), 
         .A0 (CALCULATOR_L1Results_9__0), .A1 (CALCULATOR_L1Results_8__0)) ;
    xnor2 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix380 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx379), .A0 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx381), .A1 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx383)) ;
    nand02 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix382 (.Y (
           CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx381), .A0 (
           CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothOperand_0), .A1 (nx8045)) ;
    xnor2 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix384 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx383), .A0 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothOperand_1), .A1 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_1)) ;
    inv01 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix388 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx387), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_2)) ;
    xnor2 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix390 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx389), .A0 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx391), .A1 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx395)) ;
    aoi32 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix392 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx391), .A0 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothOperand_0), .A1 (nx8045), .A2 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx154), .B0 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_1), .B1 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothOperand_1)) ;
    xnor2 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix396 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx395), .A0 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothOperand_2), .A1 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_2)) ;
    inv01 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix400 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx399), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_3)) ;
    xnor2 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix402 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx401), .A0 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx403), .A1 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx405)) ;
    xnor2 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix406 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx405), .A0 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothOperand_3), .A1 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_3)) ;
    inv01 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix410 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx409), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_4)) ;
    xnor2 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix412 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx411), .A0 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx413), .A1 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx415)) ;
    xnor2 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix416 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx415), .A0 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothOperand_4), .A1 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_4)) ;
    inv01 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix420 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx419), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_5)) ;
    xnor2 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix422 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx421), .A0 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx423), .A1 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx425)) ;
    xnor2 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix426 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx425), .A0 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothOperand_5), .A1 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_5)) ;
    inv01 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix430 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx429), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_6)) ;
    xnor2 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix432 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx431), .A0 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx433), .A1 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx435)) ;
    xnor2 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix436 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx435), .A0 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothOperand_6), .A1 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_6)) ;
    inv01 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix440 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx439), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_7)) ;
    xnor2 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix442 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx441), .A0 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx443), .A1 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx445)) ;
    xnor2 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix446 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx445), .A0 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothOperand_7), .A1 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_7)) ;
    inv01 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix450 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx449), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_8)) ;
    xnor2 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix452 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx451), .A0 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx453), .A1 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx455)) ;
    xnor2 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix456 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx455), .A0 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothOperand_8), .A1 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_8)) ;
    xor2 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix317 (.Y (
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx316), .A0 (
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx461), .A1 (
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx463)) ;
    xnor2 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix464 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx463), .A0 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothOperand_9), .A1 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_9)) ;
    xor2 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix337 (.Y (
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx336), .A0 (
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx467), .A1 (
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx471)) ;
    inv01 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix470 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx469), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_9)) ;
    xnor2 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix472 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx471), .A0 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothOperand_10), .A1 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_10)) ;
    xor2 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix357 (.Y (
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx356), .A0 (
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx475), .A1 (
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx479)) ;
    inv01 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix478 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx477), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_10)) ;
    xnor2 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix480 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx479), .A0 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothOperand_11), .A1 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_11)) ;
    xor2 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix377 (.Y (
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx376), .A0 (
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx483), .A1 (
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx487)) ;
    inv01 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix486 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx485), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_11)) ;
    xnor2 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix488 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx487), .A0 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothOperand_12), .A1 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_12)) ;
    xor2 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix397 (.Y (
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx396), .A0 (
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx491), .A1 (
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx495)) ;
    inv01 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix494 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx493), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_12)) ;
    xnor2 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix496 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx495), .A0 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothOperand_13), .A1 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_13)) ;
    xor2 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix417 (.Y (
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx416), .A0 (
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx499), .A1 (
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx503)) ;
    inv01 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix502 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx501), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_13)) ;
    xnor2 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix504 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx503), .A0 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothOperand_14), .A1 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_14)) ;
    xor2 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix437 (.Y (
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx436), .A0 (
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx507), .A1 (
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx511)) ;
    inv01 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix510 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx509), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_14)) ;
    xnor2 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix512 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx511), .A0 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothOperand_15), .A1 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_15)) ;
    xnor2 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix457 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx456), .A0 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx515), .A1 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx454)) ;
    inv01 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix518 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx517), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_15)) ;
    xor2 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix455 (.Y (
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx454), .A0 (
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothOperand_16), .A1 (
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_16)) ;
    mux21_ni CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix91 (.Y (
             CALCULATOR_L1FirstOperands_8__0), .A0 (
             CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_1), .A1 (
             CacheWindow_3__2__0), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix99 (.Y (
             CALCULATOR_L1FirstOperands_8__1), .A0 (
             CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_2), .A1 (
             CacheWindow_3__2__1), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix107 (.Y (
             CALCULATOR_L1FirstOperands_8__2), .A0 (
             CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_3), .A1 (
             CacheWindow_3__2__2), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix115 (.Y (
             CALCULATOR_L1FirstOperands_8__3), .A0 (
             CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_4), .A1 (
             CacheWindow_3__2__3), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix123 (.Y (
             CALCULATOR_L1FirstOperands_8__4), .A0 (
             CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_5), .A1 (
             CacheWindow_3__2__4), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix131 (.Y (
             CALCULATOR_L1FirstOperands_8__5), .A0 (
             CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_6), .A1 (
             CacheWindow_3__2__5), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix139 (.Y (
             CALCULATOR_L1FirstOperands_8__6), .A0 (
             CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_7), .A1 (
             CacheWindow_3__2__6), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix147 (.Y (
             CALCULATOR_L1FirstOperands_8__7), .A0 (
             CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_8), .A1 (
             CacheWindow_3__2__7), .S0 (Instr)) ;
    xor2 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix77 (.Y (CALCULATOR_L2Results_4__1), 
         .A0 (CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx529), .A1 (
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx531)) ;
    nand02 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix530 (.Y (
           CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx529), .A0 (
           CALCULATOR_L1Results_9__0), .A1 (CALCULATOR_L1Results_8__0)) ;
    xnor2 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix532 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx531), .A0 (
          CALCULATOR_L1Results_9__1), .A1 (CALCULATOR_L1Results_8__1)) ;
    xor2 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix75 (.Y (CALCULATOR_L2Results_4__2), 
         .A0 (CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx534), .A1 (
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx537)) ;
    aoi32 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix535 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx534), .A0 (
          CALCULATOR_L1Results_9__0), .A1 (CALCULATOR_L1Results_8__0), .A2 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx30), .B0 (CALCULATOR_L1Results_8__1
          ), .B1 (CALCULATOR_L1Results_9__1)) ;
    xnor2 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix538 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx537), .A0 (
          CALCULATOR_L1Results_9__2), .A1 (CALCULATOR_L1Results_8__2)) ;
    xor2 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix73 (.Y (CALCULATOR_L2Results_4__3), 
         .A0 (CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx540), .A1 (
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx544)) ;
    aoi22 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix541 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx540), .A0 (
          CALCULATOR_L1Results_8__2), .A1 (CALCULATOR_L1Results_9__2), .B0 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx40), .B1 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx24)) ;
    xnor2 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix545 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx544), .A0 (
          CALCULATOR_L1Results_9__3), .A1 (CALCULATOR_L1Results_8__3)) ;
    xor2 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix71 (.Y (CALCULATOR_L2Results_4__4), 
         .A0 (CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx547), .A1 (
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx551)) ;
    aoi22 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix548 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx547), .A0 (
          CALCULATOR_L1Results_8__3), .A1 (CALCULATOR_L1Results_9__3), .B0 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx44), .B1 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx18)) ;
    xnor2 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix552 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx551), .A0 (
          CALCULATOR_L1Results_9__4), .A1 (CALCULATOR_L1Results_8__4)) ;
    xor2 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix69 (.Y (CALCULATOR_L2Results_4__5), 
         .A0 (CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx554), .A1 (
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx558)) ;
    aoi22 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix555 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx554), .A0 (
          CALCULATOR_L1Results_8__4), .A1 (CALCULATOR_L1Results_9__4), .B0 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx48), .B1 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx12)) ;
    xnor2 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix559 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx558), .A0 (
          CALCULATOR_L1Results_9__5), .A1 (CALCULATOR_L1Results_8__5)) ;
    xor2 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix67 (.Y (CALCULATOR_L2Results_4__6), 
         .A0 (CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx561), .A1 (
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx565)) ;
    aoi22 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix562 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx561), .A0 (
          CALCULATOR_L1Results_8__5), .A1 (CALCULATOR_L1Results_9__5), .B0 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx52), .B1 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx6)) ;
    xnor2 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix566 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx565), .A0 (
          CALCULATOR_L1Results_9__6), .A1 (CALCULATOR_L1Results_8__6)) ;
    xnor2 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix65 (.Y (CALCULATOR_L2Results_4__7)
          , .A0 (CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx568), .A1 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx62)) ;
    aoi22 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix569 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx568), .A0 (
          CALCULATOR_L1Results_8__6), .A1 (CALCULATOR_L1Results_9__6), .B0 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx56), .B1 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx0)) ;
    xor2 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix63 (.Y (
         CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx62), .A0 (CALCULATOR_L1Results_9__7)
         , .A1 (CALCULATOR_L1Results_8__7)) ;
    inv01 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix155 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx154), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx383)) ;
    inv01 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix57 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx56), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx561)) ;
    inv01 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix53 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx52), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx554)) ;
    inv01 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix49 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx48), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx547)) ;
    inv01 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix45 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx44), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx540)) ;
    inv01 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix41 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx40), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx534)) ;
    inv01 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix31 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx30), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx531)) ;
    inv01 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix25 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx24), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx537)) ;
    inv01 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix19 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx18), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx544)) ;
    inv01 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix13 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx12), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx551)) ;
    inv01 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix7 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx6), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx558)) ;
    inv01 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix1 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx0), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx565)) ;
    fake_gnd CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix216 (.Y (
             CALCULATOR_L1_3_L2_2_G2_MINI_ALU_WindowCellShiftedLeft_16)) ;
    aoi21 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix77 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_10), .A0 (
          CacheFilter_3__2__1), .A1 (CacheFilter_3__2__0), .B0 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_nx4)) ;
    nor02_2x CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix5 (.Y (
             CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_nx4), .A0 (
             CacheFilter_3__2__0), .A1 (CacheFilter_3__2__1)) ;
    aoi21 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix67 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_11), .A0 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_nx328), .A1 (
          CacheFilter_3__2__2), .B0 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_nx8)) ;
    nor03_2x CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix9 (.Y (
             CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_nx8), .A0 (
             CacheFilter_3__2__2), .A1 (CacheFilter_3__2__0), .A2 (
             CacheFilter_3__2__1)) ;
    xnor2 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix59 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_12), .A0 (
          CacheFilter_3__2__3), .A1 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_nx8)) ;
    xnor2 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix51 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_13), .A0 (
          CacheFilter_3__2__4), .A1 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_nx12)) ;
    nor04 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix13 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_nx12), .A0 (
          CacheFilter_3__2__3), .A1 (CacheFilter_3__2__2), .A2 (
          CacheFilter_3__2__0), .A3 (CacheFilter_3__2__1)) ;
    xnor2 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix43 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_14), .A0 (
          CacheFilter_3__2__5), .A1 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_nx16)) ;
    nor02ii CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix17 (.Y (
            CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_nx16), .A0 (
            CacheFilter_3__2__4), .A1 (
            CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_nx12)) ;
    xnor2 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix35 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_15), .A0 (
          CacheFilter_3__2__6), .A1 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_nx20)) ;
    nor02ii CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix21 (.Y (
            CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_nx20), .A0 (
            CacheFilter_3__2__5), .A1 (
            CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_nx16)) ;
    xnor2 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix27 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_16), .A0 (
          CacheFilter_3__2__7), .A1 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_nx24)) ;
    nor02ii CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix25 (.Y (
            CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_nx24), .A0 (
            CacheFilter_3__2__6), .A1 (
            CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_nx20)) ;
    inv01 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix329 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_nx328), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_nx4)) ;
    inv02 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix383 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_nx384), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_0)) ;
    dff CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_0 (.Q (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_0), .QB (
        \$dummy [894]), .D (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .CLK (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    nor02_2x CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix567 (.Y (
             CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566), .A0 (
             RST), .A1 (
             CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644)) ;
    dff CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_1 (.Q (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_1), .QB (
        \$dummy [895]), .D (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .CLK (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_2 (.Q (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_2), .QB (
        \$dummy [896]), .D (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .CLK (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_3 (.Q (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_3), .QB (
        \$dummy [897]), .D (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .CLK (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_4 (.Q (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_4), .QB (
        \$dummy [898]), .D (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .CLK (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_5 (.Q (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_5), .QB (
        \$dummy [899]), .D (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .CLK (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_6 (.Q (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_6), .QB (
        \$dummy [900]), .D (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .CLK (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_7 (.Q (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_7), .QB (
        \$dummy [901]), .D (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .CLK (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_8 (.Q (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_8), .QB (
        \$dummy [902]), .D (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .CLK (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_9 (.Q (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_9), .QB (
        \$dummy [903]), .D (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .CLK (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_10 (.Q (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_10), .QB (
        \$dummy [904]), .D (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .CLK (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_11 (.Q (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_11), .QB (
        \$dummy [905]), .D (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .CLK (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_12 (.Q (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_12), .QB (
        \$dummy [906]), .D (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .CLK (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_13 (.Q (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_13), .QB (
        \$dummy [907]), .D (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .CLK (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_14 (.Q (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_14), .QB (
        \$dummy [908]), .D (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .CLK (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_15 (.Q (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_15), .QB (
        \$dummy [909]), .D (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .CLK (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_16 (.Q (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_16), .QB (
        \$dummy [910]), .D (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .CLK (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    inv02 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix623 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix625 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix627 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix643 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644), .A (
          nx8059)) ;
    dff CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_0 (.Q (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_0), .QB (
        \$dummy [911]), .D (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .CLK (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    nor02_2x CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix567 (.Y (
             CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566), .A0 (
             RST), .A1 (
             CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644)) ;
    dff CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_1 (.Q (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_1), .QB (
        \$dummy [912]), .D (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .CLK (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_2 (.Q (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_2), .QB (
        \$dummy [913]), .D (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .CLK (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_3 (.Q (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_3), .QB (
        \$dummy [914]), .D (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .CLK (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_4 (.Q (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_4), .QB (
        \$dummy [915]), .D (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .CLK (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_5 (.Q (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_5), .QB (
        \$dummy [916]), .D (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .CLK (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_6 (.Q (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_6), .QB (
        \$dummy [917]), .D (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .CLK (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_7 (.Q (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_7), .QB (
        \$dummy [918]), .D (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .CLK (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_8 (.Q (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_8), .QB (
        \$dummy [919]), .D (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .CLK (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_9 (.Q (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_9), .QB (
        \$dummy [920]), .D (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .CLK (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_10 (.Q (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_10), .QB (
        \$dummy [921]), .D (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .CLK (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_11 (.Q (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_11), .QB (
        \$dummy [922]), .D (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .CLK (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_12 (.Q (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_12), .QB (
        \$dummy [923]), .D (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .CLK (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_13 (.Q (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_13), .QB (
        \$dummy [924]), .D (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .CLK (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_14 (.Q (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_14), .QB (
        \$dummy [925]), .D (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .CLK (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_15 (.Q (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_15), .QB (
        \$dummy [926]), .D (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .CLK (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_16 (.Q (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_16), .QB (
        \$dummy [927]), .D (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .CLK (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    inv02 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix623 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix625 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix627 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix643 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644), .A (
          nx8065)) ;
    dff CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_0 (.Q (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_0), .QB (\$dummy [928]), .D (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .CLK (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    nor02_2x CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix567 (.Y (
             CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566), .A0 (
             RST), .A1 (
             CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    dff CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_1 (.Q (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_1), .QB (\$dummy [929]), .D (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .CLK (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_2 (.Q (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_2), .QB (\$dummy [930]), .D (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .CLK (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_3 (.Q (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_3), .QB (\$dummy [931]), .D (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .CLK (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_4 (.Q (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_4), .QB (\$dummy [932]), .D (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .CLK (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_5 (.Q (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_5), .QB (\$dummy [933]), .D (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .CLK (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_6 (.Q (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_6), .QB (\$dummy [934]), .D (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .CLK (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_7 (.Q (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_7), .QB (\$dummy [935]), .D (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .CLK (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_8 (.Q (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_8), .QB (\$dummy [936]), .D (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .CLK (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_9 (.Q (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_9), .QB (\$dummy [937]), .D (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .CLK (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_10 (.Q (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_10), .QB (\$dummy [938]), .D (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .CLK (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_11 (.Q (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_11), .QB (\$dummy [939]), .D (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .CLK (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_12 (.Q (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_12), .QB (\$dummy [940]), .D (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .CLK (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_13 (.Q (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_13), .QB (\$dummy [941]), .D (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .CLK (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_14 (.Q (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_14), .QB (\$dummy [942]), .D (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .CLK (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_15 (.Q (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_15), .QB (\$dummy [943]), .D (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .CLK (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_16 (.Q (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_16), .QB (\$dummy [944]), .D (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .CLK (
        CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    inv02 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix623 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix625 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix627 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix643 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642)) ;
    xor2 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix83 (.Y (CALCULATOR_L2Results_5__0), 
         .A0 (CALCULATOR_L1Results_11__0), .A1 (CALCULATOR_L1Results_10__0)) ;
    xnor2 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix380 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx379), .A0 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx381), .A1 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx383)) ;
    nand02 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix382 (.Y (
           CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx381), .A0 (
           CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothOperand_0), .A1 (nx8085)) ;
    xnor2 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix384 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx383), .A0 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothOperand_1), .A1 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_1)) ;
    inv01 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix388 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx387), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_2)) ;
    xnor2 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix390 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx389), .A0 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx391), .A1 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx395)) ;
    aoi32 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix392 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx391), .A0 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothOperand_0), .A1 (nx8085), .A2 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx154), .B0 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_1), .B1 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothOperand_1)) ;
    xnor2 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix396 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx395), .A0 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothOperand_2), .A1 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_2)) ;
    inv01 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix400 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx399), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_3)) ;
    xnor2 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix402 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx401), .A0 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx403), .A1 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx405)) ;
    xnor2 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix406 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx405), .A0 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothOperand_3), .A1 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_3)) ;
    inv01 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix410 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx409), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_4)) ;
    xnor2 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix412 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx411), .A0 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx413), .A1 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx415)) ;
    xnor2 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix416 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx415), .A0 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothOperand_4), .A1 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_4)) ;
    inv01 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix420 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx419), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_5)) ;
    xnor2 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix422 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx421), .A0 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx423), .A1 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx425)) ;
    xnor2 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix426 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx425), .A0 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothOperand_5), .A1 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_5)) ;
    inv01 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix430 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx429), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_6)) ;
    xnor2 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix432 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx431), .A0 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx433), .A1 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx435)) ;
    xnor2 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix436 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx435), .A0 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothOperand_6), .A1 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_6)) ;
    inv01 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix440 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx439), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_7)) ;
    xnor2 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix442 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx441), .A0 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx443), .A1 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx445)) ;
    xnor2 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix446 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx445), .A0 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothOperand_7), .A1 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_7)) ;
    inv01 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix450 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx449), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_8)) ;
    xnor2 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix452 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx451), .A0 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx453), .A1 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx455)) ;
    xnor2 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix456 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx455), .A0 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothOperand_8), .A1 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_8)) ;
    xor2 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix317 (.Y (
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx316), .A0 (
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx461), .A1 (
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx463)) ;
    xnor2 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix464 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx463), .A0 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothOperand_9), .A1 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_9)) ;
    xor2 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix337 (.Y (
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx336), .A0 (
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx467), .A1 (
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx471)) ;
    inv01 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix470 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx469), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_9)) ;
    xnor2 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix472 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx471), .A0 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothOperand_10), .A1 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_10)) ;
    xor2 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix357 (.Y (
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx356), .A0 (
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx475), .A1 (
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx479)) ;
    inv01 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix478 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx477), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_10)) ;
    xnor2 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix480 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx479), .A0 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothOperand_11), .A1 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_11)) ;
    xor2 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix377 (.Y (
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx376), .A0 (
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx483), .A1 (
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx487)) ;
    inv01 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix486 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx485), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_11)) ;
    xnor2 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix488 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx487), .A0 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothOperand_12), .A1 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_12)) ;
    xor2 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix397 (.Y (
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx396), .A0 (
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx491), .A1 (
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx495)) ;
    inv01 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix494 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx493), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_12)) ;
    xnor2 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix496 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx495), .A0 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothOperand_13), .A1 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_13)) ;
    xor2 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix417 (.Y (
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx416), .A0 (
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx499), .A1 (
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx503)) ;
    inv01 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix502 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx501), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_13)) ;
    xnor2 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix504 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx503), .A0 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothOperand_14), .A1 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_14)) ;
    xor2 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix437 (.Y (
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx436), .A0 (
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx507), .A1 (
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx511)) ;
    inv01 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix510 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx509), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_14)) ;
    xnor2 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix512 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx511), .A0 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothOperand_15), .A1 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_15)) ;
    xnor2 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix457 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx456), .A0 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx515), .A1 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx454)) ;
    inv01 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix518 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx517), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_15)) ;
    xor2 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix455 (.Y (
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx454), .A0 (
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothOperand_16), .A1 (
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_16)) ;
    mux21_ni CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix91 (.Y (
             CALCULATOR_L1FirstOperands_10__0), .A0 (
             CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_1), .A1 (
             CacheWindow_3__3__0), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix99 (.Y (
             CALCULATOR_L1FirstOperands_10__1), .A0 (
             CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_2), .A1 (
             CacheWindow_3__3__1), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix107 (.Y (
             CALCULATOR_L1FirstOperands_10__2), .A0 (
             CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_3), .A1 (
             CacheWindow_3__3__2), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix115 (.Y (
             CALCULATOR_L1FirstOperands_10__3), .A0 (
             CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_4), .A1 (
             CacheWindow_3__3__3), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix123 (.Y (
             CALCULATOR_L1FirstOperands_10__4), .A0 (
             CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_5), .A1 (
             CacheWindow_3__3__4), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix131 (.Y (
             CALCULATOR_L1FirstOperands_10__5), .A0 (
             CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_6), .A1 (
             CacheWindow_3__3__5), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix139 (.Y (
             CALCULATOR_L1FirstOperands_10__6), .A0 (
             CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_7), .A1 (
             CacheWindow_3__3__6), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix147 (.Y (
             CALCULATOR_L1FirstOperands_10__7), .A0 (
             CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_8), .A1 (
             CacheWindow_3__3__7), .S0 (Instr)) ;
    xor2 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix77 (.Y (CALCULATOR_L2Results_5__1), 
         .A0 (CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx529), .A1 (
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx531)) ;
    nand02 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix530 (.Y (
           CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx529), .A0 (
           CALCULATOR_L1Results_11__0), .A1 (CALCULATOR_L1Results_10__0)) ;
    xnor2 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix532 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx531), .A0 (
          CALCULATOR_L1Results_11__1), .A1 (CALCULATOR_L1Results_10__1)) ;
    xor2 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix75 (.Y (CALCULATOR_L2Results_5__2), 
         .A0 (CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx534), .A1 (
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx537)) ;
    aoi32 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix535 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx534), .A0 (
          CALCULATOR_L1Results_11__0), .A1 (CALCULATOR_L1Results_10__0), .A2 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx30), .B0 (
          CALCULATOR_L1Results_10__1), .B1 (CALCULATOR_L1Results_11__1)) ;
    xnor2 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix538 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx537), .A0 (
          CALCULATOR_L1Results_11__2), .A1 (CALCULATOR_L1Results_10__2)) ;
    xor2 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix73 (.Y (CALCULATOR_L2Results_5__3), 
         .A0 (CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx540), .A1 (
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx544)) ;
    aoi22 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix541 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx540), .A0 (
          CALCULATOR_L1Results_10__2), .A1 (CALCULATOR_L1Results_11__2), .B0 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx40), .B1 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx24)) ;
    xnor2 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix545 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx544), .A0 (
          CALCULATOR_L1Results_11__3), .A1 (CALCULATOR_L1Results_10__3)) ;
    xor2 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix71 (.Y (CALCULATOR_L2Results_5__4), 
         .A0 (CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx547), .A1 (
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx551)) ;
    aoi22 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix548 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx547), .A0 (
          CALCULATOR_L1Results_10__3), .A1 (CALCULATOR_L1Results_11__3), .B0 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx44), .B1 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx18)) ;
    xnor2 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix552 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx551), .A0 (
          CALCULATOR_L1Results_11__4), .A1 (CALCULATOR_L1Results_10__4)) ;
    xor2 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix69 (.Y (CALCULATOR_L2Results_5__5), 
         .A0 (CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx554), .A1 (
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx558)) ;
    aoi22 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix555 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx554), .A0 (
          CALCULATOR_L1Results_10__4), .A1 (CALCULATOR_L1Results_11__4), .B0 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx48), .B1 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx12)) ;
    xnor2 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix559 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx558), .A0 (
          CALCULATOR_L1Results_11__5), .A1 (CALCULATOR_L1Results_10__5)) ;
    xor2 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix67 (.Y (CALCULATOR_L2Results_5__6), 
         .A0 (CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx561), .A1 (
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx565)) ;
    aoi22 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix562 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx561), .A0 (
          CALCULATOR_L1Results_10__5), .A1 (CALCULATOR_L1Results_11__5), .B0 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx52), .B1 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx6)) ;
    xnor2 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix566 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx565), .A0 (
          CALCULATOR_L1Results_11__6), .A1 (CALCULATOR_L1Results_10__6)) ;
    xnor2 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix65 (.Y (CALCULATOR_L2Results_5__7)
          , .A0 (CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx568), .A1 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx62)) ;
    aoi22 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix569 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx568), .A0 (
          CALCULATOR_L1Results_10__6), .A1 (CALCULATOR_L1Results_11__6), .B0 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx56), .B1 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx0)) ;
    xor2 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix63 (.Y (
         CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx62), .A0 (CALCULATOR_L1Results_11__7
         ), .A1 (CALCULATOR_L1Results_10__7)) ;
    inv01 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix155 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx154), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx383)) ;
    inv01 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix57 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx56), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx561)) ;
    inv01 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix53 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx52), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx554)) ;
    inv01 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix49 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx48), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx547)) ;
    inv01 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix45 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx44), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx540)) ;
    inv01 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix41 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx40), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx534)) ;
    inv01 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix31 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx30), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx531)) ;
    inv01 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix25 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx24), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx537)) ;
    inv01 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix19 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx18), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx544)) ;
    inv01 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix13 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx12), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx551)) ;
    inv01 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix7 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx6), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx558)) ;
    inv01 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix1 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx0), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx565)) ;
    fake_gnd CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix216 (.Y (
             CALCULATOR_L1_3_L2_3_G2_MINI_ALU_WindowCellShiftedLeft_16)) ;
    aoi21 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix77 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_10), .A0 (
          CacheFilter_3__3__1), .A1 (CacheFilter_3__3__0), .B0 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx4)) ;
    nor02_2x CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix5 (.Y (
             CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx4), .A0 (
             CacheFilter_3__3__0), .A1 (CacheFilter_3__3__1)) ;
    aoi21 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix67 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_11), .A0 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx328), .A1 (
          CacheFilter_3__3__2), .B0 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx8)) ;
    nor03_2x CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix9 (.Y (
             CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx8), .A0 (
             CacheFilter_3__3__2), .A1 (CacheFilter_3__3__0), .A2 (
             CacheFilter_3__3__1)) ;
    xnor2 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix59 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_12), .A0 (
          CacheFilter_3__3__3), .A1 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx8)) ;
    xnor2 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix51 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_13), .A0 (
          CacheFilter_3__3__4), .A1 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx12)) ;
    nor04 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix13 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx12), .A0 (
          CacheFilter_3__3__3), .A1 (CacheFilter_3__3__2), .A2 (
          CacheFilter_3__3__0), .A3 (CacheFilter_3__3__1)) ;
    xnor2 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix43 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_14), .A0 (
          CacheFilter_3__3__5), .A1 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx16)) ;
    nor02ii CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix17 (.Y (
            CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx16), .A0 (
            CacheFilter_3__3__4), .A1 (
            CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx12)) ;
    xnor2 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix35 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_15), .A0 (
          CacheFilter_3__3__6), .A1 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx20)) ;
    nor02ii CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix21 (.Y (
            CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx20), .A0 (
            CacheFilter_3__3__5), .A1 (
            CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx16)) ;
    xnor2 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix27 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_16), .A0 (
          CacheFilter_3__3__7), .A1 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx24)) ;
    nor02ii CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix25 (.Y (
            CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx24), .A0 (
            CacheFilter_3__3__6), .A1 (
            CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx20)) ;
    inv01 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix329 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx328), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx4)) ;
    inv02 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix383 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx384), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_0)) ;
    dff CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_0 (.Q (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_0), .QB (
        \$dummy [945]), .D (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .CLK (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    nor02_2x CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix567 (.Y (
             CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566), .A0 (
             RST), .A1 (
             CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644)) ;
    dff CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_1 (.Q (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_1), .QB (
        \$dummy [946]), .D (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .CLK (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_2 (.Q (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_2), .QB (
        \$dummy [947]), .D (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .CLK (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_3 (.Q (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_3), .QB (
        \$dummy [948]), .D (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .CLK (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_4 (.Q (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_4), .QB (
        \$dummy [949]), .D (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .CLK (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_5 (.Q (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_5), .QB (
        \$dummy [950]), .D (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .CLK (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_6 (.Q (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_6), .QB (
        \$dummy [951]), .D (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .CLK (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_7 (.Q (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_7), .QB (
        \$dummy [952]), .D (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .CLK (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_8 (.Q (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_8), .QB (
        \$dummy [953]), .D (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .CLK (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_9 (.Q (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_9), .QB (
        \$dummy [954]), .D (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .CLK (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_10 (.Q (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_10), .QB (
        \$dummy [955]), .D (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .CLK (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_11 (.Q (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_11), .QB (
        \$dummy [956]), .D (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .CLK (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_12 (.Q (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_12), .QB (
        \$dummy [957]), .D (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .CLK (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_13 (.Q (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_13), .QB (
        \$dummy [958]), .D (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .CLK (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_14 (.Q (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_14), .QB (
        \$dummy [959]), .D (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .CLK (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_15 (.Q (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_15), .QB (
        \$dummy [960]), .D (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .CLK (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_16 (.Q (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_16), .QB (
        \$dummy [961]), .D (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .CLK (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    inv02 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix623 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix625 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix627 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix643 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644), .A (
          nx8099)) ;
    dff CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_0 (.Q (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_0), .QB (
        \$dummy [962]), .D (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .CLK (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    nor02_2x CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix567 (.Y (
             CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566), .A0 (
             RST), .A1 (
             CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644)) ;
    dff CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_1 (.Q (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_1), .QB (
        \$dummy [963]), .D (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .CLK (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_2 (.Q (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_2), .QB (
        \$dummy [964]), .D (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .CLK (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_3 (.Q (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_3), .QB (
        \$dummy [965]), .D (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .CLK (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_4 (.Q (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_4), .QB (
        \$dummy [966]), .D (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .CLK (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_5 (.Q (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_5), .QB (
        \$dummy [967]), .D (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .CLK (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_6 (.Q (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_6), .QB (
        \$dummy [968]), .D (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .CLK (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_7 (.Q (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_7), .QB (
        \$dummy [969]), .D (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .CLK (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_8 (.Q (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_8), .QB (
        \$dummy [970]), .D (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .CLK (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_9 (.Q (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_9), .QB (
        \$dummy [971]), .D (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .CLK (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_10 (.Q (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_10), .QB (
        \$dummy [972]), .D (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .CLK (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_11 (.Q (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_11), .QB (
        \$dummy [973]), .D (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .CLK (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_12 (.Q (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_12), .QB (
        \$dummy [974]), .D (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .CLK (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_13 (.Q (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_13), .QB (
        \$dummy [975]), .D (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .CLK (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_14 (.Q (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_14), .QB (
        \$dummy [976]), .D (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .CLK (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_15 (.Q (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_15), .QB (
        \$dummy [977]), .D (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .CLK (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_16 (.Q (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_16), .QB (
        \$dummy [978]), .D (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .CLK (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    inv02 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix623 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix625 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix627 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix643 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644), .A (
          nx8105)) ;
    dff CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_0 (.Q (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_0), .QB (\$dummy [979]), .D (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .CLK (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    nor02_2x CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix567 (.Y (
             CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566), .A0 (
             RST), .A1 (
             CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    dff CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_1 (.Q (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_1), .QB (\$dummy [980]), .D (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .CLK (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_2 (.Q (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_2), .QB (\$dummy [981]), .D (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .CLK (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_3 (.Q (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_3), .QB (\$dummy [982]), .D (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .CLK (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_4 (.Q (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_4), .QB (\$dummy [983]), .D (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .CLK (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_5 (.Q (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_5), .QB (\$dummy [984]), .D (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .CLK (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_6 (.Q (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_6), .QB (\$dummy [985]), .D (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .CLK (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_7 (.Q (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_7), .QB (\$dummy [986]), .D (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .CLK (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_8 (.Q (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_8), .QB (\$dummy [987]), .D (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .CLK (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_9 (.Q (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_9), .QB (\$dummy [988]), .D (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .CLK (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_10 (.Q (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_10), .QB (\$dummy [989]), .D (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .CLK (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_11 (.Q (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_11), .QB (\$dummy [990]), .D (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .CLK (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_12 (.Q (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_12), .QB (\$dummy [991]), .D (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .CLK (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_13 (.Q (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_13), .QB (\$dummy [992]), .D (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .CLK (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_14 (.Q (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_14), .QB (\$dummy [993]), .D (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .CLK (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_15 (.Q (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_15), .QB (\$dummy [994]), .D (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .CLK (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_16 (.Q (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_16), .QB (\$dummy [995]), .D (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .CLK (
        CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    inv02 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix623 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix625 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix627 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix643 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642)) ;
    xor2 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix83 (.Y (CALCULATOR_L3Results_0__0), 
         .A0 (CALCULATOR_L2Results_1__0), .A1 (CALCULATOR_L2Results_0__0)) ;
    xnor2 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix380 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx379), .A0 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx381), .A1 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx383)) ;
    nand02 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix382 (.Y (
           CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx381), .A0 (
           CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothOperand_0), .A1 (nx8125)) ;
    xnor2 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix384 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx383), .A0 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothOperand_1), .A1 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_1)) ;
    inv01 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix388 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx387), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_2)) ;
    xnor2 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix390 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx389), .A0 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx391), .A1 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx395)) ;
    aoi32 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix392 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx391), .A0 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothOperand_0), .A1 (nx8125), .A2 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx154), .B0 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_1), .B1 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothOperand_1)) ;
    xnor2 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix396 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx395), .A0 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothOperand_2), .A1 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_2)) ;
    inv01 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix400 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx399), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_3)) ;
    xnor2 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix402 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx401), .A0 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx403), .A1 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx405)) ;
    xnor2 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix406 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx405), .A0 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothOperand_3), .A1 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_3)) ;
    inv01 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix410 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx409), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_4)) ;
    xnor2 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix412 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx411), .A0 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx413), .A1 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx415)) ;
    xnor2 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix416 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx415), .A0 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothOperand_4), .A1 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_4)) ;
    inv01 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix420 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx419), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_5)) ;
    xnor2 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix422 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx421), .A0 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx423), .A1 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx425)) ;
    xnor2 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix426 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx425), .A0 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothOperand_5), .A1 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_5)) ;
    inv01 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix430 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx429), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_6)) ;
    xnor2 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix432 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx431), .A0 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx433), .A1 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx435)) ;
    xnor2 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix436 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx435), .A0 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothOperand_6), .A1 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_6)) ;
    inv01 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix440 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx439), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_7)) ;
    xnor2 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix442 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx441), .A0 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx443), .A1 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx445)) ;
    xnor2 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix446 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx445), .A0 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothOperand_7), .A1 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_7)) ;
    inv01 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix450 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx449), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_8)) ;
    xnor2 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix452 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx451), .A0 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx453), .A1 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx455)) ;
    xnor2 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix456 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx455), .A0 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothOperand_8), .A1 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_8)) ;
    xor2 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix317 (.Y (
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx316), .A0 (
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx461), .A1 (
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx463)) ;
    xnor2 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix464 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx463), .A0 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothOperand_9), .A1 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_9)) ;
    xor2 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix337 (.Y (
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx336), .A0 (
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx467), .A1 (
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx471)) ;
    inv01 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix470 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx469), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_9)) ;
    xnor2 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix472 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx471), .A0 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothOperand_10), .A1 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_10)) ;
    xor2 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix357 (.Y (
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx356), .A0 (
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx475), .A1 (
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx479)) ;
    inv01 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix478 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx477), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_10)) ;
    xnor2 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix480 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx479), .A0 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothOperand_11), .A1 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_11)) ;
    xor2 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix377 (.Y (
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx376), .A0 (
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx483), .A1 (
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx487)) ;
    inv01 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix486 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx485), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_11)) ;
    xnor2 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix488 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx487), .A0 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothOperand_12), .A1 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_12)) ;
    xor2 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix397 (.Y (
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx396), .A0 (
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx491), .A1 (
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx495)) ;
    inv01 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix494 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx493), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_12)) ;
    xnor2 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix496 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx495), .A0 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothOperand_13), .A1 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_13)) ;
    xor2 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix417 (.Y (
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx416), .A0 (
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx499), .A1 (
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx503)) ;
    inv01 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix502 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx501), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_13)) ;
    xnor2 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix504 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx503), .A0 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothOperand_14), .A1 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_14)) ;
    xor2 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix437 (.Y (
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx436), .A0 (
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx507), .A1 (
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx511)) ;
    inv01 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix510 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx509), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_14)) ;
    xnor2 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix512 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx511), .A0 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothOperand_15), .A1 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_15)) ;
    xnor2 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix457 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx456), .A0 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx515), .A1 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx454)) ;
    inv01 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix518 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx517), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_15)) ;
    xor2 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix455 (.Y (
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx454), .A0 (
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothOperand_16), .A1 (
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_16)) ;
    mux21_ni CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix91 (.Y (
             CALCULATOR_L1FirstOperands_1__0), .A0 (
             CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_1), .A1 (
             CacheWindow_3__4__0), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix99 (.Y (
             CALCULATOR_L1FirstOperands_1__1), .A0 (
             CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_2), .A1 (
             CacheWindow_3__4__1), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix107 (.Y (
             CALCULATOR_L1FirstOperands_1__2), .A0 (
             CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_3), .A1 (
             CacheWindow_3__4__2), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix115 (.Y (
             CALCULATOR_L1FirstOperands_1__3), .A0 (
             CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_4), .A1 (
             CacheWindow_3__4__3), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix123 (.Y (
             CALCULATOR_L1FirstOperands_1__4), .A0 (
             CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_5), .A1 (
             CacheWindow_3__4__4), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix131 (.Y (
             CALCULATOR_L1FirstOperands_1__5), .A0 (
             CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_6), .A1 (
             CacheWindow_3__4__5), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix139 (.Y (
             CALCULATOR_L1FirstOperands_1__6), .A0 (
             CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_7), .A1 (
             CacheWindow_3__4__6), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix147 (.Y (
             CALCULATOR_L1FirstOperands_1__7), .A0 (
             CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_8), .A1 (
             CacheWindow_3__4__7), .S0 (Instr)) ;
    xor2 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix77 (.Y (CALCULATOR_L3Results_0__1), 
         .A0 (CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx529), .A1 (
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx531)) ;
    nand02 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix530 (.Y (
           CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx529), .A0 (
           CALCULATOR_L2Results_1__0), .A1 (CALCULATOR_L2Results_0__0)) ;
    xnor2 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix532 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx531), .A0 (
          CALCULATOR_L2Results_1__1), .A1 (CALCULATOR_L2Results_0__1)) ;
    xor2 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix75 (.Y (CALCULATOR_L3Results_0__2), 
         .A0 (CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx534), .A1 (
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx537)) ;
    aoi32 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix535 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx534), .A0 (
          CALCULATOR_L2Results_1__0), .A1 (CALCULATOR_L2Results_0__0), .A2 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx30), .B0 (CALCULATOR_L2Results_0__1
          ), .B1 (CALCULATOR_L2Results_1__1)) ;
    xnor2 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix538 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx537), .A0 (
          CALCULATOR_L2Results_1__2), .A1 (CALCULATOR_L2Results_0__2)) ;
    xor2 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix73 (.Y (CALCULATOR_L3Results_0__3), 
         .A0 (CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx540), .A1 (
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx544)) ;
    aoi22 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix541 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx540), .A0 (
          CALCULATOR_L2Results_0__2), .A1 (CALCULATOR_L2Results_1__2), .B0 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx40), .B1 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx24)) ;
    xnor2 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix545 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx544), .A0 (
          CALCULATOR_L2Results_1__3), .A1 (CALCULATOR_L2Results_0__3)) ;
    xor2 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix71 (.Y (CALCULATOR_L3Results_0__4), 
         .A0 (CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx547), .A1 (
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx551)) ;
    aoi22 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix548 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx547), .A0 (
          CALCULATOR_L2Results_0__3), .A1 (CALCULATOR_L2Results_1__3), .B0 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx44), .B1 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx18)) ;
    xnor2 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix552 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx551), .A0 (
          CALCULATOR_L2Results_1__4), .A1 (CALCULATOR_L2Results_0__4)) ;
    xor2 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix69 (.Y (CALCULATOR_L3Results_0__5), 
         .A0 (CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx554), .A1 (
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx558)) ;
    aoi22 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix555 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx554), .A0 (
          CALCULATOR_L2Results_0__4), .A1 (CALCULATOR_L2Results_1__4), .B0 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx48), .B1 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx12)) ;
    xnor2 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix559 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx558), .A0 (
          CALCULATOR_L2Results_1__5), .A1 (CALCULATOR_L2Results_0__5)) ;
    xor2 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix67 (.Y (CALCULATOR_L3Results_0__6), 
         .A0 (CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx561), .A1 (
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx565)) ;
    aoi22 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix562 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx561), .A0 (
          CALCULATOR_L2Results_0__5), .A1 (CALCULATOR_L2Results_1__5), .B0 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx52), .B1 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx6)) ;
    xnor2 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix566 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx565), .A0 (
          CALCULATOR_L2Results_1__6), .A1 (CALCULATOR_L2Results_0__6)) ;
    xnor2 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix65 (.Y (CALCULATOR_L3Results_0__7)
          , .A0 (CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx568), .A1 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx62)) ;
    aoi22 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix569 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx568), .A0 (
          CALCULATOR_L2Results_0__6), .A1 (CALCULATOR_L2Results_1__6), .B0 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx56), .B1 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx0)) ;
    xor2 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix63 (.Y (
         CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx62), .A0 (CALCULATOR_L2Results_1__7)
         , .A1 (CALCULATOR_L2Results_0__7)) ;
    inv01 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix155 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx154), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx383)) ;
    inv01 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix57 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx56), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx561)) ;
    inv01 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix53 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx52), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx554)) ;
    inv01 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix49 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx48), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx547)) ;
    inv01 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix45 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx44), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx540)) ;
    inv01 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix41 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx40), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx534)) ;
    inv01 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix31 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx30), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx531)) ;
    inv01 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix25 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx24), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx537)) ;
    inv01 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix19 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx18), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx544)) ;
    inv01 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix13 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx12), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx551)) ;
    inv01 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix7 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx6), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx558)) ;
    inv01 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix1 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx0), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx565)) ;
    fake_gnd CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix216 (.Y (
             CALCULATOR_L1_3_L2_4_G3_MINI_ALU_WindowCellShiftedLeft_16)) ;
    aoi21 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix77 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_10), .A0 (
          CacheFilter_3__4__1), .A1 (CacheFilter_3__4__0), .B0 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_nx4)) ;
    nor02_2x CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix5 (.Y (
             CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_nx4), .A0 (
             CacheFilter_3__4__0), .A1 (CacheFilter_3__4__1)) ;
    aoi21 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix67 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_11), .A0 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_nx328), .A1 (
          CacheFilter_3__4__2), .B0 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_nx8)) ;
    nor03_2x CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix9 (.Y (
             CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_nx8), .A0 (
             CacheFilter_3__4__2), .A1 (CacheFilter_3__4__0), .A2 (
             CacheFilter_3__4__1)) ;
    xnor2 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix59 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_12), .A0 (
          CacheFilter_3__4__3), .A1 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_nx8)) ;
    xnor2 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix51 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_13), .A0 (
          CacheFilter_3__4__4), .A1 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_nx12)) ;
    nor04 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix13 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_nx12), .A0 (
          CacheFilter_3__4__3), .A1 (CacheFilter_3__4__2), .A2 (
          CacheFilter_3__4__0), .A3 (CacheFilter_3__4__1)) ;
    xnor2 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix43 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_14), .A0 (
          CacheFilter_3__4__5), .A1 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_nx16)) ;
    nor02ii CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix17 (.Y (
            CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_nx16), .A0 (
            CacheFilter_3__4__4), .A1 (
            CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_nx12)) ;
    xnor2 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix35 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_15), .A0 (
          CacheFilter_3__4__6), .A1 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_nx20)) ;
    nor02ii CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix21 (.Y (
            CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_nx20), .A0 (
            CacheFilter_3__4__5), .A1 (
            CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_nx16)) ;
    xnor2 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix27 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_16), .A0 (
          CacheFilter_3__4__7), .A1 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_nx24)) ;
    nor02ii CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix25 (.Y (
            CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_nx24), .A0 (
            CacheFilter_3__4__6), .A1 (
            CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_nx20)) ;
    inv01 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix329 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_nx328), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_nx4)) ;
    inv02 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix383 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_nx384), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_0)) ;
    dff CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_0 (.Q (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_0), .QB (
        \$dummy [996]), .D (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .CLK (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    nor02_2x CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix567 (.Y (
             CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566), .A0 (
             RST), .A1 (
             CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644)) ;
    dff CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_1 (.Q (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_1), .QB (
        \$dummy [997]), .D (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .CLK (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_2 (.Q (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_2), .QB (
        \$dummy [998]), .D (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .CLK (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_3 (.Q (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_3), .QB (
        \$dummy [999]), .D (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .CLK (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_4 (.Q (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_4), .QB (
        \$dummy [1000]), .D (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .CLK (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_5 (.Q (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_5), .QB (
        \$dummy [1001]), .D (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .CLK (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_6 (.Q (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_6), .QB (
        \$dummy [1002]), .D (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .CLK (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_7 (.Q (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_7), .QB (
        \$dummy [1003]), .D (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .CLK (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_8 (.Q (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_8), .QB (
        \$dummy [1004]), .D (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .CLK (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_9 (.Q (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_9), .QB (
        \$dummy [1005]), .D (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .CLK (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_10 (.Q (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_10), .QB (
        \$dummy [1006]), .D (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .CLK (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_11 (.Q (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_11), .QB (
        \$dummy [1007]), .D (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .CLK (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_12 (.Q (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_12), .QB (
        \$dummy [1008]), .D (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .CLK (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_13 (.Q (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_13), .QB (
        \$dummy [1009]), .D (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .CLK (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_14 (.Q (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_14), .QB (
        \$dummy [1010]), .D (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .CLK (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_15 (.Q (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_15), .QB (
        \$dummy [1011]), .D (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .CLK (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_16 (.Q (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_16), .QB (
        \$dummy [1012]), .D (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .CLK (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    inv02 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix623 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix625 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix627 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix643 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644), .A (
          nx8139)) ;
    dff CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_0 (.Q (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_0), .QB (
        \$dummy [1013]), .D (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .CLK (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    nor02_2x CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix567 (.Y (
             CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566), .A0 (
             RST), .A1 (
             CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644)) ;
    dff CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_1 (.Q (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_1), .QB (
        \$dummy [1014]), .D (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .CLK (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_2 (.Q (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_2), .QB (
        \$dummy [1015]), .D (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .CLK (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_3 (.Q (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_3), .QB (
        \$dummy [1016]), .D (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .CLK (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_4 (.Q (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_4), .QB (
        \$dummy [1017]), .D (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .CLK (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_5 (.Q (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_5), .QB (
        \$dummy [1018]), .D (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .CLK (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_6 (.Q (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_6), .QB (
        \$dummy [1019]), .D (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .CLK (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_7 (.Q (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_7), .QB (
        \$dummy [1020]), .D (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .CLK (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_8 (.Q (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_8), .QB (
        \$dummy [1021]), .D (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .CLK (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_9 (.Q (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_9), .QB (
        \$dummy [1022]), .D (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .CLK (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_10 (.Q (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_10), .QB (
        \$dummy [1023]), .D (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .CLK (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_11 (.Q (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_11), .QB (
        \$dummy [1024]), .D (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .CLK (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_12 (.Q (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_12), .QB (
        \$dummy [1025]), .D (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .CLK (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_13 (.Q (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_13), .QB (
        \$dummy [1026]), .D (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .CLK (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_14 (.Q (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_14), .QB (
        \$dummy [1027]), .D (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .CLK (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_15 (.Q (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_15), .QB (
        \$dummy [1028]), .D (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .CLK (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_16 (.Q (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_16), .QB (
        \$dummy [1029]), .D (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .CLK (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    inv02 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix623 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix625 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix627 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix643 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644), .A (
          nx8145)) ;
    dff CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_0 (.Q (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_0), .QB (\$dummy [1030]), .D (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .CLK (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    nor02_2x CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix567 (.Y (
             CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566), .A0 (
             RST), .A1 (
             CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    dff CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_1 (.Q (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_1), .QB (\$dummy [1031]), .D (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .CLK (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_2 (.Q (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_2), .QB (\$dummy [1032]), .D (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .CLK (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_3 (.Q (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_3), .QB (\$dummy [1033]), .D (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .CLK (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_4 (.Q (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_4), .QB (\$dummy [1034]), .D (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .CLK (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_5 (.Q (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_5), .QB (\$dummy [1035]), .D (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .CLK (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_6 (.Q (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_6), .QB (\$dummy [1036]), .D (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .CLK (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_7 (.Q (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_7), .QB (\$dummy [1037]), .D (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .CLK (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_8 (.Q (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_8), .QB (\$dummy [1038]), .D (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .CLK (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_9 (.Q (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_9), .QB (\$dummy [1039]), .D (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .CLK (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_10 (.Q (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_10), .QB (\$dummy [1040]), .D (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .CLK (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_11 (.Q (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_11), .QB (\$dummy [1041]), .D (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .CLK (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_12 (.Q (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_12), .QB (\$dummy [1042]), .D (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .CLK (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_13 (.Q (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_13), .QB (\$dummy [1043]), .D (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .CLK (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_14 (.Q (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_14), .QB (\$dummy [1044]), .D (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .CLK (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_15 (.Q (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_15), .QB (\$dummy [1045]), .D (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .CLK (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_16 (.Q (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_16), .QB (\$dummy [1046]), .D (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .CLK (
        CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    inv02 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix623 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix625 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix627 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix643 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642)) ;
    xor2 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix83 (.Y (CALCULATOR_L3Results_1__0), 
         .A0 (CALCULATOR_L2Results_3__0), .A1 (CALCULATOR_L2Results_2__0)) ;
    xnor2 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix380 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx379), .A0 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx381), .A1 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx383)) ;
    nand02 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix382 (.Y (
           CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx381), .A0 (
           CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothOperand_0), .A1 (nx8165)) ;
    xnor2 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix384 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx383), .A0 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothOperand_1), .A1 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_1)) ;
    inv01 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix388 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx387), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_2)) ;
    xnor2 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix390 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx389), .A0 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx391), .A1 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx395)) ;
    aoi32 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix392 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx391), .A0 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothOperand_0), .A1 (nx8165), .A2 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx154), .B0 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_1), .B1 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothOperand_1)) ;
    xnor2 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix396 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx395), .A0 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothOperand_2), .A1 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_2)) ;
    inv01 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix400 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx399), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_3)) ;
    xnor2 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix402 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx401), .A0 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx403), .A1 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx405)) ;
    xnor2 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix406 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx405), .A0 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothOperand_3), .A1 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_3)) ;
    inv01 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix410 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx409), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_4)) ;
    xnor2 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix412 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx411), .A0 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx413), .A1 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx415)) ;
    xnor2 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix416 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx415), .A0 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothOperand_4), .A1 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_4)) ;
    inv01 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix420 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx419), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_5)) ;
    xnor2 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix422 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx421), .A0 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx423), .A1 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx425)) ;
    xnor2 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix426 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx425), .A0 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothOperand_5), .A1 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_5)) ;
    inv01 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix430 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx429), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_6)) ;
    xnor2 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix432 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx431), .A0 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx433), .A1 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx435)) ;
    xnor2 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix436 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx435), .A0 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothOperand_6), .A1 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_6)) ;
    inv01 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix440 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx439), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_7)) ;
    xnor2 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix442 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx441), .A0 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx443), .A1 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx445)) ;
    xnor2 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix446 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx445), .A0 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothOperand_7), .A1 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_7)) ;
    inv01 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix450 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx449), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_8)) ;
    xnor2 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix452 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx451), .A0 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx453), .A1 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx455)) ;
    xnor2 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix456 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx455), .A0 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothOperand_8), .A1 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_8)) ;
    xor2 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix317 (.Y (
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx316), .A0 (
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx461), .A1 (
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx463)) ;
    xnor2 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix464 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx463), .A0 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothOperand_9), .A1 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_9)) ;
    xor2 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix337 (.Y (
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx336), .A0 (
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx467), .A1 (
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx471)) ;
    inv01 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix470 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx469), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_9)) ;
    xnor2 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix472 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx471), .A0 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothOperand_10), .A1 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_10)) ;
    xor2 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix357 (.Y (
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx356), .A0 (
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx475), .A1 (
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx479)) ;
    inv01 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix478 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx477), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_10)) ;
    xnor2 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix480 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx479), .A0 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothOperand_11), .A1 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_11)) ;
    xor2 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix377 (.Y (
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx376), .A0 (
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx483), .A1 (
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx487)) ;
    inv01 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix486 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx485), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_11)) ;
    xnor2 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix488 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx487), .A0 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothOperand_12), .A1 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_12)) ;
    xor2 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix397 (.Y (
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx396), .A0 (
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx491), .A1 (
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx495)) ;
    inv01 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix494 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx493), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_12)) ;
    xnor2 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix496 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx495), .A0 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothOperand_13), .A1 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_13)) ;
    xor2 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix417 (.Y (
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx416), .A0 (
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx499), .A1 (
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx503)) ;
    inv01 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix502 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx501), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_13)) ;
    xnor2 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix504 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx503), .A0 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothOperand_14), .A1 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_14)) ;
    xor2 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix437 (.Y (
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx436), .A0 (
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx507), .A1 (
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx511)) ;
    inv01 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix510 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx509), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_14)) ;
    xnor2 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix512 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx511), .A0 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothOperand_15), .A1 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_15)) ;
    xnor2 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix457 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx456), .A0 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx515), .A1 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx454)) ;
    inv01 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix518 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx517), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_15)) ;
    xor2 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix455 (.Y (
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx454), .A0 (
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothOperand_16), .A1 (
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_16)) ;
    mux21_ni CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix91 (.Y (
             CALCULATOR_L1FirstOperands_5__0), .A0 (
             CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_1), .A1 (
             CacheWindow_4__0__0), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix99 (.Y (
             CALCULATOR_L1FirstOperands_5__1), .A0 (
             CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_2), .A1 (
             CacheWindow_4__0__1), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix107 (.Y (
             CALCULATOR_L1FirstOperands_5__2), .A0 (
             CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_3), .A1 (
             CacheWindow_4__0__2), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix115 (.Y (
             CALCULATOR_L1FirstOperands_5__3), .A0 (
             CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_4), .A1 (
             CacheWindow_4__0__3), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix123 (.Y (
             CALCULATOR_L1FirstOperands_5__4), .A0 (
             CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_5), .A1 (
             CacheWindow_4__0__4), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix131 (.Y (
             CALCULATOR_L1FirstOperands_5__5), .A0 (
             CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_6), .A1 (
             CacheWindow_4__0__5), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix139 (.Y (
             CALCULATOR_L1FirstOperands_5__6), .A0 (
             CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_7), .A1 (
             CacheWindow_4__0__6), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix147 (.Y (
             CALCULATOR_L1FirstOperands_5__7), .A0 (
             CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_8), .A1 (
             CacheWindow_4__0__7), .S0 (Instr)) ;
    xor2 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix77 (.Y (CALCULATOR_L3Results_1__1), 
         .A0 (CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx529), .A1 (
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx531)) ;
    nand02 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix530 (.Y (
           CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx529), .A0 (
           CALCULATOR_L2Results_3__0), .A1 (CALCULATOR_L2Results_2__0)) ;
    xnor2 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix532 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx531), .A0 (
          CALCULATOR_L2Results_3__1), .A1 (CALCULATOR_L2Results_2__1)) ;
    xor2 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix75 (.Y (CALCULATOR_L3Results_1__2), 
         .A0 (CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx534), .A1 (
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx537)) ;
    aoi32 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix535 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx534), .A0 (
          CALCULATOR_L2Results_3__0), .A1 (CALCULATOR_L2Results_2__0), .A2 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx30), .B0 (CALCULATOR_L2Results_2__1
          ), .B1 (CALCULATOR_L2Results_3__1)) ;
    xnor2 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix538 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx537), .A0 (
          CALCULATOR_L2Results_3__2), .A1 (CALCULATOR_L2Results_2__2)) ;
    xor2 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix73 (.Y (CALCULATOR_L3Results_1__3), 
         .A0 (CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx540), .A1 (
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx544)) ;
    aoi22 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix541 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx540), .A0 (
          CALCULATOR_L2Results_2__2), .A1 (CALCULATOR_L2Results_3__2), .B0 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx40), .B1 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx24)) ;
    xnor2 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix545 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx544), .A0 (
          CALCULATOR_L2Results_3__3), .A1 (CALCULATOR_L2Results_2__3)) ;
    xor2 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix71 (.Y (CALCULATOR_L3Results_1__4), 
         .A0 (CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx547), .A1 (
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx551)) ;
    aoi22 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix548 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx547), .A0 (
          CALCULATOR_L2Results_2__3), .A1 (CALCULATOR_L2Results_3__3), .B0 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx44), .B1 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx18)) ;
    xnor2 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix552 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx551), .A0 (
          CALCULATOR_L2Results_3__4), .A1 (CALCULATOR_L2Results_2__4)) ;
    xor2 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix69 (.Y (CALCULATOR_L3Results_1__5), 
         .A0 (CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx554), .A1 (
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx558)) ;
    aoi22 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix555 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx554), .A0 (
          CALCULATOR_L2Results_2__4), .A1 (CALCULATOR_L2Results_3__4), .B0 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx48), .B1 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx12)) ;
    xnor2 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix559 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx558), .A0 (
          CALCULATOR_L2Results_3__5), .A1 (CALCULATOR_L2Results_2__5)) ;
    xor2 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix67 (.Y (CALCULATOR_L3Results_1__6), 
         .A0 (CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx561), .A1 (
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx565)) ;
    aoi22 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix562 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx561), .A0 (
          CALCULATOR_L2Results_2__5), .A1 (CALCULATOR_L2Results_3__5), .B0 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx52), .B1 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx6)) ;
    xnor2 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix566 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx565), .A0 (
          CALCULATOR_L2Results_3__6), .A1 (CALCULATOR_L2Results_2__6)) ;
    xnor2 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix65 (.Y (CALCULATOR_L3Results_1__7)
          , .A0 (CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx568), .A1 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx62)) ;
    aoi22 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix569 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx568), .A0 (
          CALCULATOR_L2Results_2__6), .A1 (CALCULATOR_L2Results_3__6), .B0 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx56), .B1 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx0)) ;
    xor2 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix63 (.Y (
         CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx62), .A0 (CALCULATOR_L2Results_3__7)
         , .A1 (CALCULATOR_L2Results_2__7)) ;
    inv01 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix155 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx154), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx383)) ;
    inv01 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix57 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx56), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx561)) ;
    inv01 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix53 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx52), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx554)) ;
    inv01 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix49 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx48), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx547)) ;
    inv01 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix45 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx44), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx540)) ;
    inv01 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix41 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx40), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx534)) ;
    inv01 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix31 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx30), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx531)) ;
    inv01 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix25 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx24), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx537)) ;
    inv01 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix19 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx18), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx544)) ;
    inv01 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix13 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx12), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx551)) ;
    inv01 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix7 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx6), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx558)) ;
    inv01 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix1 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx0), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx565)) ;
    fake_gnd CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix216 (.Y (
             CALCULATOR_L1_4_L2_0_G3_MINI_ALU_WindowCellShiftedLeft_16)) ;
    aoi21 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix77 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_10), .A0 (
          CacheFilter_4__0__1), .A1 (CacheFilter_4__0__0), .B0 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_nx4)) ;
    nor02_2x CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix5 (.Y (
             CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_nx4), .A0 (
             CacheFilter_4__0__0), .A1 (CacheFilter_4__0__1)) ;
    aoi21 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix67 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_11), .A0 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_nx328), .A1 (
          CacheFilter_4__0__2), .B0 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_nx8)) ;
    nor03_2x CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix9 (.Y (
             CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_nx8), .A0 (
             CacheFilter_4__0__2), .A1 (CacheFilter_4__0__0), .A2 (
             CacheFilter_4__0__1)) ;
    xnor2 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix59 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_12), .A0 (
          CacheFilter_4__0__3), .A1 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_nx8)) ;
    xnor2 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix51 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_13), .A0 (
          CacheFilter_4__0__4), .A1 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_nx12)) ;
    nor04 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix13 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_nx12), .A0 (
          CacheFilter_4__0__3), .A1 (CacheFilter_4__0__2), .A2 (
          CacheFilter_4__0__0), .A3 (CacheFilter_4__0__1)) ;
    xnor2 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix43 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_14), .A0 (
          CacheFilter_4__0__5), .A1 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_nx16)) ;
    nor02ii CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix17 (.Y (
            CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_nx16), .A0 (
            CacheFilter_4__0__4), .A1 (
            CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_nx12)) ;
    xnor2 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix35 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_15), .A0 (
          CacheFilter_4__0__6), .A1 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_nx20)) ;
    nor02ii CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix21 (.Y (
            CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_nx20), .A0 (
            CacheFilter_4__0__5), .A1 (
            CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_nx16)) ;
    xnor2 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix27 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_16), .A0 (
          CacheFilter_4__0__7), .A1 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_nx24)) ;
    nor02ii CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix25 (.Y (
            CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_nx24), .A0 (
            CacheFilter_4__0__6), .A1 (
            CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_nx20)) ;
    inv01 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix329 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_nx328), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_nx4)) ;
    inv02 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix383 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_nx384), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_0)) ;
    dff CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_0 (.Q (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_0), .QB (
        \$dummy [1047]), .D (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .CLK (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    nor02_2x CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix567 (.Y (
             CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566), .A0 (
             RST), .A1 (
             CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644)) ;
    dff CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_1 (.Q (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_1), .QB (
        \$dummy [1048]), .D (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .CLK (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_2 (.Q (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_2), .QB (
        \$dummy [1049]), .D (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .CLK (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_3 (.Q (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_3), .QB (
        \$dummy [1050]), .D (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .CLK (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_4 (.Q (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_4), .QB (
        \$dummy [1051]), .D (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .CLK (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_5 (.Q (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_5), .QB (
        \$dummy [1052]), .D (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .CLK (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_6 (.Q (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_6), .QB (
        \$dummy [1053]), .D (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .CLK (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_7 (.Q (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_7), .QB (
        \$dummy [1054]), .D (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .CLK (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_8 (.Q (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_8), .QB (
        \$dummy [1055]), .D (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .CLK (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_9 (.Q (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_9), .QB (
        \$dummy [1056]), .D (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .CLK (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_10 (.Q (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_10), .QB (
        \$dummy [1057]), .D (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .CLK (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_11 (.Q (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_11), .QB (
        \$dummy [1058]), .D (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .CLK (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_12 (.Q (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_12), .QB (
        \$dummy [1059]), .D (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .CLK (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_13 (.Q (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_13), .QB (
        \$dummy [1060]), .D (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .CLK (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_14 (.Q (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_14), .QB (
        \$dummy [1061]), .D (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .CLK (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_15 (.Q (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_15), .QB (
        \$dummy [1062]), .D (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .CLK (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_16 (.Q (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_16), .QB (
        \$dummy [1063]), .D (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .CLK (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    inv02 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix623 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix625 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix627 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix643 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644), .A (
          nx8179)) ;
    dff CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_0 (.Q (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_0), .QB (
        \$dummy [1064]), .D (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .CLK (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    nor02_2x CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix567 (.Y (
             CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566), .A0 (
             RST), .A1 (
             CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644)) ;
    dff CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_1 (.Q (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_1), .QB (
        \$dummy [1065]), .D (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .CLK (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_2 (.Q (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_2), .QB (
        \$dummy [1066]), .D (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .CLK (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_3 (.Q (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_3), .QB (
        \$dummy [1067]), .D (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .CLK (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_4 (.Q (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_4), .QB (
        \$dummy [1068]), .D (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .CLK (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_5 (.Q (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_5), .QB (
        \$dummy [1069]), .D (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .CLK (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_6 (.Q (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_6), .QB (
        \$dummy [1070]), .D (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .CLK (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_7 (.Q (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_7), .QB (
        \$dummy [1071]), .D (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .CLK (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_8 (.Q (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_8), .QB (
        \$dummy [1072]), .D (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .CLK (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_9 (.Q (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_9), .QB (
        \$dummy [1073]), .D (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .CLK (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_10 (.Q (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_10), .QB (
        \$dummy [1074]), .D (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .CLK (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_11 (.Q (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_11), .QB (
        \$dummy [1075]), .D (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .CLK (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_12 (.Q (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_12), .QB (
        \$dummy [1076]), .D (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .CLK (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_13 (.Q (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_13), .QB (
        \$dummy [1077]), .D (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .CLK (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_14 (.Q (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_14), .QB (
        \$dummy [1078]), .D (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .CLK (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_15 (.Q (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_15), .QB (
        \$dummy [1079]), .D (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .CLK (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_16 (.Q (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_16), .QB (
        \$dummy [1080]), .D (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .CLK (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    inv02 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix623 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix625 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix627 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix643 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644), .A (
          nx8185)) ;
    dff CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_0 (.Q (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_0), .QB (\$dummy [1081]), .D (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .CLK (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    nor02_2x CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix567 (.Y (
             CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566), .A0 (
             RST), .A1 (
             CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    dff CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_1 (.Q (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_1), .QB (\$dummy [1082]), .D (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .CLK (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_2 (.Q (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_2), .QB (\$dummy [1083]), .D (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .CLK (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_3 (.Q (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_3), .QB (\$dummy [1084]), .D (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .CLK (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_4 (.Q (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_4), .QB (\$dummy [1085]), .D (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .CLK (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_5 (.Q (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_5), .QB (\$dummy [1086]), .D (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .CLK (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_6 (.Q (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_6), .QB (\$dummy [1087]), .D (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .CLK (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_7 (.Q (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_7), .QB (\$dummy [1088]), .D (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .CLK (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_8 (.Q (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_8), .QB (\$dummy [1089]), .D (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .CLK (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_9 (.Q (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_9), .QB (\$dummy [1090]), .D (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .CLK (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_10 (.Q (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_10), .QB (\$dummy [1091]), .D (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .CLK (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_11 (.Q (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_11), .QB (\$dummy [1092]), .D (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .CLK (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_12 (.Q (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_12), .QB (\$dummy [1093]), .D (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .CLK (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_13 (.Q (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_13), .QB (\$dummy [1094]), .D (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .CLK (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_14 (.Q (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_14), .QB (\$dummy [1095]), .D (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .CLK (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_15 (.Q (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_15), .QB (\$dummy [1096]), .D (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .CLK (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_16 (.Q (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_16), .QB (\$dummy [1097]), .D (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .CLK (
        CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    inv02 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix623 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix625 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix627 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix643 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642)) ;
    xor2 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix83 (.Y (CALCULATOR_L3Results_2__0), 
         .A0 (CALCULATOR_L2Results_5__0), .A1 (CALCULATOR_L2Results_4__0)) ;
    xnor2 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix380 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx379), .A0 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx381), .A1 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx383)) ;
    nand02 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix382 (.Y (
           CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx381), .A0 (
           CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothOperand_0), .A1 (nx8205)) ;
    xnor2 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix384 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx383), .A0 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothOperand_1), .A1 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_1)) ;
    inv01 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix388 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx387), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_2)) ;
    xnor2 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix390 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx389), .A0 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx391), .A1 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx395)) ;
    aoi32 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix392 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx391), .A0 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothOperand_0), .A1 (nx8205), .A2 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx154), .B0 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_1), .B1 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothOperand_1)) ;
    xnor2 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix396 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx395), .A0 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothOperand_2), .A1 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_2)) ;
    inv01 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix400 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx399), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_3)) ;
    xnor2 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix402 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx401), .A0 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx403), .A1 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx405)) ;
    xnor2 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix406 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx405), .A0 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothOperand_3), .A1 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_3)) ;
    inv01 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix410 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx409), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_4)) ;
    xnor2 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix412 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx411), .A0 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx413), .A1 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx415)) ;
    xnor2 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix416 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx415), .A0 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothOperand_4), .A1 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_4)) ;
    inv01 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix420 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx419), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_5)) ;
    xnor2 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix422 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx421), .A0 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx423), .A1 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx425)) ;
    xnor2 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix426 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx425), .A0 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothOperand_5), .A1 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_5)) ;
    inv01 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix430 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx429), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_6)) ;
    xnor2 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix432 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx431), .A0 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx433), .A1 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx435)) ;
    xnor2 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix436 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx435), .A0 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothOperand_6), .A1 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_6)) ;
    inv01 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix440 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx439), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_7)) ;
    xnor2 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix442 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx441), .A0 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx443), .A1 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx445)) ;
    xnor2 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix446 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx445), .A0 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothOperand_7), .A1 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_7)) ;
    inv01 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix450 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx449), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_8)) ;
    xnor2 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix452 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx451), .A0 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx453), .A1 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx455)) ;
    xnor2 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix456 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx455), .A0 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothOperand_8), .A1 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_8)) ;
    xor2 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix317 (.Y (
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx316), .A0 (
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx461), .A1 (
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx463)) ;
    xnor2 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix464 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx463), .A0 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothOperand_9), .A1 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_9)) ;
    xor2 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix337 (.Y (
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx336), .A0 (
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx467), .A1 (
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx471)) ;
    inv01 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix470 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx469), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_9)) ;
    xnor2 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix472 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx471), .A0 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothOperand_10), .A1 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_10)) ;
    xor2 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix357 (.Y (
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx356), .A0 (
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx475), .A1 (
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx479)) ;
    inv01 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix478 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx477), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_10)) ;
    xnor2 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix480 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx479), .A0 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothOperand_11), .A1 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_11)) ;
    xor2 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix377 (.Y (
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx376), .A0 (
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx483), .A1 (
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx487)) ;
    inv01 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix486 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx485), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_11)) ;
    xnor2 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix488 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx487), .A0 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothOperand_12), .A1 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_12)) ;
    xor2 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix397 (.Y (
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx396), .A0 (
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx491), .A1 (
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx495)) ;
    inv01 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix494 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx493), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_12)) ;
    xnor2 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix496 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx495), .A0 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothOperand_13), .A1 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_13)) ;
    xor2 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix417 (.Y (
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx416), .A0 (
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx499), .A1 (
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx503)) ;
    inv01 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix502 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx501), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_13)) ;
    xnor2 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix504 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx503), .A0 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothOperand_14), .A1 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_14)) ;
    xor2 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix437 (.Y (
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx436), .A0 (
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx507), .A1 (
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx511)) ;
    inv01 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix510 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx509), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_14)) ;
    xnor2 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix512 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx511), .A0 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothOperand_15), .A1 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_15)) ;
    xnor2 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix457 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx456), .A0 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx515), .A1 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx454)) ;
    inv01 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix518 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx517), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_15)) ;
    xor2 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix455 (.Y (
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx454), .A0 (
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothOperand_16), .A1 (
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_16)) ;
    mux21_ni CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix91 (.Y (
             CALCULATOR_L1FirstOperands_9__0), .A0 (
             CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_1), .A1 (
             CacheWindow_4__1__0), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix99 (.Y (
             CALCULATOR_L1FirstOperands_9__1), .A0 (
             CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_2), .A1 (
             CacheWindow_4__1__1), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix107 (.Y (
             CALCULATOR_L1FirstOperands_9__2), .A0 (
             CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_3), .A1 (
             CacheWindow_4__1__2), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix115 (.Y (
             CALCULATOR_L1FirstOperands_9__3), .A0 (
             CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_4), .A1 (
             CacheWindow_4__1__3), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix123 (.Y (
             CALCULATOR_L1FirstOperands_9__4), .A0 (
             CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_5), .A1 (
             CacheWindow_4__1__4), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix131 (.Y (
             CALCULATOR_L1FirstOperands_9__5), .A0 (
             CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_6), .A1 (
             CacheWindow_4__1__5), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix139 (.Y (
             CALCULATOR_L1FirstOperands_9__6), .A0 (
             CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_7), .A1 (
             CacheWindow_4__1__6), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix147 (.Y (
             CALCULATOR_L1FirstOperands_9__7), .A0 (
             CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_8), .A1 (
             CacheWindow_4__1__7), .S0 (Instr)) ;
    xor2 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix77 (.Y (CALCULATOR_L3Results_2__1), 
         .A0 (CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx529), .A1 (
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx531)) ;
    nand02 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix530 (.Y (
           CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx529), .A0 (
           CALCULATOR_L2Results_5__0), .A1 (CALCULATOR_L2Results_4__0)) ;
    xnor2 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix532 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx531), .A0 (
          CALCULATOR_L2Results_5__1), .A1 (CALCULATOR_L2Results_4__1)) ;
    xor2 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix75 (.Y (CALCULATOR_L3Results_2__2), 
         .A0 (CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx534), .A1 (
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx537)) ;
    aoi32 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix535 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx534), .A0 (
          CALCULATOR_L2Results_5__0), .A1 (CALCULATOR_L2Results_4__0), .A2 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx30), .B0 (CALCULATOR_L2Results_4__1
          ), .B1 (CALCULATOR_L2Results_5__1)) ;
    xnor2 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix538 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx537), .A0 (
          CALCULATOR_L2Results_5__2), .A1 (CALCULATOR_L2Results_4__2)) ;
    xor2 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix73 (.Y (CALCULATOR_L3Results_2__3), 
         .A0 (CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx540), .A1 (
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx544)) ;
    aoi22 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix541 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx540), .A0 (
          CALCULATOR_L2Results_4__2), .A1 (CALCULATOR_L2Results_5__2), .B0 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx40), .B1 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx24)) ;
    xnor2 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix545 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx544), .A0 (
          CALCULATOR_L2Results_5__3), .A1 (CALCULATOR_L2Results_4__3)) ;
    xor2 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix71 (.Y (CALCULATOR_L3Results_2__4), 
         .A0 (CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx547), .A1 (
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx551)) ;
    aoi22 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix548 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx547), .A0 (
          CALCULATOR_L2Results_4__3), .A1 (CALCULATOR_L2Results_5__3), .B0 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx44), .B1 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx18)) ;
    xnor2 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix552 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx551), .A0 (
          CALCULATOR_L2Results_5__4), .A1 (CALCULATOR_L2Results_4__4)) ;
    xor2 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix69 (.Y (CALCULATOR_L3Results_2__5), 
         .A0 (CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx554), .A1 (
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx558)) ;
    aoi22 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix555 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx554), .A0 (
          CALCULATOR_L2Results_4__4), .A1 (CALCULATOR_L2Results_5__4), .B0 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx48), .B1 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx12)) ;
    xnor2 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix559 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx558), .A0 (
          CALCULATOR_L2Results_5__5), .A1 (CALCULATOR_L2Results_4__5)) ;
    xor2 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix67 (.Y (CALCULATOR_L3Results_2__6), 
         .A0 (CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx561), .A1 (
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx565)) ;
    aoi22 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix562 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx561), .A0 (
          CALCULATOR_L2Results_4__5), .A1 (CALCULATOR_L2Results_5__5), .B0 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx52), .B1 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx6)) ;
    xnor2 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix566 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx565), .A0 (
          CALCULATOR_L2Results_5__6), .A1 (CALCULATOR_L2Results_4__6)) ;
    xnor2 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix65 (.Y (CALCULATOR_L3Results_2__7)
          , .A0 (CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx568), .A1 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx62)) ;
    aoi22 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix569 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx568), .A0 (
          CALCULATOR_L2Results_4__6), .A1 (CALCULATOR_L2Results_5__6), .B0 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx56), .B1 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx0)) ;
    xor2 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix63 (.Y (
         CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx62), .A0 (CALCULATOR_L2Results_5__7)
         , .A1 (CALCULATOR_L2Results_4__7)) ;
    inv01 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix155 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx154), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx383)) ;
    inv01 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix57 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx56), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx561)) ;
    inv01 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix53 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx52), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx554)) ;
    inv01 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix49 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx48), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx547)) ;
    inv01 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix45 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx44), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx540)) ;
    inv01 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix41 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx40), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx534)) ;
    inv01 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix31 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx30), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx531)) ;
    inv01 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix25 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx24), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx537)) ;
    inv01 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix19 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx18), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx544)) ;
    inv01 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix13 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx12), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx551)) ;
    inv01 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix7 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx6), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx558)) ;
    inv01 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix1 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx0), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx565)) ;
    fake_gnd CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix216 (.Y (
             CALCULATOR_L1_4_L2_1_G3_MINI_ALU_WindowCellShiftedLeft_16)) ;
    aoi21 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix77 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_10), .A0 (
          CacheFilter_4__1__1), .A1 (CacheFilter_4__1__0), .B0 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_nx4)) ;
    nor02_2x CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix5 (.Y (
             CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_nx4), .A0 (
             CacheFilter_4__1__0), .A1 (CacheFilter_4__1__1)) ;
    aoi21 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix67 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_11), .A0 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_nx328), .A1 (
          CacheFilter_4__1__2), .B0 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_nx8)) ;
    nor03_2x CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix9 (.Y (
             CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_nx8), .A0 (
             CacheFilter_4__1__2), .A1 (CacheFilter_4__1__0), .A2 (
             CacheFilter_4__1__1)) ;
    xnor2 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix59 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_12), .A0 (
          CacheFilter_4__1__3), .A1 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_nx8)) ;
    xnor2 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix51 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_13), .A0 (
          CacheFilter_4__1__4), .A1 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_nx12)) ;
    nor04 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix13 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_nx12), .A0 (
          CacheFilter_4__1__3), .A1 (CacheFilter_4__1__2), .A2 (
          CacheFilter_4__1__0), .A3 (CacheFilter_4__1__1)) ;
    xnor2 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix43 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_14), .A0 (
          CacheFilter_4__1__5), .A1 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_nx16)) ;
    nor02ii CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix17 (.Y (
            CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_nx16), .A0 (
            CacheFilter_4__1__4), .A1 (
            CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_nx12)) ;
    xnor2 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix35 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_15), .A0 (
          CacheFilter_4__1__6), .A1 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_nx20)) ;
    nor02ii CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix21 (.Y (
            CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_nx20), .A0 (
            CacheFilter_4__1__5), .A1 (
            CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_nx16)) ;
    xnor2 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix27 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_16), .A0 (
          CacheFilter_4__1__7), .A1 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_nx24)) ;
    nor02ii CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix25 (.Y (
            CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_nx24), .A0 (
            CacheFilter_4__1__6), .A1 (
            CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_nx20)) ;
    inv01 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix329 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_nx328), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_nx4)) ;
    inv02 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix383 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_nx384), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_0)) ;
    dff CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_0 (.Q (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_0), .QB (
        \$dummy [1098]), .D (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .CLK (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    nor02_2x CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix567 (.Y (
             CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566), .A0 (
             RST), .A1 (
             CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644)) ;
    dff CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_1 (.Q (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_1), .QB (
        \$dummy [1099]), .D (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .CLK (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_2 (.Q (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_2), .QB (
        \$dummy [1100]), .D (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .CLK (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_3 (.Q (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_3), .QB (
        \$dummy [1101]), .D (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .CLK (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_4 (.Q (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_4), .QB (
        \$dummy [1102]), .D (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .CLK (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_5 (.Q (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_5), .QB (
        \$dummy [1103]), .D (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .CLK (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_6 (.Q (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_6), .QB (
        \$dummy [1104]), .D (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .CLK (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_7 (.Q (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_7), .QB (
        \$dummy [1105]), .D (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .CLK (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_8 (.Q (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_8), .QB (
        \$dummy [1106]), .D (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .CLK (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_9 (.Q (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_9), .QB (
        \$dummy [1107]), .D (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .CLK (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_10 (.Q (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_10), .QB (
        \$dummy [1108]), .D (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .CLK (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_11 (.Q (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_11), .QB (
        \$dummy [1109]), .D (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .CLK (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_12 (.Q (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_12), .QB (
        \$dummy [1110]), .D (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .CLK (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_13 (.Q (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_13), .QB (
        \$dummy [1111]), .D (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .CLK (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_14 (.Q (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_14), .QB (
        \$dummy [1112]), .D (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .CLK (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_15 (.Q (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_15), .QB (
        \$dummy [1113]), .D (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .CLK (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_16 (.Q (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_16), .QB (
        \$dummy [1114]), .D (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .CLK (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    inv02 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix623 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix625 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix627 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix643 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644), .A (
          nx8219)) ;
    dff CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_0 (.Q (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_0), .QB (
        \$dummy [1115]), .D (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .CLK (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    nor02_2x CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix567 (.Y (
             CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566), .A0 (
             RST), .A1 (
             CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644)) ;
    dff CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_1 (.Q (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_1), .QB (
        \$dummy [1116]), .D (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .CLK (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_2 (.Q (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_2), .QB (
        \$dummy [1117]), .D (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .CLK (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_3 (.Q (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_3), .QB (
        \$dummy [1118]), .D (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .CLK (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_4 (.Q (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_4), .QB (
        \$dummy [1119]), .D (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .CLK (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_5 (.Q (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_5), .QB (
        \$dummy [1120]), .D (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .CLK (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_6 (.Q (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_6), .QB (
        \$dummy [1121]), .D (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .CLK (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_7 (.Q (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_7), .QB (
        \$dummy [1122]), .D (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .CLK (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_8 (.Q (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_8), .QB (
        \$dummy [1123]), .D (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .CLK (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_9 (.Q (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_9), .QB (
        \$dummy [1124]), .D (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .CLK (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_10 (.Q (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_10), .QB (
        \$dummy [1125]), .D (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .CLK (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_11 (.Q (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_11), .QB (
        \$dummy [1126]), .D (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .CLK (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_12 (.Q (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_12), .QB (
        \$dummy [1127]), .D (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .CLK (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_13 (.Q (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_13), .QB (
        \$dummy [1128]), .D (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .CLK (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_14 (.Q (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_14), .QB (
        \$dummy [1129]), .D (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .CLK (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_15 (.Q (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_15), .QB (
        \$dummy [1130]), .D (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .CLK (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_16 (.Q (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_16), .QB (
        \$dummy [1131]), .D (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .CLK (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    inv02 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix623 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix625 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix627 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix643 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644), .A (
          nx8225)) ;
    dff CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_0 (.Q (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_0), .QB (\$dummy [1132]), .D (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .CLK (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    nor02_2x CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix567 (.Y (
             CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566), .A0 (
             RST), .A1 (
             CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    dff CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_1 (.Q (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_1), .QB (\$dummy [1133]), .D (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .CLK (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_2 (.Q (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_2), .QB (\$dummy [1134]), .D (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .CLK (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_3 (.Q (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_3), .QB (\$dummy [1135]), .D (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .CLK (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_4 (.Q (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_4), .QB (\$dummy [1136]), .D (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .CLK (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_5 (.Q (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_5), .QB (\$dummy [1137]), .D (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .CLK (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_6 (.Q (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_6), .QB (\$dummy [1138]), .D (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .CLK (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_7 (.Q (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_7), .QB (\$dummy [1139]), .D (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .CLK (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_8 (.Q (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_8), .QB (\$dummy [1140]), .D (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .CLK (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_9 (.Q (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_9), .QB (\$dummy [1141]), .D (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .CLK (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_10 (.Q (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_10), .QB (\$dummy [1142]), .D (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .CLK (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_11 (.Q (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_11), .QB (\$dummy [1143]), .D (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .CLK (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_12 (.Q (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_12), .QB (\$dummy [1144]), .D (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .CLK (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_13 (.Q (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_13), .QB (\$dummy [1145]), .D (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .CLK (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_14 (.Q (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_14), .QB (\$dummy [1146]), .D (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .CLK (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_15 (.Q (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_15), .QB (\$dummy [1147]), .D (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .CLK (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_16 (.Q (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_16), .QB (\$dummy [1148]), .D (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .CLK (
        CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    inv02 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix623 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix625 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix627 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix643 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642)) ;
    xor2 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix83 (.Y (CALCULATOR_L4Results_0__0), 
         .A0 (CALCULATOR_L3Results_1__0), .A1 (CALCULATOR_L3Results_0__0)) ;
    xnor2 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix380 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx379), .A0 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx381), .A1 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx383)) ;
    nand02 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix382 (.Y (
           CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx381), .A0 (
           CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothOperand_0), .A1 (nx8245)) ;
    xnor2 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix384 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx383), .A0 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothOperand_1), .A1 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_1)) ;
    inv01 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix388 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx387), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_2)) ;
    xnor2 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix390 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx389), .A0 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx391), .A1 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx395)) ;
    aoi32 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix392 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx391), .A0 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothOperand_0), .A1 (nx8245), .A2 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx154), .B0 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_1), .B1 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothOperand_1)) ;
    xnor2 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix396 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx395), .A0 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothOperand_2), .A1 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_2)) ;
    inv01 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix400 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx399), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_3)) ;
    xnor2 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix402 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx401), .A0 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx403), .A1 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx405)) ;
    xnor2 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix406 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx405), .A0 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothOperand_3), .A1 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_3)) ;
    inv01 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix410 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx409), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_4)) ;
    xnor2 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix412 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx411), .A0 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx413), .A1 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx415)) ;
    xnor2 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix416 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx415), .A0 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothOperand_4), .A1 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_4)) ;
    inv01 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix420 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx419), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_5)) ;
    xnor2 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix422 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx421), .A0 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx423), .A1 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx425)) ;
    xnor2 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix426 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx425), .A0 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothOperand_5), .A1 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_5)) ;
    inv01 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix430 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx429), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_6)) ;
    xnor2 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix432 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx431), .A0 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx433), .A1 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx435)) ;
    xnor2 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix436 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx435), .A0 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothOperand_6), .A1 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_6)) ;
    inv01 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix440 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx439), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_7)) ;
    xnor2 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix442 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx441), .A0 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx443), .A1 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx445)) ;
    xnor2 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix446 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx445), .A0 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothOperand_7), .A1 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_7)) ;
    inv01 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix450 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx449), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_8)) ;
    xnor2 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix452 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx451), .A0 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx453), .A1 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx455)) ;
    xnor2 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix456 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx455), .A0 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothOperand_8), .A1 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_8)) ;
    xor2 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix317 (.Y (
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx316), .A0 (
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx461), .A1 (
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx463)) ;
    xnor2 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix464 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx463), .A0 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothOperand_9), .A1 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_9)) ;
    xor2 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix337 (.Y (
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx336), .A0 (
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx467), .A1 (
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx471)) ;
    inv01 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix470 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx469), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_9)) ;
    xnor2 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix472 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx471), .A0 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothOperand_10), .A1 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_10)) ;
    xor2 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix357 (.Y (
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx356), .A0 (
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx475), .A1 (
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx479)) ;
    inv01 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix478 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx477), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_10)) ;
    xnor2 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix480 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx479), .A0 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothOperand_11), .A1 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_11)) ;
    xor2 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix377 (.Y (
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx376), .A0 (
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx483), .A1 (
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx487)) ;
    inv01 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix486 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx485), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_11)) ;
    xnor2 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix488 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx487), .A0 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothOperand_12), .A1 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_12)) ;
    xor2 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix397 (.Y (
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx396), .A0 (
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx491), .A1 (
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx495)) ;
    inv01 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix494 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx493), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_12)) ;
    xnor2 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix496 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx495), .A0 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothOperand_13), .A1 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_13)) ;
    xor2 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix417 (.Y (
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx416), .A0 (
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx499), .A1 (
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx503)) ;
    inv01 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix502 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx501), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_13)) ;
    xnor2 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix504 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx503), .A0 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothOperand_14), .A1 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_14)) ;
    xor2 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix437 (.Y (
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx436), .A0 (
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx507), .A1 (
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx511)) ;
    inv01 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix510 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx509), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_14)) ;
    xnor2 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix512 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx511), .A0 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothOperand_15), .A1 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_15)) ;
    xnor2 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix457 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx456), .A0 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx515), .A1 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx454)) ;
    inv01 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix518 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx517), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_15)) ;
    xor2 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix455 (.Y (
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx454), .A0 (
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothOperand_16), .A1 (
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_16)) ;
    mux21_ni CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix91 (.Y (
             CALCULATOR_L1FirstOperands_3__0), .A0 (
             CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_1), .A1 (
             CacheWindow_4__2__0), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix99 (.Y (
             CALCULATOR_L1FirstOperands_3__1), .A0 (
             CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_2), .A1 (
             CacheWindow_4__2__1), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix107 (.Y (
             CALCULATOR_L1FirstOperands_3__2), .A0 (
             CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_3), .A1 (
             CacheWindow_4__2__2), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix115 (.Y (
             CALCULATOR_L1FirstOperands_3__3), .A0 (
             CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_4), .A1 (
             CacheWindow_4__2__3), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix123 (.Y (
             CALCULATOR_L1FirstOperands_3__4), .A0 (
             CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_5), .A1 (
             CacheWindow_4__2__4), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix131 (.Y (
             CALCULATOR_L1FirstOperands_3__5), .A0 (
             CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_6), .A1 (
             CacheWindow_4__2__5), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix139 (.Y (
             CALCULATOR_L1FirstOperands_3__6), .A0 (
             CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_7), .A1 (
             CacheWindow_4__2__6), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix147 (.Y (
             CALCULATOR_L1FirstOperands_3__7), .A0 (
             CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_8), .A1 (
             CacheWindow_4__2__7), .S0 (Instr)) ;
    xor2 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix77 (.Y (CALCULATOR_L4Results_0__1), 
         .A0 (CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx529), .A1 (
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx531)) ;
    nand02 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix530 (.Y (
           CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx529), .A0 (
           CALCULATOR_L3Results_1__0), .A1 (CALCULATOR_L3Results_0__0)) ;
    xnor2 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix532 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx531), .A0 (
          CALCULATOR_L3Results_1__1), .A1 (CALCULATOR_L3Results_0__1)) ;
    xor2 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix75 (.Y (CALCULATOR_L4Results_0__2), 
         .A0 (CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx534), .A1 (
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx537)) ;
    aoi32 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix535 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx534), .A0 (
          CALCULATOR_L3Results_1__0), .A1 (CALCULATOR_L3Results_0__0), .A2 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx30), .B0 (CALCULATOR_L3Results_0__1
          ), .B1 (CALCULATOR_L3Results_1__1)) ;
    xnor2 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix538 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx537), .A0 (
          CALCULATOR_L3Results_1__2), .A1 (CALCULATOR_L3Results_0__2)) ;
    xor2 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix73 (.Y (CALCULATOR_L4Results_0__3), 
         .A0 (CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx540), .A1 (
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx544)) ;
    aoi22 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix541 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx540), .A0 (
          CALCULATOR_L3Results_0__2), .A1 (CALCULATOR_L3Results_1__2), .B0 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx40), .B1 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx24)) ;
    xnor2 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix545 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx544), .A0 (
          CALCULATOR_L3Results_1__3), .A1 (CALCULATOR_L3Results_0__3)) ;
    xor2 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix71 (.Y (CALCULATOR_L4Results_0__4), 
         .A0 (CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx547), .A1 (
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx551)) ;
    aoi22 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix548 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx547), .A0 (
          CALCULATOR_L3Results_0__3), .A1 (CALCULATOR_L3Results_1__3), .B0 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx44), .B1 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx18)) ;
    xnor2 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix552 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx551), .A0 (
          CALCULATOR_L3Results_1__4), .A1 (CALCULATOR_L3Results_0__4)) ;
    xor2 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix69 (.Y (CALCULATOR_L4Results_0__5), 
         .A0 (CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx554), .A1 (
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx558)) ;
    aoi22 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix555 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx554), .A0 (
          CALCULATOR_L3Results_0__4), .A1 (CALCULATOR_L3Results_1__4), .B0 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx48), .B1 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx12)) ;
    xnor2 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix559 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx558), .A0 (
          CALCULATOR_L3Results_1__5), .A1 (CALCULATOR_L3Results_0__5)) ;
    xor2 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix67 (.Y (CALCULATOR_L4Results_0__6), 
         .A0 (CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx561), .A1 (
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx565)) ;
    aoi22 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix562 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx561), .A0 (
          CALCULATOR_L3Results_0__5), .A1 (CALCULATOR_L3Results_1__5), .B0 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx52), .B1 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx6)) ;
    xnor2 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix566 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx565), .A0 (
          CALCULATOR_L3Results_1__6), .A1 (CALCULATOR_L3Results_0__6)) ;
    xnor2 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix65 (.Y (CALCULATOR_L4Results_0__7)
          , .A0 (CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx568), .A1 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx62)) ;
    aoi22 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix569 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx568), .A0 (
          CALCULATOR_L3Results_0__6), .A1 (CALCULATOR_L3Results_1__6), .B0 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx56), .B1 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx0)) ;
    xor2 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix63 (.Y (
         CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx62), .A0 (CALCULATOR_L3Results_1__7)
         , .A1 (CALCULATOR_L3Results_0__7)) ;
    inv01 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix155 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx154), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx383)) ;
    inv01 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix57 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx56), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx561)) ;
    inv01 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix53 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx52), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx554)) ;
    inv01 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix49 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx48), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx547)) ;
    inv01 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix45 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx44), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx540)) ;
    inv01 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix41 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx40), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx534)) ;
    inv01 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix31 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx30), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx531)) ;
    inv01 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix25 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx24), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx537)) ;
    inv01 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix19 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx18), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx544)) ;
    inv01 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix13 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx12), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx551)) ;
    inv01 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix7 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx6), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx558)) ;
    inv01 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix1 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx0), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx565)) ;
    fake_gnd CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix216 (.Y (
             CALCULATOR_L1_4_L2_2_G4_MINI_ALU_WindowCellShiftedLeft_16)) ;
    aoi21 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix77 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDin_10), .A0 (
          CacheFilter_4__2__1), .A1 (CacheFilter_4__2__0), .B0 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_nx4)) ;
    nor02_2x CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix5 (.Y (
             CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_nx4), .A0 (
             CacheFilter_4__2__0), .A1 (CacheFilter_4__2__1)) ;
    aoi21 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix67 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDin_11), .A0 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_nx328), .A1 (
          CacheFilter_4__2__2), .B0 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_nx8)) ;
    nor03_2x CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix9 (.Y (
             CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_nx8), .A0 (
             CacheFilter_4__2__2), .A1 (CacheFilter_4__2__0), .A2 (
             CacheFilter_4__2__1)) ;
    xnor2 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix59 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDin_12), .A0 (
          CacheFilter_4__2__3), .A1 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_nx8)) ;
    xnor2 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix51 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDin_13), .A0 (
          CacheFilter_4__2__4), .A1 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_nx12)) ;
    nor04 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix13 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_nx12), .A0 (
          CacheFilter_4__2__3), .A1 (CacheFilter_4__2__2), .A2 (
          CacheFilter_4__2__0), .A3 (CacheFilter_4__2__1)) ;
    xnor2 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix43 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDin_14), .A0 (
          CacheFilter_4__2__5), .A1 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_nx16)) ;
    nor02ii CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix17 (.Y (
            CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_nx16), .A0 (
            CacheFilter_4__2__4), .A1 (
            CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_nx12)) ;
    xnor2 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix35 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDin_15), .A0 (
          CacheFilter_4__2__6), .A1 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_nx20)) ;
    nor02ii CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix21 (.Y (
            CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_nx20), .A0 (
            CacheFilter_4__2__5), .A1 (
            CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_nx16)) ;
    xnor2 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix27 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDin_16), .A0 (
          CacheFilter_4__2__7), .A1 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_nx24)) ;
    nor02ii CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix25 (.Y (
            CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_nx24), .A0 (
            CacheFilter_4__2__6), .A1 (
            CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_nx20)) ;
    inv01 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix329 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_nx328), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_nx4)) ;
    inv02 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix383 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_nx384), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_0)) ;
    dff CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_0 (.Q (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_0), .QB (
        \$dummy [1149]), .D (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .CLK (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    nor02_2x CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix567 (.Y (
             CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566), .A0 (
             RST), .A1 (
             CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644)) ;
    dff CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_1 (.Q (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_1), .QB (
        \$dummy [1150]), .D (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .CLK (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_2 (.Q (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_2), .QB (
        \$dummy [1151]), .D (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .CLK (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_3 (.Q (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_3), .QB (
        \$dummy [1152]), .D (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .CLK (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_4 (.Q (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_4), .QB (
        \$dummy [1153]), .D (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .CLK (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_5 (.Q (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_5), .QB (
        \$dummy [1154]), .D (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .CLK (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_6 (.Q (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_6), .QB (
        \$dummy [1155]), .D (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .CLK (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_7 (.Q (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_7), .QB (
        \$dummy [1156]), .D (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .CLK (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_8 (.Q (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_8), .QB (
        \$dummy [1157]), .D (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .CLK (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_9 (.Q (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_9), .QB (
        \$dummy [1158]), .D (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .CLK (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_10 (.Q (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_10), .QB (
        \$dummy [1159]), .D (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .CLK (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_11 (.Q (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_11), .QB (
        \$dummy [1160]), .D (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .CLK (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_12 (.Q (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_12), .QB (
        \$dummy [1161]), .D (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .CLK (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_13 (.Q (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_13), .QB (
        \$dummy [1162]), .D (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .CLK (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_14 (.Q (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_14), .QB (
        \$dummy [1163]), .D (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .CLK (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_15 (.Q (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_15), .QB (
        \$dummy [1164]), .D (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .CLK (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_16 (.Q (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_16), .QB (
        \$dummy [1165]), .D (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .CLK (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    inv02 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix623 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix625 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix627 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix643 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644), .A (
          nx8259)) ;
    dff CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_0 (.Q (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_0), .QB (
        \$dummy [1166]), .D (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .CLK (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    nor02_2x CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix567 (.Y (
             CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566), .A0 (
             RST), .A1 (
             CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644)) ;
    dff CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_1 (.Q (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_1), .QB (
        \$dummy [1167]), .D (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .CLK (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_2 (.Q (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_2), .QB (
        \$dummy [1168]), .D (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .CLK (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_3 (.Q (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_3), .QB (
        \$dummy [1169]), .D (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .CLK (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_4 (.Q (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_4), .QB (
        \$dummy [1170]), .D (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .CLK (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_5 (.Q (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_5), .QB (
        \$dummy [1171]), .D (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .CLK (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_6 (.Q (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_6), .QB (
        \$dummy [1172]), .D (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .CLK (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_7 (.Q (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_7), .QB (
        \$dummy [1173]), .D (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .CLK (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_8 (.Q (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_8), .QB (
        \$dummy [1174]), .D (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .CLK (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_9 (.Q (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_9), .QB (
        \$dummy [1175]), .D (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .CLK (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_10 (.Q (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_10), .QB (
        \$dummy [1176]), .D (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .CLK (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_11 (.Q (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_11), .QB (
        \$dummy [1177]), .D (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .CLK (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_12 (.Q (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_12), .QB (
        \$dummy [1178]), .D (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .CLK (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_13 (.Q (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_13), .QB (
        \$dummy [1179]), .D (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .CLK (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_14 (.Q (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_14), .QB (
        \$dummy [1180]), .D (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .CLK (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_15 (.Q (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_15), .QB (
        \$dummy [1181]), .D (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .CLK (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_16 (.Q (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_16), .QB (
        \$dummy [1182]), .D (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .CLK (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    inv02 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix623 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix625 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix627 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix643 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644), .A (
          nx8265)) ;
    dff CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_0 (.Q (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_0), .QB (\$dummy [1183]), .D (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .CLK (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    nor02_2x CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix567 (.Y (
             CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566), .A0 (
             RST), .A1 (
             CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    dff CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_1 (.Q (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_1), .QB (\$dummy [1184]), .D (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .CLK (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_2 (.Q (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_2), .QB (\$dummy [1185]), .D (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .CLK (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_3 (.Q (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_3), .QB (\$dummy [1186]), .D (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .CLK (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_4 (.Q (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_4), .QB (\$dummy [1187]), .D (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .CLK (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_5 (.Q (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_5), .QB (\$dummy [1188]), .D (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .CLK (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_6 (.Q (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_6), .QB (\$dummy [1189]), .D (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .CLK (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_7 (.Q (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_7), .QB (\$dummy [1190]), .D (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .CLK (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_8 (.Q (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_8), .QB (\$dummy [1191]), .D (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .CLK (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_9 (.Q (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_9), .QB (\$dummy [1192]), .D (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .CLK (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_10 (.Q (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_10), .QB (\$dummy [1193]), .D (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .CLK (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_11 (.Q (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_11), .QB (\$dummy [1194]), .D (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .CLK (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_12 (.Q (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_12), .QB (\$dummy [1195]), .D (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .CLK (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_13 (.Q (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_13), .QB (\$dummy [1196]), .D (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .CLK (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_14 (.Q (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_14), .QB (\$dummy [1197]), .D (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .CLK (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_15 (.Q (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_15), .QB (\$dummy [1198]), .D (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .CLK (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_16 (.Q (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_16), .QB (\$dummy [1199]), .D (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .CLK (
        CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    inv02 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix623 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix625 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix627 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix643 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642)) ;
    xor2 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix83 (.Y (
         CALCULATOR_L5FirstOperands_1__0), .A0 (CALCULATOR_L3Results_2__0), .A1 (
         CALCULATOR_L4Results_0__0)) ;
    xnor2 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix380 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx379), .A0 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx381), .A1 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx383)) ;
    nand02 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix382 (.Y (
           CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx381), .A0 (
           CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothOperand_0), .A1 (nx8285)) ;
    xnor2 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix384 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx383), .A0 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothOperand_1), .A1 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_1)) ;
    inv01 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix388 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx387), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_2)) ;
    xnor2 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix390 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx389), .A0 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx391), .A1 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx395)) ;
    aoi32 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix392 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx391), .A0 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothOperand_0), .A1 (nx8285), .A2 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx154), .B0 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_1), .B1 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothOperand_1)) ;
    xnor2 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix396 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx395), .A0 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothOperand_2), .A1 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_2)) ;
    inv01 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix400 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx399), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_3)) ;
    xnor2 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix402 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx401), .A0 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx403), .A1 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx405)) ;
    xnor2 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix406 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx405), .A0 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothOperand_3), .A1 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_3)) ;
    inv01 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix410 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx409), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_4)) ;
    xnor2 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix412 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx411), .A0 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx413), .A1 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx415)) ;
    xnor2 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix416 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx415), .A0 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothOperand_4), .A1 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_4)) ;
    inv01 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix420 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx419), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_5)) ;
    xnor2 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix422 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx421), .A0 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx423), .A1 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx425)) ;
    xnor2 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix426 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx425), .A0 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothOperand_5), .A1 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_5)) ;
    inv01 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix430 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx429), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_6)) ;
    xnor2 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix432 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx431), .A0 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx433), .A1 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx435)) ;
    xnor2 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix436 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx435), .A0 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothOperand_6), .A1 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_6)) ;
    inv01 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix440 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx439), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_7)) ;
    xnor2 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix442 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx441), .A0 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx443), .A1 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx445)) ;
    xnor2 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix446 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx445), .A0 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothOperand_7), .A1 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_7)) ;
    inv01 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix450 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx449), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_8)) ;
    xnor2 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix452 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx451), .A0 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx453), .A1 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx455)) ;
    xnor2 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix456 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx455), .A0 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothOperand_8), .A1 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_8)) ;
    xor2 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix317 (.Y (
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx316), .A0 (
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx461), .A1 (
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx463)) ;
    xnor2 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix464 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx463), .A0 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothOperand_9), .A1 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_9)) ;
    xor2 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix337 (.Y (
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx336), .A0 (
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx467), .A1 (
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx471)) ;
    inv01 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix470 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx469), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_9)) ;
    xnor2 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix472 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx471), .A0 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothOperand_10), .A1 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_10)) ;
    xor2 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix357 (.Y (
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx356), .A0 (
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx475), .A1 (
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx479)) ;
    inv01 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix478 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx477), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_10)) ;
    xnor2 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix480 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx479), .A0 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothOperand_11), .A1 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_11)) ;
    xor2 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix377 (.Y (
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx376), .A0 (
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx483), .A1 (
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx487)) ;
    inv01 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix486 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx485), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_11)) ;
    xnor2 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix488 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx487), .A0 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothOperand_12), .A1 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_12)) ;
    xor2 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix397 (.Y (
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx396), .A0 (
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx491), .A1 (
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx495)) ;
    inv01 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix494 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx493), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_12)) ;
    xnor2 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix496 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx495), .A0 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothOperand_13), .A1 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_13)) ;
    xor2 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix417 (.Y (
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx416), .A0 (
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx499), .A1 (
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx503)) ;
    inv01 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix502 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx501), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_13)) ;
    xnor2 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix504 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx503), .A0 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothOperand_14), .A1 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_14)) ;
    xor2 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix437 (.Y (
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx436), .A0 (
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx507), .A1 (
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx511)) ;
    inv01 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix510 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx509), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_14)) ;
    xnor2 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix512 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx511), .A0 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothOperand_15), .A1 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_15)) ;
    xnor2 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix457 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx456), .A0 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx515), .A1 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx454)) ;
    inv01 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix518 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx517), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_15)) ;
    xor2 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix455 (.Y (
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx454), .A0 (
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothOperand_16), .A1 (
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_16)) ;
    mux21_ni CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix91 (.Y (
             CALCULATOR_L1FirstOperands_7__0), .A0 (
             CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_1), .A1 (
             CacheWindow_4__3__0), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix99 (.Y (
             CALCULATOR_L1FirstOperands_7__1), .A0 (
             CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_2), .A1 (
             CacheWindow_4__3__1), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix107 (.Y (
             CALCULATOR_L1FirstOperands_7__2), .A0 (
             CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_3), .A1 (
             CacheWindow_4__3__2), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix115 (.Y (
             CALCULATOR_L1FirstOperands_7__3), .A0 (
             CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_4), .A1 (
             CacheWindow_4__3__3), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix123 (.Y (
             CALCULATOR_L1FirstOperands_7__4), .A0 (
             CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_5), .A1 (
             CacheWindow_4__3__4), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix131 (.Y (
             CALCULATOR_L1FirstOperands_7__5), .A0 (
             CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_6), .A1 (
             CacheWindow_4__3__5), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix139 (.Y (
             CALCULATOR_L1FirstOperands_7__6), .A0 (
             CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_7), .A1 (
             CacheWindow_4__3__6), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix147 (.Y (
             CALCULATOR_L1FirstOperands_7__7), .A0 (
             CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_8), .A1 (
             CacheWindow_4__3__7), .S0 (Instr)) ;
    xor2 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix77 (.Y (
         CALCULATOR_L5FirstOperands_1__1), .A0 (
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx529), .A1 (
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx531)) ;
    nand02 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix530 (.Y (
           CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx529), .A0 (
           CALCULATOR_L3Results_2__0), .A1 (CALCULATOR_L4Results_0__0)) ;
    xnor2 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix532 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx531), .A0 (
          CALCULATOR_L3Results_2__1), .A1 (CALCULATOR_L4Results_0__1)) ;
    xor2 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix75 (.Y (
         CALCULATOR_L5FirstOperands_1__2), .A0 (
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx534), .A1 (
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx537)) ;
    aoi32 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix535 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx534), .A0 (
          CALCULATOR_L3Results_2__0), .A1 (CALCULATOR_L4Results_0__0), .A2 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx30), .B0 (CALCULATOR_L4Results_0__1
          ), .B1 (CALCULATOR_L3Results_2__1)) ;
    xnor2 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix538 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx537), .A0 (
          CALCULATOR_L3Results_2__2), .A1 (CALCULATOR_L4Results_0__2)) ;
    xor2 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix73 (.Y (
         CALCULATOR_L5FirstOperands_1__3), .A0 (
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx540), .A1 (
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx544)) ;
    aoi22 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix541 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx540), .A0 (
          CALCULATOR_L4Results_0__2), .A1 (CALCULATOR_L3Results_2__2), .B0 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx40), .B1 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx24)) ;
    xnor2 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix545 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx544), .A0 (
          CALCULATOR_L3Results_2__3), .A1 (CALCULATOR_L4Results_0__3)) ;
    xor2 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix71 (.Y (
         CALCULATOR_L5FirstOperands_1__4), .A0 (
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx547), .A1 (
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx551)) ;
    aoi22 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix548 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx547), .A0 (
          CALCULATOR_L4Results_0__3), .A1 (CALCULATOR_L3Results_2__3), .B0 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx44), .B1 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx18)) ;
    xnor2 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix552 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx551), .A0 (
          CALCULATOR_L3Results_2__4), .A1 (CALCULATOR_L4Results_0__4)) ;
    xor2 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix69 (.Y (
         CALCULATOR_L5FirstOperands_1__5), .A0 (
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx554), .A1 (
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx558)) ;
    aoi22 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix555 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx554), .A0 (
          CALCULATOR_L4Results_0__4), .A1 (CALCULATOR_L3Results_2__4), .B0 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx48), .B1 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx12)) ;
    xnor2 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix559 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx558), .A0 (
          CALCULATOR_L3Results_2__5), .A1 (CALCULATOR_L4Results_0__5)) ;
    xor2 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix67 (.Y (
         CALCULATOR_L5FirstOperands_1__6), .A0 (
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx561), .A1 (
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx565)) ;
    aoi22 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix562 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx561), .A0 (
          CALCULATOR_L4Results_0__5), .A1 (CALCULATOR_L3Results_2__5), .B0 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx52), .B1 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx6)) ;
    xnor2 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix566 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx565), .A0 (
          CALCULATOR_L3Results_2__6), .A1 (CALCULATOR_L4Results_0__6)) ;
    xnor2 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix65 (.Y (
          CALCULATOR_L5FirstOperands_1__7), .A0 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx568), .A1 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx62)) ;
    aoi22 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix569 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx568), .A0 (
          CALCULATOR_L4Results_0__6), .A1 (CALCULATOR_L3Results_2__6), .B0 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx56), .B1 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx0)) ;
    xor2 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix63 (.Y (
         CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx62), .A0 (CALCULATOR_L3Results_2__7)
         , .A1 (CALCULATOR_L4Results_0__7)) ;
    inv01 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix155 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx154), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx383)) ;
    inv01 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix57 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx56), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx561)) ;
    inv01 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix53 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx52), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx554)) ;
    inv01 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix49 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx48), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx547)) ;
    inv01 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix45 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx44), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx540)) ;
    inv01 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix41 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx40), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx534)) ;
    inv01 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix31 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx30), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx531)) ;
    inv01 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix25 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx24), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx537)) ;
    inv01 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix19 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx18), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx544)) ;
    inv01 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix13 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx12), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx551)) ;
    inv01 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix7 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx6), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx558)) ;
    inv01 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix1 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx0), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx565)) ;
    fake_gnd CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix216 (.Y (
             CALCULATOR_L1_4_L2_3_G5_MINI_ALU_WindowCellShiftedLeft_16)) ;
    aoi21 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix77 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_10), .A0 (
          CacheFilter_4__3__1), .A1 (CacheFilter_4__3__0), .B0 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_nx4)) ;
    nor02_2x CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix5 (.Y (
             CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_nx4), .A0 (
             CacheFilter_4__3__0), .A1 (CacheFilter_4__3__1)) ;
    aoi21 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix67 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_11), .A0 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_nx328), .A1 (
          CacheFilter_4__3__2), .B0 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_nx8)) ;
    nor03_2x CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix9 (.Y (
             CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_nx8), .A0 (
             CacheFilter_4__3__2), .A1 (CacheFilter_4__3__0), .A2 (
             CacheFilter_4__3__1)) ;
    xnor2 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix59 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_12), .A0 (
          CacheFilter_4__3__3), .A1 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_nx8)) ;
    xnor2 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix51 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_13), .A0 (
          CacheFilter_4__3__4), .A1 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_nx12)) ;
    nor04 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix13 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_nx12), .A0 (
          CacheFilter_4__3__3), .A1 (CacheFilter_4__3__2), .A2 (
          CacheFilter_4__3__0), .A3 (CacheFilter_4__3__1)) ;
    xnor2 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix43 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_14), .A0 (
          CacheFilter_4__3__5), .A1 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_nx16)) ;
    nor02ii CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix17 (.Y (
            CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_nx16), .A0 (
            CacheFilter_4__3__4), .A1 (
            CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_nx12)) ;
    xnor2 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix35 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_15), .A0 (
          CacheFilter_4__3__6), .A1 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_nx20)) ;
    nor02ii CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix21 (.Y (
            CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_nx20), .A0 (
            CacheFilter_4__3__5), .A1 (
            CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_nx16)) ;
    xnor2 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix27 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_16), .A0 (
          CacheFilter_4__3__7), .A1 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_nx24)) ;
    nor02ii CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix25 (.Y (
            CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_nx24), .A0 (
            CacheFilter_4__3__6), .A1 (
            CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_nx20)) ;
    inv01 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix329 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_nx328), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_nx4)) ;
    inv02 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix383 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_nx384), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_0)) ;
    dff CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_0 (.Q (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_0), .QB (
        \$dummy [1200]), .D (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .CLK (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    nor02_2x CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix567 (.Y (
             CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566), .A0 (
             RST), .A1 (
             CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644)) ;
    dff CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_1 (.Q (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_1), .QB (
        \$dummy [1201]), .D (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .CLK (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_2 (.Q (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_2), .QB (
        \$dummy [1202]), .D (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .CLK (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_3 (.Q (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_3), .QB (
        \$dummy [1203]), .D (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .CLK (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_4 (.Q (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_4), .QB (
        \$dummy [1204]), .D (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .CLK (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_5 (.Q (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_5), .QB (
        \$dummy [1205]), .D (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .CLK (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_6 (.Q (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_6), .QB (
        \$dummy [1206]), .D (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .CLK (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_7 (.Q (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_7), .QB (
        \$dummy [1207]), .D (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .CLK (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_8 (.Q (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_8), .QB (
        \$dummy [1208]), .D (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .CLK (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_9 (.Q (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_9), .QB (
        \$dummy [1209]), .D (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .CLK (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_10 (.Q (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_10), .QB (
        \$dummy [1210]), .D (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .CLK (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_11 (.Q (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_11), .QB (
        \$dummy [1211]), .D (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .CLK (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_12 (.Q (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_12), .QB (
        \$dummy [1212]), .D (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .CLK (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_13 (.Q (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_13), .QB (
        \$dummy [1213]), .D (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .CLK (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_14 (.Q (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_14), .QB (
        \$dummy [1214]), .D (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .CLK (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_15 (.Q (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_15), .QB (
        \$dummy [1215]), .D (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .CLK (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_16 (.Q (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_16), .QB (
        \$dummy [1216]), .D (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .CLK (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    inv02 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix623 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix625 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix627 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix643 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644), .A (
          nx8299)) ;
    dff CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_0 (.Q (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_0), .QB (
        \$dummy [1217]), .D (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .CLK (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    nor02_2x CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix567 (.Y (
             CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566), .A0 (
             RST), .A1 (
             CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644)) ;
    dff CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_1 (.Q (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_1), .QB (
        \$dummy [1218]), .D (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .CLK (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_2 (.Q (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_2), .QB (
        \$dummy [1219]), .D (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .CLK (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_3 (.Q (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_3), .QB (
        \$dummy [1220]), .D (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .CLK (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_4 (.Q (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_4), .QB (
        \$dummy [1221]), .D (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .CLK (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_5 (.Q (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_5), .QB (
        \$dummy [1222]), .D (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .CLK (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_6 (.Q (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_6), .QB (
        \$dummy [1223]), .D (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .CLK (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_7 (.Q (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_7), .QB (
        \$dummy [1224]), .D (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .CLK (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_8 (.Q (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_8), .QB (
        \$dummy [1225]), .D (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .CLK (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_9 (.Q (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_9), .QB (
        \$dummy [1226]), .D (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .CLK (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_10 (.Q (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_10), .QB (
        \$dummy [1227]), .D (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .CLK (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_11 (.Q (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_11), .QB (
        \$dummy [1228]), .D (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .CLK (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_12 (.Q (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_12), .QB (
        \$dummy [1229]), .D (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .CLK (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_13 (.Q (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_13), .QB (
        \$dummy [1230]), .D (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .CLK (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_14 (.Q (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_14), .QB (
        \$dummy [1231]), .D (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .CLK (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_15 (.Q (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_15), .QB (
        \$dummy [1232]), .D (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .CLK (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_16 (.Q (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_16), .QB (
        \$dummy [1233]), .D (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .CLK (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    inv02 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix623 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix625 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix627 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix643 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644), .A (
          nx8305)) ;
    dff CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_0 (.Q (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_0), .QB (\$dummy [1234]), .D (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .CLK (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    nor02_2x CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix567 (.Y (
             CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566), .A0 (
             RST), .A1 (
             CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    dff CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_1 (.Q (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_1), .QB (\$dummy [1235]), .D (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .CLK (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_2 (.Q (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_2), .QB (\$dummy [1236]), .D (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .CLK (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_3 (.Q (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_3), .QB (\$dummy [1237]), .D (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .CLK (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_4 (.Q (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_4), .QB (\$dummy [1238]), .D (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .CLK (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_5 (.Q (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_5), .QB (\$dummy [1239]), .D (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .CLK (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_6 (.Q (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_6), .QB (\$dummy [1240]), .D (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .CLK (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_7 (.Q (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_7), .QB (\$dummy [1241]), .D (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .CLK (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_8 (.Q (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_8), .QB (\$dummy [1242]), .D (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .CLK (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_9 (.Q (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_9), .QB (\$dummy [1243]), .D (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .CLK (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_10 (.Q (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_10), .QB (\$dummy [1244]), .D (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .CLK (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_11 (.Q (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_11), .QB (\$dummy [1245]), .D (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .CLK (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_12 (.Q (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_12), .QB (\$dummy [1246]), .D (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .CLK (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_13 (.Q (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_13), .QB (\$dummy [1247]), .D (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .CLK (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_14 (.Q (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_14), .QB (\$dummy [1248]), .D (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .CLK (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_15 (.Q (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_15), .QB (\$dummy [1249]), .D (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .CLK (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_16 (.Q (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_16), .QB (\$dummy [1250]), .D (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .CLK (
        CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    inv02 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix623 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix625 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix627 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix643 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642)) ;
    xor2 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix83 (.Y (CALCULATOR_L5Results_1__0), 
         .A0 (CALCULATOR_L5SecondOperands_1__0), .A1 (
         CALCULATOR_L5FirstOperands_1__0)) ;
    xnor2 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix380 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx379), .A0 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx381), .A1 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx383)) ;
    nand02 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix382 (.Y (
           CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx381), .A0 (
           CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothOperand_0), .A1 (nx8325)) ;
    xnor2 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix384 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx383), .A0 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothOperand_1), .A1 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_1)) ;
    inv01 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix388 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx387), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_2)) ;
    xnor2 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix390 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx389), .A0 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx391), .A1 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx395)) ;
    aoi32 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix392 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx391), .A0 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothOperand_0), .A1 (nx8325), .A2 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx154), .B0 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_1), .B1 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothOperand_1)) ;
    xnor2 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix396 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx395), .A0 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothOperand_2), .A1 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_2)) ;
    inv01 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix400 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx399), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_3)) ;
    xnor2 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix402 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx401), .A0 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx403), .A1 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx405)) ;
    xnor2 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix406 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx405), .A0 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothOperand_3), .A1 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_3)) ;
    inv01 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix410 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx409), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_4)) ;
    xnor2 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix412 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx411), .A0 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx413), .A1 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx415)) ;
    xnor2 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix416 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx415), .A0 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothOperand_4), .A1 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_4)) ;
    inv01 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix420 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx419), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_5)) ;
    xnor2 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix422 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx421), .A0 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx423), .A1 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx425)) ;
    xnor2 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix426 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx425), .A0 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothOperand_5), .A1 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_5)) ;
    inv01 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix430 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx429), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_6)) ;
    xnor2 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix432 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx431), .A0 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx433), .A1 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx435)) ;
    xnor2 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix436 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx435), .A0 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothOperand_6), .A1 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_6)) ;
    inv01 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix440 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx439), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_7)) ;
    xnor2 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix442 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx441), .A0 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx443), .A1 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx445)) ;
    xnor2 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix446 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx445), .A0 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothOperand_7), .A1 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_7)) ;
    inv01 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix450 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx449), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_8)) ;
    xnor2 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix452 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx451), .A0 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx453), .A1 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx455)) ;
    xnor2 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix456 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx455), .A0 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothOperand_8), .A1 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_8)) ;
    xor2 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix317 (.Y (
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx316), .A0 (
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx461), .A1 (
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx463)) ;
    xnor2 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix464 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx463), .A0 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothOperand_9), .A1 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_9)) ;
    xor2 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix337 (.Y (
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx336), .A0 (
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx467), .A1 (
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx471)) ;
    inv01 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix470 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx469), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_9)) ;
    xnor2 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix472 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx471), .A0 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothOperand_10), .A1 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_10)) ;
    xor2 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix357 (.Y (
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx356), .A0 (
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx475), .A1 (
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx479)) ;
    inv01 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix478 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx477), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_10)) ;
    xnor2 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix480 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx479), .A0 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothOperand_11), .A1 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_11)) ;
    xor2 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix377 (.Y (
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx376), .A0 (
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx483), .A1 (
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx487)) ;
    inv01 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix486 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx485), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_11)) ;
    xnor2 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix488 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx487), .A0 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothOperand_12), .A1 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_12)) ;
    xor2 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix397 (.Y (
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx396), .A0 (
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx491), .A1 (
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx495)) ;
    inv01 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix494 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx493), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_12)) ;
    xnor2 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix496 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx495), .A0 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothOperand_13), .A1 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_13)) ;
    xor2 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix417 (.Y (
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx416), .A0 (
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx499), .A1 (
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx503)) ;
    inv01 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix502 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx501), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_13)) ;
    xnor2 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix504 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx503), .A0 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothOperand_14), .A1 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_14)) ;
    xor2 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix437 (.Y (
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx436), .A0 (
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx507), .A1 (
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx511)) ;
    inv01 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix510 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx509), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_14)) ;
    xnor2 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix512 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx511), .A0 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothOperand_15), .A1 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_15)) ;
    xnor2 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix457 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx456), .A0 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx515), .A1 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx454)) ;
    inv01 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix518 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx517), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_15)) ;
    xor2 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix455 (.Y (
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx454), .A0 (
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothOperand_16), .A1 (
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_16)) ;
    mux21_ni CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix91 (.Y (
             CALCULATOR_L5SecondOperands_1__0), .A0 (
             CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_1), .A1 (
             CacheWindow_4__4__0), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix99 (.Y (
             CALCULATOR_L5SecondOperands_1__1), .A0 (
             CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_2), .A1 (
             CacheWindow_4__4__1), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix107 (.Y (
             CALCULATOR_L5SecondOperands_1__2), .A0 (
             CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_3), .A1 (
             CacheWindow_4__4__2), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix115 (.Y (
             CALCULATOR_L5SecondOperands_1__3), .A0 (
             CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_4), .A1 (
             CacheWindow_4__4__3), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix123 (.Y (
             CALCULATOR_L5SecondOperands_1__4), .A0 (
             CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_5), .A1 (
             CacheWindow_4__4__4), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix131 (.Y (
             CALCULATOR_L5SecondOperands_1__5), .A0 (
             CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_6), .A1 (
             CacheWindow_4__4__5), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix139 (.Y (
             CALCULATOR_L5SecondOperands_1__6), .A0 (
             CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_7), .A1 (
             CacheWindow_4__4__6), .S0 (Instr)) ;
    mux21_ni CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix147 (.Y (
             CALCULATOR_L5SecondOperands_1__7), .A0 (
             CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_8), .A1 (
             CacheWindow_4__4__7), .S0 (Instr)) ;
    xor2 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix77 (.Y (CALCULATOR_L5Results_1__1), 
         .A0 (CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx529), .A1 (
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx531)) ;
    nand02 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix530 (.Y (
           CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx529), .A0 (
           CALCULATOR_L5SecondOperands_1__0), .A1 (
           CALCULATOR_L5FirstOperands_1__0)) ;
    xnor2 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix532 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx531), .A0 (
          CALCULATOR_L5SecondOperands_1__1), .A1 (
          CALCULATOR_L5FirstOperands_1__1)) ;
    xor2 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix75 (.Y (CALCULATOR_L5Results_1__2), 
         .A0 (CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx534), .A1 (
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx537)) ;
    aoi32 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix535 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx534), .A0 (
          CALCULATOR_L5SecondOperands_1__0), .A1 (
          CALCULATOR_L5FirstOperands_1__0), .A2 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx30), .B0 (
          CALCULATOR_L5FirstOperands_1__1), .B1 (
          CALCULATOR_L5SecondOperands_1__1)) ;
    xnor2 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix538 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx537), .A0 (
          CALCULATOR_L5SecondOperands_1__2), .A1 (
          CALCULATOR_L5FirstOperands_1__2)) ;
    xor2 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix73 (.Y (CALCULATOR_L5Results_1__3), 
         .A0 (CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx540), .A1 (
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx544)) ;
    aoi22 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix541 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx540), .A0 (
          CALCULATOR_L5FirstOperands_1__2), .A1 (
          CALCULATOR_L5SecondOperands_1__2), .B0 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx40), .B1 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx24)) ;
    xnor2 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix545 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx544), .A0 (
          CALCULATOR_L5SecondOperands_1__3), .A1 (
          CALCULATOR_L5FirstOperands_1__3)) ;
    xor2 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix71 (.Y (CALCULATOR_L5Results_1__4), 
         .A0 (CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx547), .A1 (
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx551)) ;
    aoi22 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix548 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx547), .A0 (
          CALCULATOR_L5FirstOperands_1__3), .A1 (
          CALCULATOR_L5SecondOperands_1__3), .B0 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx44), .B1 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx18)) ;
    xnor2 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix552 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx551), .A0 (
          CALCULATOR_L5SecondOperands_1__4), .A1 (
          CALCULATOR_L5FirstOperands_1__4)) ;
    xor2 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix69 (.Y (CALCULATOR_L5Results_1__5), 
         .A0 (CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx554), .A1 (
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx558)) ;
    aoi22 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix555 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx554), .A0 (
          CALCULATOR_L5FirstOperands_1__4), .A1 (
          CALCULATOR_L5SecondOperands_1__4), .B0 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx48), .B1 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx12)) ;
    xnor2 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix559 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx558), .A0 (
          CALCULATOR_L5SecondOperands_1__5), .A1 (
          CALCULATOR_L5FirstOperands_1__5)) ;
    xor2 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix67 (.Y (CALCULATOR_L5Results_1__6), 
         .A0 (CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx561), .A1 (
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx565)) ;
    aoi22 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix562 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx561), .A0 (
          CALCULATOR_L5FirstOperands_1__5), .A1 (
          CALCULATOR_L5SecondOperands_1__5), .B0 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx52), .B1 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx6)) ;
    xnor2 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix566 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx565), .A0 (
          CALCULATOR_L5SecondOperands_1__6), .A1 (
          CALCULATOR_L5FirstOperands_1__6)) ;
    xnor2 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix65 (.Y (CALCULATOR_L5Results_1__7)
          , .A0 (CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx568), .A1 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx62)) ;
    aoi22 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix569 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx568), .A0 (
          CALCULATOR_L5FirstOperands_1__6), .A1 (
          CALCULATOR_L5SecondOperands_1__6), .B0 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx56), .B1 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx0)) ;
    xor2 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix63 (.Y (
         CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx62), .A0 (
         CALCULATOR_L5SecondOperands_1__7), .A1 (CALCULATOR_L5FirstOperands_1__7
         )) ;
    inv01 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix155 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx154), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx383)) ;
    inv01 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix57 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx56), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx561)) ;
    inv01 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix53 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx52), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx554)) ;
    inv01 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix49 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx48), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx547)) ;
    inv01 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix45 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx44), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx540)) ;
    inv01 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix41 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx40), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx534)) ;
    inv01 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix31 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx30), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx531)) ;
    inv01 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix25 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx24), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx537)) ;
    inv01 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix19 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx18), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx544)) ;
    inv01 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix13 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx12), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx551)) ;
    inv01 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix7 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx6), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx558)) ;
    inv01 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix1 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx0), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx565)) ;
    fake_gnd CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix216 (.Y (
             CALCULATOR_L1_4_L2_4_G5_MINI_ALU_WindowCellShiftedLeft_16)) ;
    aoi21 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix77 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_10), .A0 (
          CacheFilter_4__4__1), .A1 (CacheFilter_4__4__0), .B0 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_nx4)) ;
    nor02_2x CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix5 (.Y (
             CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_nx4), .A0 (
             CacheFilter_4__4__0), .A1 (CacheFilter_4__4__1)) ;
    aoi21 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix67 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_11), .A0 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_nx328), .A1 (
          CacheFilter_4__4__2), .B0 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_nx8)) ;
    nor03_2x CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix9 (.Y (
             CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_nx8), .A0 (
             CacheFilter_4__4__2), .A1 (CacheFilter_4__4__0), .A2 (
             CacheFilter_4__4__1)) ;
    xnor2 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix59 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_12), .A0 (
          CacheFilter_4__4__3), .A1 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_nx8)) ;
    xnor2 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix51 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_13), .A0 (
          CacheFilter_4__4__4), .A1 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_nx12)) ;
    nor04 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix13 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_nx12), .A0 (
          CacheFilter_4__4__3), .A1 (CacheFilter_4__4__2), .A2 (
          CacheFilter_4__4__0), .A3 (CacheFilter_4__4__1)) ;
    xnor2 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix43 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_14), .A0 (
          CacheFilter_4__4__5), .A1 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_nx16)) ;
    nor02ii CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix17 (.Y (
            CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_nx16), .A0 (
            CacheFilter_4__4__4), .A1 (
            CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_nx12)) ;
    xnor2 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix35 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_15), .A0 (
          CacheFilter_4__4__6), .A1 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_nx20)) ;
    nor02ii CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix21 (.Y (
            CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_nx20), .A0 (
            CacheFilter_4__4__5), .A1 (
            CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_nx16)) ;
    xnor2 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix27 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_16), .A0 (
          CacheFilter_4__4__7), .A1 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_nx24)) ;
    nor02ii CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix25 (.Y (
            CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_nx24), .A0 (
            CacheFilter_4__4__6), .A1 (
            CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_nx20)) ;
    inv01 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix329 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_nx328), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_nx4)) ;
    inv02 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix383 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_nx384), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_0)) ;
    dff CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_0 (.Q (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_0), .QB (
        \$dummy [1251]), .D (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .CLK (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    nor02_2x CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix567 (.Y (
             CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566), .A0 (
             RST), .A1 (
             CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644)) ;
    dff CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_1 (.Q (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_1), .QB (
        \$dummy [1252]), .D (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .CLK (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_2 (.Q (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_2), .QB (
        \$dummy [1253]), .D (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .CLK (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_3 (.Q (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_3), .QB (
        \$dummy [1254]), .D (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .CLK (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_4 (.Q (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_4), .QB (
        \$dummy [1255]), .D (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .CLK (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_5 (.Q (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_5), .QB (
        \$dummy [1256]), .D (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .CLK (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_6 (.Q (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_6), .QB (
        \$dummy [1257]), .D (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .CLK (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_7 (.Q (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_7), .QB (
        \$dummy [1258]), .D (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .CLK (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_8 (.Q (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_8), .QB (
        \$dummy [1259]), .D (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .CLK (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_9 (.Q (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_9), .QB (
        \$dummy [1260]), .D (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .CLK (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_10 (.Q (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_10), .QB (
        \$dummy [1261]), .D (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .CLK (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_11 (.Q (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_11), .QB (
        \$dummy [1262]), .D (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .CLK (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_12 (.Q (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_12), .QB (
        \$dummy [1263]), .D (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .CLK (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_13 (.Q (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_13), .QB (
        \$dummy [1264]), .D (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .CLK (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_14 (.Q (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_14), .QB (
        \$dummy [1265]), .D (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .CLK (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_15 (.Q (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_15), .QB (
        \$dummy [1266]), .D (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .CLK (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_16 (.Q (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_16), .QB (
        \$dummy [1267]), .D (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .CLK (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    inv02 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix623 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix625 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix627 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix643 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644), .A (
          nx8339)) ;
    dff CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_0 (.Q (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_0), .QB (
        \$dummy [1268]), .D (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .CLK (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    nor02_2x CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix567 (.Y (
             CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566), .A0 (
             RST), .A1 (
             CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644)) ;
    dff CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_1 (.Q (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_1), .QB (
        \$dummy [1269]), .D (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .CLK (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_2 (.Q (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_2), .QB (
        \$dummy [1270]), .D (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .CLK (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_3 (.Q (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_3), .QB (
        \$dummy [1271]), .D (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .CLK (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_4 (.Q (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_4), .QB (
        \$dummy [1272]), .D (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .CLK (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_5 (.Q (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_5), .QB (
        \$dummy [1273]), .D (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .CLK (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_6 (.Q (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_6), .QB (
        \$dummy [1274]), .D (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .CLK (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_7 (.Q (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_7), .QB (
        \$dummy [1275]), .D (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .CLK (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_8 (.Q (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_8), .QB (
        \$dummy [1276]), .D (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .CLK (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_9 (.Q (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_9), .QB (
        \$dummy [1277]), .D (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .CLK (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_10 (.Q (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_10), .QB (
        \$dummy [1278]), .D (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .CLK (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_11 (.Q (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_11), .QB (
        \$dummy [1279]), .D (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .CLK (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_12 (.Q (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_12), .QB (
        \$dummy [1280]), .D (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .CLK (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_13 (.Q (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_13), .QB (
        \$dummy [1281]), .D (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .CLK (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_14 (.Q (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_14), .QB (
        \$dummy [1282]), .D (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .CLK (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_15 (.Q (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_15), .QB (
        \$dummy [1283]), .D (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .CLK (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_16 (.Q (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_16), .QB (
        \$dummy [1284]), .D (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .CLK (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    inv02 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix623 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix625 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix627 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix643 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644), .A (
          nx8345)) ;
    dff CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_0 (.Q (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_0), .QB (\$dummy [1285]), .D (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .CLK (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    nor02_2x CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix567 (.Y (
             CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566), .A0 (
             RST), .A1 (
             CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    dff CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_1 (.Q (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_1), .QB (\$dummy [1286]), .D (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .CLK (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_2 (.Q (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_2), .QB (\$dummy [1287]), .D (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .CLK (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_3 (.Q (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_3), .QB (\$dummy [1288]), .D (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .CLK (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_4 (.Q (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_4), .QB (\$dummy [1289]), .D (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .CLK (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_5 (.Q (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_5), .QB (\$dummy [1290]), .D (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .CLK (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_6 (.Q (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_6), .QB (\$dummy [1291]), .D (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .CLK (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_7 (.Q (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_7), .QB (\$dummy [1292]), .D (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .CLK (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_8 (.Q (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_8), .QB (\$dummy [1293]), .D (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .CLK (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_9 (.Q (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_9), .QB (\$dummy [1294]), .D (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .CLK (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_10 (.Q (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_10), .QB (\$dummy [1295]), .D (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .CLK (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_11 (.Q (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_11), .QB (\$dummy [1296]), .D (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .CLK (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_12 (.Q (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_12), .QB (\$dummy [1297]), .D (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .CLK (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_13 (.Q (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_13), .QB (\$dummy [1298]), .D (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .CLK (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_14 (.Q (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_14), .QB (\$dummy [1299]), .D (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .CLK (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_15 (.Q (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_15), .QB (\$dummy [1300]), .D (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .CLK (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_16 (.Q (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_16), .QB (\$dummy [1301]), .D (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .CLK (
        CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    inv02 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix623 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix625 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix627 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628), .A (CLK
          )) ;
    inv02 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix643 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642)) ;
    inv01 CACHE_ix942 (.Y (CACHE_EN_dup_1491), .A (CACHE_nx941)) ;
    inv01 CACHE_ix944 (.Y (CACHE_EN_dup_1359), .A (CACHE_nx941)) ;
    inv01 CACHE_ix946 (.Y (CACHE_EN_dup_1227), .A (CACHE_nx941)) ;
    inv01 CACHE_ix948 (.Y (CACHE_EN_dup_1161), .A (CACHE_nx941)) ;
    inv01 CACHE_ix950 (.Y (CACHE_EN_dup_1095), .A (CACHE_nx941)) ;
    inv01 CACHE_ix952 (.Y (CACHE_EN), .A (CACHE_nx941)) ;
    inv01 CACHE_ix956 (.Y (CACHE_EN_dup_1502), .A (CACHE_nx955)) ;
    inv01 CACHE_ix958 (.Y (CACHE_EN_dup_1370), .A (CACHE_nx955)) ;
    inv01 CACHE_ix960 (.Y (CACHE_EN_dup_1238), .A (CACHE_nx955)) ;
    inv01 CACHE_ix962 (.Y (CACHE_EN_dup_1172), .A (CACHE_nx955)) ;
    inv01 CACHE_ix964 (.Y (CACHE_EN_dup_1106), .A (CACHE_nx955)) ;
    inv01 CACHE_ix966 (.Y (CACHE_EN_dup_1084), .A (CACHE_nx955)) ;
    inv02 CACHE_ix974 (.Y (CACHE_RST_dup_1073), .A (nx8457)) ;
    inv02 CACHE_ix976 (.Y (CACHE_RST_dup_1094), .A (nx8457)) ;
    inv02 CACHE_ix978 (.Y (CACHE_RST_dup_1116), .A (nx8457)) ;
    inv02 CACHE_ix980 (.Y (CACHE_RST_dup_1138), .A (nx8457)) ;
    inv02 CACHE_ix982 (.Y (CACHE_RST_dup_1160), .A (nx8457)) ;
    inv02 CACHE_ix984 (.Y (CACHE_RST_dup_1182), .A (nx8457)) ;
    inv02 CACHE_ix986 (.Y (CACHE_RST_dup_1204), .A (nx8457)) ;
    inv02 CACHE_ix988 (.Y (CACHE_RST_dup_1226), .A (nx8461)) ;
    inv02 CACHE_ix990 (.Y (CACHE_RST_dup_1248), .A (nx8461)) ;
    inv02 CACHE_ix992 (.Y (CACHE_RST_dup_1270), .A (nx8461)) ;
    inv02 CACHE_ix994 (.Y (CACHE_RST_dup_1292), .A (nx8461)) ;
    inv02 CACHE_ix996 (.Y (CACHE_RST_dup_1314), .A (nx8461)) ;
    inv02 CACHE_ix998 (.Y (CACHE_RST_dup_1336), .A (nx8461)) ;
    inv02 CACHE_ix1000 (.Y (CACHE_RST_dup_1358), .A (nx8461)) ;
    inv02 CACHE_ix1002 (.Y (CACHE_RST_dup_1380), .A (nx8465)) ;
    inv02 CACHE_ix1004 (.Y (CACHE_RST_dup_1402), .A (nx8465)) ;
    inv02 CACHE_ix1006 (.Y (CACHE_RST_dup_1424), .A (nx8465)) ;
    inv02 CACHE_ix1008 (.Y (CACHE_RST_dup_1446), .A (nx8465)) ;
    inv02 CACHE_ix1010 (.Y (CACHE_RST_dup_1468), .A (nx8465)) ;
    inv02 CACHE_ix1012 (.Y (CACHE_RST_dup_1490), .A (nx8465)) ;
    inv02 CACHE_ix1014 (.Y (CACHE_RST_dup_1512), .A (nx8465)) ;
    inv02 CACHE_ix1016 (.Y (CACHE_RST_dup_1534), .A (nx8469)) ;
    inv02 CACHE_ix1018 (.Y (CACHE_RST_dup_1556), .A (nx8469)) ;
    inv02 CACHE_ix1020 (.Y (CACHE_RST_dup_1578), .A (nx8469)) ;
    inv02 CACHE_ix1022 (.Y (CACHE_RST_dup_1600), .A (nx8469)) ;
    inv01 CACHE_ix1024 (.Y (CACHE_nx1025), .A (CacheFilterWR)) ;
    inv01 CACHE_ix1026 (.Y (CACHE_EN_dup_1293), .A (CACHE_nx1025)) ;
    inv01 CACHE_ix1028 (.Y (CACHE_EN_dup_1403), .A (CACHE_nx1025)) ;
    inv01 CACHE_ix1030 (.Y (CACHE_EN_dup_1513), .A (CACHE_nx1025)) ;
    inv01 CACHE_ix1032 (.Y (CACHE_nx1033), .A (CacheWindowWR)) ;
    inv01 CACHE_ix1034 (.Y (CACHE_EN_dup_1304), .A (CACHE_nx1033)) ;
    inv01 CACHE_ix1036 (.Y (CACHE_EN_dup_1414), .A (CACHE_nx1033)) ;
    inv01 CACHE_ix1038 (.Y (CACHE_EN_dup_1524), .A (CACHE_nx1033)) ;
    inv02 CACHE_ix1040 (.Y (CACHE_nx1041), .A (CacheRST)) ;
    inv02 CACHE_ix1042 (.Y (CACHE_nx1043), .A (nx8833)) ;
    inv02 CACHE_ix1044 (.Y (CACHE_nx1045), .A (nx8833)) ;
    inv02 CACHE_ix1046 (.Y (CACHE_nx1047), .A (nx8833)) ;
    dff CACHE_L0_0_L1_0_Fij_reg_Dout_0 (.Q (CacheFilter_0__0__0), .QB (
        \$dummy [1302]), .D (CACHE_L0_0_L1_0_Fij_nx212), .CLK (CLK)) ;
    nor02_2x CACHE_L0_0_L1_0_Fij_ix297 (.Y (CACHE_L0_0_L1_0_Fij_nx296), .A0 (
             nx8357), .A1 (CACHE_L0_0_L1_0_Fij_nx331)) ;
    dff CACHE_L0_0_L1_0_Fij_reg_Dout_1 (.Q (CacheFilter_0__0__1), .QB (
        \$dummy [1303]), .D (CACHE_L0_0_L1_0_Fij_nx222), .CLK (CLK)) ;
    dff CACHE_L0_0_L1_0_Fij_reg_Dout_2 (.Q (CacheFilter_0__0__2), .QB (
        \$dummy [1304]), .D (CACHE_L0_0_L1_0_Fij_nx232), .CLK (CLK)) ;
    dff CACHE_L0_0_L1_0_Fij_reg_Dout_3 (.Q (CacheFilter_0__0__3), .QB (
        \$dummy [1305]), .D (CACHE_L0_0_L1_0_Fij_nx242), .CLK (CLK)) ;
    dff CACHE_L0_0_L1_0_Fij_reg_Dout_4 (.Q (CacheFilter_0__0__4), .QB (
        \$dummy [1306]), .D (CACHE_L0_0_L1_0_Fij_nx252), .CLK (CLK)) ;
    dff CACHE_L0_0_L1_0_Fij_reg_Dout_5 (.Q (CacheFilter_0__0__5), .QB (
        \$dummy [1307]), .D (CACHE_L0_0_L1_0_Fij_nx262), .CLK (CLK)) ;
    dff CACHE_L0_0_L1_0_Fij_reg_Dout_6 (.Q (CacheFilter_0__0__6), .QB (
        \$dummy [1308]), .D (CACHE_L0_0_L1_0_Fij_nx272), .CLK (CLK)) ;
    dff CACHE_L0_0_L1_0_Fij_reg_Dout_7 (.Q (CacheFilter_0__0__7), .QB (
        \$dummy [1309]), .D (CACHE_L0_0_L1_0_Fij_nx282), .CLK (CLK)) ;
    buf02 CACHE_L0_0_L1_0_Fij_ix330 (.Y (CACHE_L0_0_L1_0_Fij_nx331), .A (
          CACHE_EN)) ;
    buf02 CACHE_L0_0_L1_0_Fij_ix332 (.Y (CACHE_L0_0_L1_0_Fij_nx333), .A (
          CACHE_EN)) ;
    dff CACHE_L0_0_L1_0_Wij_reg_Dout_0 (.Q (CacheWindow_0__0__0), .QB (
        \$dummy [1310]), .D (CACHE_L0_0_L1_0_Wij_nx212), .CLK (CLK)) ;
    nor02_2x CACHE_L0_0_L1_0_Wij_ix297 (.Y (CACHE_L0_0_L1_0_Wij_nx296), .A0 (
             nx8357), .A1 (CACHE_L0_0_L1_0_Wij_nx331)) ;
    dff CACHE_L0_0_L1_0_Wij_reg_Dout_1 (.Q (CacheWindow_0__0__1), .QB (
        \$dummy [1311]), .D (CACHE_L0_0_L1_0_Wij_nx222), .CLK (CLK)) ;
    dff CACHE_L0_0_L1_0_Wij_reg_Dout_2 (.Q (CacheWindow_0__0__2), .QB (
        \$dummy [1312]), .D (CACHE_L0_0_L1_0_Wij_nx232), .CLK (CLK)) ;
    dff CACHE_L0_0_L1_0_Wij_reg_Dout_3 (.Q (CacheWindow_0__0__3), .QB (
        \$dummy [1313]), .D (CACHE_L0_0_L1_0_Wij_nx242), .CLK (CLK)) ;
    dff CACHE_L0_0_L1_0_Wij_reg_Dout_4 (.Q (CacheWindow_0__0__4), .QB (
        \$dummy [1314]), .D (CACHE_L0_0_L1_0_Wij_nx252), .CLK (CLK)) ;
    dff CACHE_L0_0_L1_0_Wij_reg_Dout_5 (.Q (CacheWindow_0__0__5), .QB (
        \$dummy [1315]), .D (CACHE_L0_0_L1_0_Wij_nx262), .CLK (CLK)) ;
    dff CACHE_L0_0_L1_0_Wij_reg_Dout_6 (.Q (CacheWindow_0__0__6), .QB (
        \$dummy [1316]), .D (CACHE_L0_0_L1_0_Wij_nx272), .CLK (CLK)) ;
    dff CACHE_L0_0_L1_0_Wij_reg_Dout_7 (.Q (CacheWindow_0__0__7), .QB (
        \$dummy [1317]), .D (CACHE_L0_0_L1_0_Wij_nx282), .CLK (CLK)) ;
    buf02 CACHE_L0_0_L1_0_Wij_ix330 (.Y (CACHE_L0_0_L1_0_Wij_nx331), .A (
          CACHE_EN_dup_1084)) ;
    buf02 CACHE_L0_0_L1_0_Wij_ix332 (.Y (CACHE_L0_0_L1_0_Wij_nx333), .A (
          CACHE_EN_dup_1084)) ;
    dff CACHE_L0_0_L1_1_Fij_reg_Dout_0 (.Q (CacheFilter_0__1__0), .QB (
        \$dummy [1318]), .D (CACHE_L0_0_L1_1_Fij_nx212), .CLK (CLK)) ;
    nor02_2x CACHE_L0_0_L1_1_Fij_ix297 (.Y (CACHE_L0_0_L1_1_Fij_nx296), .A0 (
             nx8361), .A1 (CACHE_L0_0_L1_1_Fij_nx331)) ;
    dff CACHE_L0_0_L1_1_Fij_reg_Dout_1 (.Q (CacheFilter_0__1__1), .QB (
        \$dummy [1319]), .D (CACHE_L0_0_L1_1_Fij_nx222), .CLK (CLK)) ;
    dff CACHE_L0_0_L1_1_Fij_reg_Dout_2 (.Q (CacheFilter_0__1__2), .QB (
        \$dummy [1320]), .D (CACHE_L0_0_L1_1_Fij_nx232), .CLK (CLK)) ;
    dff CACHE_L0_0_L1_1_Fij_reg_Dout_3 (.Q (CacheFilter_0__1__3), .QB (
        \$dummy [1321]), .D (CACHE_L0_0_L1_1_Fij_nx242), .CLK (CLK)) ;
    dff CACHE_L0_0_L1_1_Fij_reg_Dout_4 (.Q (CacheFilter_0__1__4), .QB (
        \$dummy [1322]), .D (CACHE_L0_0_L1_1_Fij_nx252), .CLK (CLK)) ;
    dff CACHE_L0_0_L1_1_Fij_reg_Dout_5 (.Q (CacheFilter_0__1__5), .QB (
        \$dummy [1323]), .D (CACHE_L0_0_L1_1_Fij_nx262), .CLK (CLK)) ;
    dff CACHE_L0_0_L1_1_Fij_reg_Dout_6 (.Q (CacheFilter_0__1__6), .QB (
        \$dummy [1324]), .D (CACHE_L0_0_L1_1_Fij_nx272), .CLK (CLK)) ;
    dff CACHE_L0_0_L1_1_Fij_reg_Dout_7 (.Q (CacheFilter_0__1__7), .QB (
        \$dummy [1325]), .D (CACHE_L0_0_L1_1_Fij_nx282), .CLK (CLK)) ;
    buf02 CACHE_L0_0_L1_1_Fij_ix330 (.Y (CACHE_L0_0_L1_1_Fij_nx331), .A (
          CACHE_EN_dup_1095)) ;
    buf02 CACHE_L0_0_L1_1_Fij_ix332 (.Y (CACHE_L0_0_L1_1_Fij_nx333), .A (
          CACHE_EN_dup_1095)) ;
    dff CACHE_L0_0_L1_1_Wij_reg_Dout_0 (.Q (CacheWindow_0__1__0), .QB (
        \$dummy [1326]), .D (CACHE_L0_0_L1_1_Wij_nx212), .CLK (CLK)) ;
    nor02_2x CACHE_L0_0_L1_1_Wij_ix297 (.Y (CACHE_L0_0_L1_1_Wij_nx296), .A0 (
             nx8361), .A1 (CACHE_L0_0_L1_1_Wij_nx331)) ;
    dff CACHE_L0_0_L1_1_Wij_reg_Dout_1 (.Q (CacheWindow_0__1__1), .QB (
        \$dummy [1327]), .D (CACHE_L0_0_L1_1_Wij_nx222), .CLK (CLK)) ;
    dff CACHE_L0_0_L1_1_Wij_reg_Dout_2 (.Q (CacheWindow_0__1__2), .QB (
        \$dummy [1328]), .D (CACHE_L0_0_L1_1_Wij_nx232), .CLK (CLK)) ;
    dff CACHE_L0_0_L1_1_Wij_reg_Dout_3 (.Q (CacheWindow_0__1__3), .QB (
        \$dummy [1329]), .D (CACHE_L0_0_L1_1_Wij_nx242), .CLK (CLK)) ;
    dff CACHE_L0_0_L1_1_Wij_reg_Dout_4 (.Q (CacheWindow_0__1__4), .QB (
        \$dummy [1330]), .D (CACHE_L0_0_L1_1_Wij_nx252), .CLK (CLK)) ;
    dff CACHE_L0_0_L1_1_Wij_reg_Dout_5 (.Q (CacheWindow_0__1__5), .QB (
        \$dummy [1331]), .D (CACHE_L0_0_L1_1_Wij_nx262), .CLK (CLK)) ;
    dff CACHE_L0_0_L1_1_Wij_reg_Dout_6 (.Q (CacheWindow_0__1__6), .QB (
        \$dummy [1332]), .D (CACHE_L0_0_L1_1_Wij_nx272), .CLK (CLK)) ;
    dff CACHE_L0_0_L1_1_Wij_reg_Dout_7 (.Q (CacheWindow_0__1__7), .QB (
        \$dummy [1333]), .D (CACHE_L0_0_L1_1_Wij_nx282), .CLK (CLK)) ;
    buf02 CACHE_L0_0_L1_1_Wij_ix330 (.Y (CACHE_L0_0_L1_1_Wij_nx331), .A (
          CACHE_EN_dup_1106)) ;
    buf02 CACHE_L0_0_L1_1_Wij_ix332 (.Y (CACHE_L0_0_L1_1_Wij_nx333), .A (
          CACHE_EN_dup_1106)) ;
    dff CACHE_L0_0_L1_2_Fij_reg_Dout_0 (.Q (CacheFilter_0__2__0), .QB (
        \$dummy [1334]), .D (CACHE_L0_0_L1_2_Fij_nx212), .CLK (CLK)) ;
    nor02_2x CACHE_L0_0_L1_2_Fij_ix297 (.Y (CACHE_L0_0_L1_2_Fij_nx296), .A0 (
             nx8365), .A1 (CACHE_L0_0_L1_2_Fij_nx331)) ;
    dff CACHE_L0_0_L1_2_Fij_reg_Dout_1 (.Q (CacheFilter_0__2__1), .QB (
        \$dummy [1335]), .D (CACHE_L0_0_L1_2_Fij_nx222), .CLK (CLK)) ;
    dff CACHE_L0_0_L1_2_Fij_reg_Dout_2 (.Q (CacheFilter_0__2__2), .QB (
        \$dummy [1336]), .D (CACHE_L0_0_L1_2_Fij_nx232), .CLK (CLK)) ;
    dff CACHE_L0_0_L1_2_Fij_reg_Dout_3 (.Q (CacheFilter_0__2__3), .QB (
        \$dummy [1337]), .D (CACHE_L0_0_L1_2_Fij_nx242), .CLK (CLK)) ;
    dff CACHE_L0_0_L1_2_Fij_reg_Dout_4 (.Q (CacheFilter_0__2__4), .QB (
        \$dummy [1338]), .D (CACHE_L0_0_L1_2_Fij_nx252), .CLK (CLK)) ;
    dff CACHE_L0_0_L1_2_Fij_reg_Dout_5 (.Q (CacheFilter_0__2__5), .QB (
        \$dummy [1339]), .D (CACHE_L0_0_L1_2_Fij_nx262), .CLK (CLK)) ;
    dff CACHE_L0_0_L1_2_Fij_reg_Dout_6 (.Q (CacheFilter_0__2__6), .QB (
        \$dummy [1340]), .D (CACHE_L0_0_L1_2_Fij_nx272), .CLK (CLK)) ;
    dff CACHE_L0_0_L1_2_Fij_reg_Dout_7 (.Q (CacheFilter_0__2__7), .QB (
        \$dummy [1341]), .D (CACHE_L0_0_L1_2_Fij_nx282), .CLK (CLK)) ;
    buf02 CACHE_L0_0_L1_2_Fij_ix330 (.Y (CACHE_L0_0_L1_2_Fij_nx331), .A (
          CACHE_EN_dup_1095)) ;
    buf02 CACHE_L0_0_L1_2_Fij_ix332 (.Y (CACHE_L0_0_L1_2_Fij_nx333), .A (
          CACHE_EN_dup_1095)) ;
    dff CACHE_L0_0_L1_2_Wij_reg_Dout_0 (.Q (CacheWindow_0__2__0), .QB (
        \$dummy [1342]), .D (CACHE_L0_0_L1_2_Wij_nx212), .CLK (CLK)) ;
    nor02_2x CACHE_L0_0_L1_2_Wij_ix297 (.Y (CACHE_L0_0_L1_2_Wij_nx296), .A0 (
             nx8365), .A1 (CACHE_L0_0_L1_2_Wij_nx331)) ;
    dff CACHE_L0_0_L1_2_Wij_reg_Dout_1 (.Q (CacheWindow_0__2__1), .QB (
        \$dummy [1343]), .D (CACHE_L0_0_L1_2_Wij_nx222), .CLK (CLK)) ;
    dff CACHE_L0_0_L1_2_Wij_reg_Dout_2 (.Q (CacheWindow_0__2__2), .QB (
        \$dummy [1344]), .D (CACHE_L0_0_L1_2_Wij_nx232), .CLK (CLK)) ;
    dff CACHE_L0_0_L1_2_Wij_reg_Dout_3 (.Q (CacheWindow_0__2__3), .QB (
        \$dummy [1345]), .D (CACHE_L0_0_L1_2_Wij_nx242), .CLK (CLK)) ;
    dff CACHE_L0_0_L1_2_Wij_reg_Dout_4 (.Q (CacheWindow_0__2__4), .QB (
        \$dummy [1346]), .D (CACHE_L0_0_L1_2_Wij_nx252), .CLK (CLK)) ;
    dff CACHE_L0_0_L1_2_Wij_reg_Dout_5 (.Q (CacheWindow_0__2__5), .QB (
        \$dummy [1347]), .D (CACHE_L0_0_L1_2_Wij_nx262), .CLK (CLK)) ;
    dff CACHE_L0_0_L1_2_Wij_reg_Dout_6 (.Q (CacheWindow_0__2__6), .QB (
        \$dummy [1348]), .D (CACHE_L0_0_L1_2_Wij_nx272), .CLK (CLK)) ;
    dff CACHE_L0_0_L1_2_Wij_reg_Dout_7 (.Q (CacheWindow_0__2__7), .QB (
        \$dummy [1349]), .D (CACHE_L0_0_L1_2_Wij_nx282), .CLK (CLK)) ;
    buf02 CACHE_L0_0_L1_2_Wij_ix330 (.Y (CACHE_L0_0_L1_2_Wij_nx331), .A (
          CACHE_EN_dup_1106)) ;
    buf02 CACHE_L0_0_L1_2_Wij_ix332 (.Y (CACHE_L0_0_L1_2_Wij_nx333), .A (
          CACHE_EN_dup_1106)) ;
    dff CACHE_L0_0_L1_3_Fij_reg_Dout_0 (.Q (CacheFilter_0__3__0), .QB (
        \$dummy [1350]), .D (CACHE_L0_0_L1_3_Fij_nx212), .CLK (CLK)) ;
    nor02_2x CACHE_L0_0_L1_3_Fij_ix297 (.Y (CACHE_L0_0_L1_3_Fij_nx296), .A0 (
             nx8369), .A1 (CACHE_L0_0_L1_3_Fij_nx331)) ;
    dff CACHE_L0_0_L1_3_Fij_reg_Dout_1 (.Q (CacheFilter_0__3__1), .QB (
        \$dummy [1351]), .D (CACHE_L0_0_L1_3_Fij_nx222), .CLK (CLK)) ;
    dff CACHE_L0_0_L1_3_Fij_reg_Dout_2 (.Q (CacheFilter_0__3__2), .QB (
        \$dummy [1352]), .D (CACHE_L0_0_L1_3_Fij_nx232), .CLK (CLK)) ;
    dff CACHE_L0_0_L1_3_Fij_reg_Dout_3 (.Q (CacheFilter_0__3__3), .QB (
        \$dummy [1353]), .D (CACHE_L0_0_L1_3_Fij_nx242), .CLK (CLK)) ;
    dff CACHE_L0_0_L1_3_Fij_reg_Dout_4 (.Q (CacheFilter_0__3__4), .QB (
        \$dummy [1354]), .D (CACHE_L0_0_L1_3_Fij_nx252), .CLK (CLK)) ;
    dff CACHE_L0_0_L1_3_Fij_reg_Dout_5 (.Q (CacheFilter_0__3__5), .QB (
        \$dummy [1355]), .D (CACHE_L0_0_L1_3_Fij_nx262), .CLK (CLK)) ;
    dff CACHE_L0_0_L1_3_Fij_reg_Dout_6 (.Q (CacheFilter_0__3__6), .QB (
        \$dummy [1356]), .D (CACHE_L0_0_L1_3_Fij_nx272), .CLK (CLK)) ;
    dff CACHE_L0_0_L1_3_Fij_reg_Dout_7 (.Q (CacheFilter_0__3__7), .QB (
        \$dummy [1357]), .D (CACHE_L0_0_L1_3_Fij_nx282), .CLK (CLK)) ;
    buf02 CACHE_L0_0_L1_3_Fij_ix330 (.Y (CACHE_L0_0_L1_3_Fij_nx331), .A (
          CACHE_EN_dup_1095)) ;
    buf02 CACHE_L0_0_L1_3_Fij_ix332 (.Y (CACHE_L0_0_L1_3_Fij_nx333), .A (
          CACHE_EN_dup_1095)) ;
    dff CACHE_L0_0_L1_3_Wij_reg_Dout_0 (.Q (CacheWindow_0__3__0), .QB (
        \$dummy [1358]), .D (CACHE_L0_0_L1_3_Wij_nx212), .CLK (CLK)) ;
    nor02_2x CACHE_L0_0_L1_3_Wij_ix297 (.Y (CACHE_L0_0_L1_3_Wij_nx296), .A0 (
             nx8369), .A1 (CACHE_L0_0_L1_3_Wij_nx331)) ;
    dff CACHE_L0_0_L1_3_Wij_reg_Dout_1 (.Q (CacheWindow_0__3__1), .QB (
        \$dummy [1359]), .D (CACHE_L0_0_L1_3_Wij_nx222), .CLK (CLK)) ;
    dff CACHE_L0_0_L1_3_Wij_reg_Dout_2 (.Q (CacheWindow_0__3__2), .QB (
        \$dummy [1360]), .D (CACHE_L0_0_L1_3_Wij_nx232), .CLK (CLK)) ;
    dff CACHE_L0_0_L1_3_Wij_reg_Dout_3 (.Q (CacheWindow_0__3__3), .QB (
        \$dummy [1361]), .D (CACHE_L0_0_L1_3_Wij_nx242), .CLK (CLK)) ;
    dff CACHE_L0_0_L1_3_Wij_reg_Dout_4 (.Q (CacheWindow_0__3__4), .QB (
        \$dummy [1362]), .D (CACHE_L0_0_L1_3_Wij_nx252), .CLK (CLK)) ;
    dff CACHE_L0_0_L1_3_Wij_reg_Dout_5 (.Q (CacheWindow_0__3__5), .QB (
        \$dummy [1363]), .D (CACHE_L0_0_L1_3_Wij_nx262), .CLK (CLK)) ;
    dff CACHE_L0_0_L1_3_Wij_reg_Dout_6 (.Q (CacheWindow_0__3__6), .QB (
        \$dummy [1364]), .D (CACHE_L0_0_L1_3_Wij_nx272), .CLK (CLK)) ;
    dff CACHE_L0_0_L1_3_Wij_reg_Dout_7 (.Q (CacheWindow_0__3__7), .QB (
        \$dummy [1365]), .D (CACHE_L0_0_L1_3_Wij_nx282), .CLK (CLK)) ;
    buf02 CACHE_L0_0_L1_3_Wij_ix330 (.Y (CACHE_L0_0_L1_3_Wij_nx331), .A (
          CACHE_EN_dup_1106)) ;
    buf02 CACHE_L0_0_L1_3_Wij_ix332 (.Y (CACHE_L0_0_L1_3_Wij_nx333), .A (
          CACHE_EN_dup_1106)) ;
    dff CACHE_L0_0_L1_4_Fij_reg_Dout_0 (.Q (CacheFilter_0__4__0), .QB (
        \$dummy [1366]), .D (CACHE_L0_0_L1_4_Fij_nx212), .CLK (CLK)) ;
    nor02_2x CACHE_L0_0_L1_4_Fij_ix297 (.Y (CACHE_L0_0_L1_4_Fij_nx296), .A0 (
             nx8373), .A1 (CACHE_L0_0_L1_4_Fij_nx331)) ;
    dff CACHE_L0_0_L1_4_Fij_reg_Dout_1 (.Q (CacheFilter_0__4__1), .QB (
        \$dummy [1367]), .D (CACHE_L0_0_L1_4_Fij_nx222), .CLK (CLK)) ;
    dff CACHE_L0_0_L1_4_Fij_reg_Dout_2 (.Q (CacheFilter_0__4__2), .QB (
        \$dummy [1368]), .D (CACHE_L0_0_L1_4_Fij_nx232), .CLK (CLK)) ;
    dff CACHE_L0_0_L1_4_Fij_reg_Dout_3 (.Q (CacheFilter_0__4__3), .QB (
        \$dummy [1369]), .D (CACHE_L0_0_L1_4_Fij_nx242), .CLK (CLK)) ;
    dff CACHE_L0_0_L1_4_Fij_reg_Dout_4 (.Q (CacheFilter_0__4__4), .QB (
        \$dummy [1370]), .D (CACHE_L0_0_L1_4_Fij_nx252), .CLK (CLK)) ;
    dff CACHE_L0_0_L1_4_Fij_reg_Dout_5 (.Q (CacheFilter_0__4__5), .QB (
        \$dummy [1371]), .D (CACHE_L0_0_L1_4_Fij_nx262), .CLK (CLK)) ;
    dff CACHE_L0_0_L1_4_Fij_reg_Dout_6 (.Q (CacheFilter_0__4__6), .QB (
        \$dummy [1372]), .D (CACHE_L0_0_L1_4_Fij_nx272), .CLK (CLK)) ;
    dff CACHE_L0_0_L1_4_Fij_reg_Dout_7 (.Q (CacheFilter_0__4__7), .QB (
        \$dummy [1373]), .D (CACHE_L0_0_L1_4_Fij_nx282), .CLK (CLK)) ;
    buf02 CACHE_L0_0_L1_4_Fij_ix330 (.Y (CACHE_L0_0_L1_4_Fij_nx331), .A (
          CACHE_EN_dup_1161)) ;
    buf02 CACHE_L0_0_L1_4_Fij_ix332 (.Y (CACHE_L0_0_L1_4_Fij_nx333), .A (
          CACHE_EN_dup_1161)) ;
    dff CACHE_L0_0_L1_4_Wij_reg_Dout_0 (.Q (CacheWindow_0__4__0), .QB (
        \$dummy [1374]), .D (CACHE_L0_0_L1_4_Wij_nx212), .CLK (CLK)) ;
    nor02_2x CACHE_L0_0_L1_4_Wij_ix297 (.Y (CACHE_L0_0_L1_4_Wij_nx296), .A0 (
             nx8373), .A1 (CACHE_L0_0_L1_4_Wij_nx331)) ;
    dff CACHE_L0_0_L1_4_Wij_reg_Dout_1 (.Q (CacheWindow_0__4__1), .QB (
        \$dummy [1375]), .D (CACHE_L0_0_L1_4_Wij_nx222), .CLK (CLK)) ;
    dff CACHE_L0_0_L1_4_Wij_reg_Dout_2 (.Q (CacheWindow_0__4__2), .QB (
        \$dummy [1376]), .D (CACHE_L0_0_L1_4_Wij_nx232), .CLK (CLK)) ;
    dff CACHE_L0_0_L1_4_Wij_reg_Dout_3 (.Q (CacheWindow_0__4__3), .QB (
        \$dummy [1377]), .D (CACHE_L0_0_L1_4_Wij_nx242), .CLK (CLK)) ;
    dff CACHE_L0_0_L1_4_Wij_reg_Dout_4 (.Q (CacheWindow_0__4__4), .QB (
        \$dummy [1378]), .D (CACHE_L0_0_L1_4_Wij_nx252), .CLK (CLK)) ;
    dff CACHE_L0_0_L1_4_Wij_reg_Dout_5 (.Q (CacheWindow_0__4__5), .QB (
        \$dummy [1379]), .D (CACHE_L0_0_L1_4_Wij_nx262), .CLK (CLK)) ;
    dff CACHE_L0_0_L1_4_Wij_reg_Dout_6 (.Q (CacheWindow_0__4__6), .QB (
        \$dummy [1380]), .D (CACHE_L0_0_L1_4_Wij_nx272), .CLK (CLK)) ;
    dff CACHE_L0_0_L1_4_Wij_reg_Dout_7 (.Q (CacheWindow_0__4__7), .QB (
        \$dummy [1381]), .D (CACHE_L0_0_L1_4_Wij_nx282), .CLK (CLK)) ;
    buf02 CACHE_L0_0_L1_4_Wij_ix330 (.Y (CACHE_L0_0_L1_4_Wij_nx331), .A (
          CACHE_EN_dup_1172)) ;
    buf02 CACHE_L0_0_L1_4_Wij_ix332 (.Y (CACHE_L0_0_L1_4_Wij_nx333), .A (
          CACHE_EN_dup_1172)) ;
    dff CACHE_L0_1_L1_0_Fij_reg_Dout_0 (.Q (CacheFilter_1__0__0), .QB (
        \$dummy [1382]), .D (CACHE_L0_1_L1_0_Fij_nx212), .CLK (CLK)) ;
    nor02_2x CACHE_L0_1_L1_0_Fij_ix297 (.Y (CACHE_L0_1_L1_0_Fij_nx296), .A0 (
             nx8377), .A1 (CACHE_L0_1_L1_0_Fij_nx331)) ;
    dff CACHE_L0_1_L1_0_Fij_reg_Dout_1 (.Q (CacheFilter_1__0__1), .QB (
        \$dummy [1383]), .D (CACHE_L0_1_L1_0_Fij_nx222), .CLK (CLK)) ;
    dff CACHE_L0_1_L1_0_Fij_reg_Dout_2 (.Q (CacheFilter_1__0__2), .QB (
        \$dummy [1384]), .D (CACHE_L0_1_L1_0_Fij_nx232), .CLK (CLK)) ;
    dff CACHE_L0_1_L1_0_Fij_reg_Dout_3 (.Q (CacheFilter_1__0__3), .QB (
        \$dummy [1385]), .D (CACHE_L0_1_L1_0_Fij_nx242), .CLK (CLK)) ;
    dff CACHE_L0_1_L1_0_Fij_reg_Dout_4 (.Q (CacheFilter_1__0__4), .QB (
        \$dummy [1386]), .D (CACHE_L0_1_L1_0_Fij_nx252), .CLK (CLK)) ;
    dff CACHE_L0_1_L1_0_Fij_reg_Dout_5 (.Q (CacheFilter_1__0__5), .QB (
        \$dummy [1387]), .D (CACHE_L0_1_L1_0_Fij_nx262), .CLK (CLK)) ;
    dff CACHE_L0_1_L1_0_Fij_reg_Dout_6 (.Q (CacheFilter_1__0__6), .QB (
        \$dummy [1388]), .D (CACHE_L0_1_L1_0_Fij_nx272), .CLK (CLK)) ;
    dff CACHE_L0_1_L1_0_Fij_reg_Dout_7 (.Q (CacheFilter_1__0__7), .QB (
        \$dummy [1389]), .D (CACHE_L0_1_L1_0_Fij_nx282), .CLK (CLK)) ;
    buf02 CACHE_L0_1_L1_0_Fij_ix330 (.Y (CACHE_L0_1_L1_0_Fij_nx331), .A (
          CACHE_EN_dup_1161)) ;
    buf02 CACHE_L0_1_L1_0_Fij_ix332 (.Y (CACHE_L0_1_L1_0_Fij_nx333), .A (
          CACHE_EN_dup_1161)) ;
    dff CACHE_L0_1_L1_0_Wij_reg_Dout_0 (.Q (CacheWindow_1__0__0), .QB (
        \$dummy [1390]), .D (CACHE_L0_1_L1_0_Wij_nx212), .CLK (CLK)) ;
    nor02_2x CACHE_L0_1_L1_0_Wij_ix297 (.Y (CACHE_L0_1_L1_0_Wij_nx296), .A0 (
             nx8377), .A1 (CACHE_L0_1_L1_0_Wij_nx331)) ;
    dff CACHE_L0_1_L1_0_Wij_reg_Dout_1 (.Q (CacheWindow_1__0__1), .QB (
        \$dummy [1391]), .D (CACHE_L0_1_L1_0_Wij_nx222), .CLK (CLK)) ;
    dff CACHE_L0_1_L1_0_Wij_reg_Dout_2 (.Q (CacheWindow_1__0__2), .QB (
        \$dummy [1392]), .D (CACHE_L0_1_L1_0_Wij_nx232), .CLK (CLK)) ;
    dff CACHE_L0_1_L1_0_Wij_reg_Dout_3 (.Q (CacheWindow_1__0__3), .QB (
        \$dummy [1393]), .D (CACHE_L0_1_L1_0_Wij_nx242), .CLK (CLK)) ;
    dff CACHE_L0_1_L1_0_Wij_reg_Dout_4 (.Q (CacheWindow_1__0__4), .QB (
        \$dummy [1394]), .D (CACHE_L0_1_L1_0_Wij_nx252), .CLK (CLK)) ;
    dff CACHE_L0_1_L1_0_Wij_reg_Dout_5 (.Q (CacheWindow_1__0__5), .QB (
        \$dummy [1395]), .D (CACHE_L0_1_L1_0_Wij_nx262), .CLK (CLK)) ;
    dff CACHE_L0_1_L1_0_Wij_reg_Dout_6 (.Q (CacheWindow_1__0__6), .QB (
        \$dummy [1396]), .D (CACHE_L0_1_L1_0_Wij_nx272), .CLK (CLK)) ;
    dff CACHE_L0_1_L1_0_Wij_reg_Dout_7 (.Q (CacheWindow_1__0__7), .QB (
        \$dummy [1397]), .D (CACHE_L0_1_L1_0_Wij_nx282), .CLK (CLK)) ;
    buf02 CACHE_L0_1_L1_0_Wij_ix330 (.Y (CACHE_L0_1_L1_0_Wij_nx331), .A (
          CACHE_EN_dup_1172)) ;
    buf02 CACHE_L0_1_L1_0_Wij_ix332 (.Y (CACHE_L0_1_L1_0_Wij_nx333), .A (
          CACHE_EN_dup_1172)) ;
    dff CACHE_L0_1_L1_1_Fij_reg_Dout_0 (.Q (CacheFilter_1__1__0), .QB (
        \$dummy [1398]), .D (CACHE_L0_1_L1_1_Fij_nx212), .CLK (CLK)) ;
    nor02_2x CACHE_L0_1_L1_1_Fij_ix297 (.Y (CACHE_L0_1_L1_1_Fij_nx296), .A0 (
             nx8381), .A1 (CACHE_L0_1_L1_1_Fij_nx331)) ;
    dff CACHE_L0_1_L1_1_Fij_reg_Dout_1 (.Q (CacheFilter_1__1__1), .QB (
        \$dummy [1399]), .D (CACHE_L0_1_L1_1_Fij_nx222), .CLK (CLK)) ;
    dff CACHE_L0_1_L1_1_Fij_reg_Dout_2 (.Q (CacheFilter_1__1__2), .QB (
        \$dummy [1400]), .D (CACHE_L0_1_L1_1_Fij_nx232), .CLK (CLK)) ;
    dff CACHE_L0_1_L1_1_Fij_reg_Dout_3 (.Q (CacheFilter_1__1__3), .QB (
        \$dummy [1401]), .D (CACHE_L0_1_L1_1_Fij_nx242), .CLK (CLK)) ;
    dff CACHE_L0_1_L1_1_Fij_reg_Dout_4 (.Q (CacheFilter_1__1__4), .QB (
        \$dummy [1402]), .D (CACHE_L0_1_L1_1_Fij_nx252), .CLK (CLK)) ;
    dff CACHE_L0_1_L1_1_Fij_reg_Dout_5 (.Q (CacheFilter_1__1__5), .QB (
        \$dummy [1403]), .D (CACHE_L0_1_L1_1_Fij_nx262), .CLK (CLK)) ;
    dff CACHE_L0_1_L1_1_Fij_reg_Dout_6 (.Q (CacheFilter_1__1__6), .QB (
        \$dummy [1404]), .D (CACHE_L0_1_L1_1_Fij_nx272), .CLK (CLK)) ;
    dff CACHE_L0_1_L1_1_Fij_reg_Dout_7 (.Q (CacheFilter_1__1__7), .QB (
        \$dummy [1405]), .D (CACHE_L0_1_L1_1_Fij_nx282), .CLK (CLK)) ;
    buf02 CACHE_L0_1_L1_1_Fij_ix330 (.Y (CACHE_L0_1_L1_1_Fij_nx331), .A (
          CACHE_EN_dup_1161)) ;
    buf02 CACHE_L0_1_L1_1_Fij_ix332 (.Y (CACHE_L0_1_L1_1_Fij_nx333), .A (
          CACHE_EN_dup_1161)) ;
    dff CACHE_L0_1_L1_1_Wij_reg_Dout_0 (.Q (CacheWindow_1__1__0), .QB (
        \$dummy [1406]), .D (CACHE_L0_1_L1_1_Wij_nx212), .CLK (CLK)) ;
    nor02_2x CACHE_L0_1_L1_1_Wij_ix297 (.Y (CACHE_L0_1_L1_1_Wij_nx296), .A0 (
             nx8381), .A1 (CACHE_L0_1_L1_1_Wij_nx331)) ;
    dff CACHE_L0_1_L1_1_Wij_reg_Dout_1 (.Q (CacheWindow_1__1__1), .QB (
        \$dummy [1407]), .D (CACHE_L0_1_L1_1_Wij_nx222), .CLK (CLK)) ;
    dff CACHE_L0_1_L1_1_Wij_reg_Dout_2 (.Q (CacheWindow_1__1__2), .QB (
        \$dummy [1408]), .D (CACHE_L0_1_L1_1_Wij_nx232), .CLK (CLK)) ;
    dff CACHE_L0_1_L1_1_Wij_reg_Dout_3 (.Q (CacheWindow_1__1__3), .QB (
        \$dummy [1409]), .D (CACHE_L0_1_L1_1_Wij_nx242), .CLK (CLK)) ;
    dff CACHE_L0_1_L1_1_Wij_reg_Dout_4 (.Q (CacheWindow_1__1__4), .QB (
        \$dummy [1410]), .D (CACHE_L0_1_L1_1_Wij_nx252), .CLK (CLK)) ;
    dff CACHE_L0_1_L1_1_Wij_reg_Dout_5 (.Q (CacheWindow_1__1__5), .QB (
        \$dummy [1411]), .D (CACHE_L0_1_L1_1_Wij_nx262), .CLK (CLK)) ;
    dff CACHE_L0_1_L1_1_Wij_reg_Dout_6 (.Q (CacheWindow_1__1__6), .QB (
        \$dummy [1412]), .D (CACHE_L0_1_L1_1_Wij_nx272), .CLK (CLK)) ;
    dff CACHE_L0_1_L1_1_Wij_reg_Dout_7 (.Q (CacheWindow_1__1__7), .QB (
        \$dummy [1413]), .D (CACHE_L0_1_L1_1_Wij_nx282), .CLK (CLK)) ;
    buf02 CACHE_L0_1_L1_1_Wij_ix330 (.Y (CACHE_L0_1_L1_1_Wij_nx331), .A (
          CACHE_EN_dup_1172)) ;
    buf02 CACHE_L0_1_L1_1_Wij_ix332 (.Y (CACHE_L0_1_L1_1_Wij_nx333), .A (
          CACHE_EN_dup_1172)) ;
    dff CACHE_L0_1_L1_2_Fij_reg_Dout_0 (.Q (CacheFilter_1__2__0), .QB (
        \$dummy [1414]), .D (CACHE_L0_1_L1_2_Fij_nx212), .CLK (CLK)) ;
    nor02_2x CACHE_L0_1_L1_2_Fij_ix297 (.Y (CACHE_L0_1_L1_2_Fij_nx296), .A0 (
             nx8385), .A1 (CACHE_L0_1_L1_2_Fij_nx331)) ;
    dff CACHE_L0_1_L1_2_Fij_reg_Dout_1 (.Q (CacheFilter_1__2__1), .QB (
        \$dummy [1415]), .D (CACHE_L0_1_L1_2_Fij_nx222), .CLK (CLK)) ;
    dff CACHE_L0_1_L1_2_Fij_reg_Dout_2 (.Q (CacheFilter_1__2__2), .QB (
        \$dummy [1416]), .D (CACHE_L0_1_L1_2_Fij_nx232), .CLK (CLK)) ;
    dff CACHE_L0_1_L1_2_Fij_reg_Dout_3 (.Q (CacheFilter_1__2__3), .QB (
        \$dummy [1417]), .D (CACHE_L0_1_L1_2_Fij_nx242), .CLK (CLK)) ;
    dff CACHE_L0_1_L1_2_Fij_reg_Dout_4 (.Q (CacheFilter_1__2__4), .QB (
        \$dummy [1418]), .D (CACHE_L0_1_L1_2_Fij_nx252), .CLK (CLK)) ;
    dff CACHE_L0_1_L1_2_Fij_reg_Dout_5 (.Q (CacheFilter_1__2__5), .QB (
        \$dummy [1419]), .D (CACHE_L0_1_L1_2_Fij_nx262), .CLK (CLK)) ;
    dff CACHE_L0_1_L1_2_Fij_reg_Dout_6 (.Q (CacheFilter_1__2__6), .QB (
        \$dummy [1420]), .D (CACHE_L0_1_L1_2_Fij_nx272), .CLK (CLK)) ;
    dff CACHE_L0_1_L1_2_Fij_reg_Dout_7 (.Q (CacheFilter_1__2__7), .QB (
        \$dummy [1421]), .D (CACHE_L0_1_L1_2_Fij_nx282), .CLK (CLK)) ;
    buf02 CACHE_L0_1_L1_2_Fij_ix330 (.Y (CACHE_L0_1_L1_2_Fij_nx331), .A (
          CACHE_EN_dup_1227)) ;
    buf02 CACHE_L0_1_L1_2_Fij_ix332 (.Y (CACHE_L0_1_L1_2_Fij_nx333), .A (
          CACHE_EN_dup_1227)) ;
    dff CACHE_L0_1_L1_2_Wij_reg_Dout_0 (.Q (CacheWindow_1__2__0), .QB (
        \$dummy [1422]), .D (CACHE_L0_1_L1_2_Wij_nx212), .CLK (CLK)) ;
    nor02_2x CACHE_L0_1_L1_2_Wij_ix297 (.Y (CACHE_L0_1_L1_2_Wij_nx296), .A0 (
             nx8385), .A1 (CACHE_L0_1_L1_2_Wij_nx331)) ;
    dff CACHE_L0_1_L1_2_Wij_reg_Dout_1 (.Q (CacheWindow_1__2__1), .QB (
        \$dummy [1423]), .D (CACHE_L0_1_L1_2_Wij_nx222), .CLK (CLK)) ;
    dff CACHE_L0_1_L1_2_Wij_reg_Dout_2 (.Q (CacheWindow_1__2__2), .QB (
        \$dummy [1424]), .D (CACHE_L0_1_L1_2_Wij_nx232), .CLK (CLK)) ;
    dff CACHE_L0_1_L1_2_Wij_reg_Dout_3 (.Q (CacheWindow_1__2__3), .QB (
        \$dummy [1425]), .D (CACHE_L0_1_L1_2_Wij_nx242), .CLK (CLK)) ;
    dff CACHE_L0_1_L1_2_Wij_reg_Dout_4 (.Q (CacheWindow_1__2__4), .QB (
        \$dummy [1426]), .D (CACHE_L0_1_L1_2_Wij_nx252), .CLK (CLK)) ;
    dff CACHE_L0_1_L1_2_Wij_reg_Dout_5 (.Q (CacheWindow_1__2__5), .QB (
        \$dummy [1427]), .D (CACHE_L0_1_L1_2_Wij_nx262), .CLK (CLK)) ;
    dff CACHE_L0_1_L1_2_Wij_reg_Dout_6 (.Q (CacheWindow_1__2__6), .QB (
        \$dummy [1428]), .D (CACHE_L0_1_L1_2_Wij_nx272), .CLK (CLK)) ;
    dff CACHE_L0_1_L1_2_Wij_reg_Dout_7 (.Q (CacheWindow_1__2__7), .QB (
        \$dummy [1429]), .D (CACHE_L0_1_L1_2_Wij_nx282), .CLK (CLK)) ;
    buf02 CACHE_L0_1_L1_2_Wij_ix330 (.Y (CACHE_L0_1_L1_2_Wij_nx331), .A (
          CACHE_EN_dup_1238)) ;
    buf02 CACHE_L0_1_L1_2_Wij_ix332 (.Y (CACHE_L0_1_L1_2_Wij_nx333), .A (
          CACHE_EN_dup_1238)) ;
    dff CACHE_L0_1_L1_3_Fij_reg_Dout_0 (.Q (CacheFilter_1__3__0), .QB (
        \$dummy [1430]), .D (CACHE_L0_1_L1_3_Fij_nx212), .CLK (CLK)) ;
    nor02_2x CACHE_L0_1_L1_3_Fij_ix297 (.Y (CACHE_L0_1_L1_3_Fij_nx296), .A0 (
             nx8389), .A1 (CACHE_L0_1_L1_3_Fij_nx331)) ;
    dff CACHE_L0_1_L1_3_Fij_reg_Dout_1 (.Q (CacheFilter_1__3__1), .QB (
        \$dummy [1431]), .D (CACHE_L0_1_L1_3_Fij_nx222), .CLK (CLK)) ;
    dff CACHE_L0_1_L1_3_Fij_reg_Dout_2 (.Q (CacheFilter_1__3__2), .QB (
        \$dummy [1432]), .D (CACHE_L0_1_L1_3_Fij_nx232), .CLK (CLK)) ;
    dff CACHE_L0_1_L1_3_Fij_reg_Dout_3 (.Q (CacheFilter_1__3__3), .QB (
        \$dummy [1433]), .D (CACHE_L0_1_L1_3_Fij_nx242), .CLK (CLK)) ;
    dff CACHE_L0_1_L1_3_Fij_reg_Dout_4 (.Q (CacheFilter_1__3__4), .QB (
        \$dummy [1434]), .D (CACHE_L0_1_L1_3_Fij_nx252), .CLK (CLK)) ;
    dff CACHE_L0_1_L1_3_Fij_reg_Dout_5 (.Q (CacheFilter_1__3__5), .QB (
        \$dummy [1435]), .D (CACHE_L0_1_L1_3_Fij_nx262), .CLK (CLK)) ;
    dff CACHE_L0_1_L1_3_Fij_reg_Dout_6 (.Q (CacheFilter_1__3__6), .QB (
        \$dummy [1436]), .D (CACHE_L0_1_L1_3_Fij_nx272), .CLK (CLK)) ;
    dff CACHE_L0_1_L1_3_Fij_reg_Dout_7 (.Q (CacheFilter_1__3__7), .QB (
        \$dummy [1437]), .D (CACHE_L0_1_L1_3_Fij_nx282), .CLK (CLK)) ;
    buf02 CACHE_L0_1_L1_3_Fij_ix330 (.Y (CACHE_L0_1_L1_3_Fij_nx331), .A (
          CACHE_EN_dup_1227)) ;
    buf02 CACHE_L0_1_L1_3_Fij_ix332 (.Y (CACHE_L0_1_L1_3_Fij_nx333), .A (
          CACHE_EN_dup_1227)) ;
    dff CACHE_L0_1_L1_3_Wij_reg_Dout_0 (.Q (CacheWindow_1__3__0), .QB (
        \$dummy [1438]), .D (CACHE_L0_1_L1_3_Wij_nx212), .CLK (CLK)) ;
    nor02_2x CACHE_L0_1_L1_3_Wij_ix297 (.Y (CACHE_L0_1_L1_3_Wij_nx296), .A0 (
             nx8389), .A1 (CACHE_L0_1_L1_3_Wij_nx331)) ;
    dff CACHE_L0_1_L1_3_Wij_reg_Dout_1 (.Q (CacheWindow_1__3__1), .QB (
        \$dummy [1439]), .D (CACHE_L0_1_L1_3_Wij_nx222), .CLK (CLK)) ;
    dff CACHE_L0_1_L1_3_Wij_reg_Dout_2 (.Q (CacheWindow_1__3__2), .QB (
        \$dummy [1440]), .D (CACHE_L0_1_L1_3_Wij_nx232), .CLK (CLK)) ;
    dff CACHE_L0_1_L1_3_Wij_reg_Dout_3 (.Q (CacheWindow_1__3__3), .QB (
        \$dummy [1441]), .D (CACHE_L0_1_L1_3_Wij_nx242), .CLK (CLK)) ;
    dff CACHE_L0_1_L1_3_Wij_reg_Dout_4 (.Q (CacheWindow_1__3__4), .QB (
        \$dummy [1442]), .D (CACHE_L0_1_L1_3_Wij_nx252), .CLK (CLK)) ;
    dff CACHE_L0_1_L1_3_Wij_reg_Dout_5 (.Q (CacheWindow_1__3__5), .QB (
        \$dummy [1443]), .D (CACHE_L0_1_L1_3_Wij_nx262), .CLK (CLK)) ;
    dff CACHE_L0_1_L1_3_Wij_reg_Dout_6 (.Q (CacheWindow_1__3__6), .QB (
        \$dummy [1444]), .D (CACHE_L0_1_L1_3_Wij_nx272), .CLK (CLK)) ;
    dff CACHE_L0_1_L1_3_Wij_reg_Dout_7 (.Q (CacheWindow_1__3__7), .QB (
        \$dummy [1445]), .D (CACHE_L0_1_L1_3_Wij_nx282), .CLK (CLK)) ;
    buf02 CACHE_L0_1_L1_3_Wij_ix330 (.Y (CACHE_L0_1_L1_3_Wij_nx331), .A (
          CACHE_EN_dup_1238)) ;
    buf02 CACHE_L0_1_L1_3_Wij_ix332 (.Y (CACHE_L0_1_L1_3_Wij_nx333), .A (
          CACHE_EN_dup_1238)) ;
    dff CACHE_L0_1_L1_4_Fij_reg_Dout_0 (.Q (CacheFilter_1__4__0), .QB (
        \$dummy [1446]), .D (CACHE_L0_1_L1_4_Fij_nx212), .CLK (CLK)) ;
    nor02_2x CACHE_L0_1_L1_4_Fij_ix297 (.Y (CACHE_L0_1_L1_4_Fij_nx296), .A0 (
             nx8393), .A1 (CACHE_L0_1_L1_4_Fij_nx331)) ;
    dff CACHE_L0_1_L1_4_Fij_reg_Dout_1 (.Q (CacheFilter_1__4__1), .QB (
        \$dummy [1447]), .D (CACHE_L0_1_L1_4_Fij_nx222), .CLK (CLK)) ;
    dff CACHE_L0_1_L1_4_Fij_reg_Dout_2 (.Q (CacheFilter_1__4__2), .QB (
        \$dummy [1448]), .D (CACHE_L0_1_L1_4_Fij_nx232), .CLK (CLK)) ;
    dff CACHE_L0_1_L1_4_Fij_reg_Dout_3 (.Q (CacheFilter_1__4__3), .QB (
        \$dummy [1449]), .D (CACHE_L0_1_L1_4_Fij_nx242), .CLK (CLK)) ;
    dff CACHE_L0_1_L1_4_Fij_reg_Dout_4 (.Q (CacheFilter_1__4__4), .QB (
        \$dummy [1450]), .D (CACHE_L0_1_L1_4_Fij_nx252), .CLK (CLK)) ;
    dff CACHE_L0_1_L1_4_Fij_reg_Dout_5 (.Q (CacheFilter_1__4__5), .QB (
        \$dummy [1451]), .D (CACHE_L0_1_L1_4_Fij_nx262), .CLK (CLK)) ;
    dff CACHE_L0_1_L1_4_Fij_reg_Dout_6 (.Q (CacheFilter_1__4__6), .QB (
        \$dummy [1452]), .D (CACHE_L0_1_L1_4_Fij_nx272), .CLK (CLK)) ;
    dff CACHE_L0_1_L1_4_Fij_reg_Dout_7 (.Q (CacheFilter_1__4__7), .QB (
        \$dummy [1453]), .D (CACHE_L0_1_L1_4_Fij_nx282), .CLK (CLK)) ;
    buf02 CACHE_L0_1_L1_4_Fij_ix330 (.Y (CACHE_L0_1_L1_4_Fij_nx331), .A (
          CACHE_EN_dup_1227)) ;
    buf02 CACHE_L0_1_L1_4_Fij_ix332 (.Y (CACHE_L0_1_L1_4_Fij_nx333), .A (
          CACHE_EN_dup_1227)) ;
    dff CACHE_L0_1_L1_4_Wij_reg_Dout_0 (.Q (CacheWindow_1__4__0), .QB (
        \$dummy [1454]), .D (CACHE_L0_1_L1_4_Wij_nx212), .CLK (CLK)) ;
    nor02_2x CACHE_L0_1_L1_4_Wij_ix297 (.Y (CACHE_L0_1_L1_4_Wij_nx296), .A0 (
             nx8393), .A1 (CACHE_L0_1_L1_4_Wij_nx331)) ;
    dff CACHE_L0_1_L1_4_Wij_reg_Dout_1 (.Q (CacheWindow_1__4__1), .QB (
        \$dummy [1455]), .D (CACHE_L0_1_L1_4_Wij_nx222), .CLK (CLK)) ;
    dff CACHE_L0_1_L1_4_Wij_reg_Dout_2 (.Q (CacheWindow_1__4__2), .QB (
        \$dummy [1456]), .D (CACHE_L0_1_L1_4_Wij_nx232), .CLK (CLK)) ;
    dff CACHE_L0_1_L1_4_Wij_reg_Dout_3 (.Q (CacheWindow_1__4__3), .QB (
        \$dummy [1457]), .D (CACHE_L0_1_L1_4_Wij_nx242), .CLK (CLK)) ;
    dff CACHE_L0_1_L1_4_Wij_reg_Dout_4 (.Q (CacheWindow_1__4__4), .QB (
        \$dummy [1458]), .D (CACHE_L0_1_L1_4_Wij_nx252), .CLK (CLK)) ;
    dff CACHE_L0_1_L1_4_Wij_reg_Dout_5 (.Q (CacheWindow_1__4__5), .QB (
        \$dummy [1459]), .D (CACHE_L0_1_L1_4_Wij_nx262), .CLK (CLK)) ;
    dff CACHE_L0_1_L1_4_Wij_reg_Dout_6 (.Q (CacheWindow_1__4__6), .QB (
        \$dummy [1460]), .D (CACHE_L0_1_L1_4_Wij_nx272), .CLK (CLK)) ;
    dff CACHE_L0_1_L1_4_Wij_reg_Dout_7 (.Q (CacheWindow_1__4__7), .QB (
        \$dummy [1461]), .D (CACHE_L0_1_L1_4_Wij_nx282), .CLK (CLK)) ;
    buf02 CACHE_L0_1_L1_4_Wij_ix330 (.Y (CACHE_L0_1_L1_4_Wij_nx331), .A (
          CACHE_EN_dup_1238)) ;
    buf02 CACHE_L0_1_L1_4_Wij_ix332 (.Y (CACHE_L0_1_L1_4_Wij_nx333), .A (
          CACHE_EN_dup_1238)) ;
    dff CACHE_L0_2_L1_0_Fij_reg_Dout_0 (.Q (CacheFilter_2__0__0), .QB (
        \$dummy [1462]), .D (CACHE_L0_2_L1_0_Fij_nx212), .CLK (CLK)) ;
    nor02_2x CACHE_L0_2_L1_0_Fij_ix297 (.Y (CACHE_L0_2_L1_0_Fij_nx296), .A0 (
             nx8397), .A1 (CACHE_L0_2_L1_0_Fij_nx331)) ;
    dff CACHE_L0_2_L1_0_Fij_reg_Dout_1 (.Q (CacheFilter_2__0__1), .QB (
        \$dummy [1463]), .D (CACHE_L0_2_L1_0_Fij_nx222), .CLK (CLK)) ;
    dff CACHE_L0_2_L1_0_Fij_reg_Dout_2 (.Q (CacheFilter_2__0__2), .QB (
        \$dummy [1464]), .D (CACHE_L0_2_L1_0_Fij_nx232), .CLK (CLK)) ;
    dff CACHE_L0_2_L1_0_Fij_reg_Dout_3 (.Q (CacheFilter_2__0__3), .QB (
        \$dummy [1465]), .D (CACHE_L0_2_L1_0_Fij_nx242), .CLK (CLK)) ;
    dff CACHE_L0_2_L1_0_Fij_reg_Dout_4 (.Q (CacheFilter_2__0__4), .QB (
        \$dummy [1466]), .D (CACHE_L0_2_L1_0_Fij_nx252), .CLK (CLK)) ;
    dff CACHE_L0_2_L1_0_Fij_reg_Dout_5 (.Q (CacheFilter_2__0__5), .QB (
        \$dummy [1467]), .D (CACHE_L0_2_L1_0_Fij_nx262), .CLK (CLK)) ;
    dff CACHE_L0_2_L1_0_Fij_reg_Dout_6 (.Q (CacheFilter_2__0__6), .QB (
        \$dummy [1468]), .D (CACHE_L0_2_L1_0_Fij_nx272), .CLK (CLK)) ;
    dff CACHE_L0_2_L1_0_Fij_reg_Dout_7 (.Q (CacheFilter_2__0__7), .QB (
        \$dummy [1469]), .D (CACHE_L0_2_L1_0_Fij_nx282), .CLK (CLK)) ;
    buf02 CACHE_L0_2_L1_0_Fij_ix330 (.Y (CACHE_L0_2_L1_0_Fij_nx331), .A (
          CACHE_EN_dup_1293)) ;
    buf02 CACHE_L0_2_L1_0_Fij_ix332 (.Y (CACHE_L0_2_L1_0_Fij_nx333), .A (
          CACHE_EN_dup_1293)) ;
    dff CACHE_L0_2_L1_0_Wij_reg_Dout_0 (.Q (CacheWindow_2__0__0), .QB (
        \$dummy [1470]), .D (CACHE_L0_2_L1_0_Wij_nx212), .CLK (CLK)) ;
    nor02_2x CACHE_L0_2_L1_0_Wij_ix297 (.Y (CACHE_L0_2_L1_0_Wij_nx296), .A0 (
             nx8397), .A1 (CACHE_L0_2_L1_0_Wij_nx331)) ;
    dff CACHE_L0_2_L1_0_Wij_reg_Dout_1 (.Q (CacheWindow_2__0__1), .QB (
        \$dummy [1471]), .D (CACHE_L0_2_L1_0_Wij_nx222), .CLK (CLK)) ;
    dff CACHE_L0_2_L1_0_Wij_reg_Dout_2 (.Q (CacheWindow_2__0__2), .QB (
        \$dummy [1472]), .D (CACHE_L0_2_L1_0_Wij_nx232), .CLK (CLK)) ;
    dff CACHE_L0_2_L1_0_Wij_reg_Dout_3 (.Q (CacheWindow_2__0__3), .QB (
        \$dummy [1473]), .D (CACHE_L0_2_L1_0_Wij_nx242), .CLK (CLK)) ;
    dff CACHE_L0_2_L1_0_Wij_reg_Dout_4 (.Q (CacheWindow_2__0__4), .QB (
        \$dummy [1474]), .D (CACHE_L0_2_L1_0_Wij_nx252), .CLK (CLK)) ;
    dff CACHE_L0_2_L1_0_Wij_reg_Dout_5 (.Q (CacheWindow_2__0__5), .QB (
        \$dummy [1475]), .D (CACHE_L0_2_L1_0_Wij_nx262), .CLK (CLK)) ;
    dff CACHE_L0_2_L1_0_Wij_reg_Dout_6 (.Q (CacheWindow_2__0__6), .QB (
        \$dummy [1476]), .D (CACHE_L0_2_L1_0_Wij_nx272), .CLK (CLK)) ;
    dff CACHE_L0_2_L1_0_Wij_reg_Dout_7 (.Q (CacheWindow_2__0__7), .QB (
        \$dummy [1477]), .D (CACHE_L0_2_L1_0_Wij_nx282), .CLK (CLK)) ;
    buf02 CACHE_L0_2_L1_0_Wij_ix330 (.Y (CACHE_L0_2_L1_0_Wij_nx331), .A (
          CACHE_EN_dup_1304)) ;
    buf02 CACHE_L0_2_L1_0_Wij_ix332 (.Y (CACHE_L0_2_L1_0_Wij_nx333), .A (
          CACHE_EN_dup_1304)) ;
    dff CACHE_L0_2_L1_1_Fij_reg_Dout_0 (.Q (CacheFilter_2__1__0), .QB (
        \$dummy [1478]), .D (CACHE_L0_2_L1_1_Fij_nx212), .CLK (CLK)) ;
    nor02_2x CACHE_L0_2_L1_1_Fij_ix297 (.Y (CACHE_L0_2_L1_1_Fij_nx296), .A0 (
             nx8401), .A1 (CACHE_L0_2_L1_1_Fij_nx331)) ;
    dff CACHE_L0_2_L1_1_Fij_reg_Dout_1 (.Q (CacheFilter_2__1__1), .QB (
        \$dummy [1479]), .D (CACHE_L0_2_L1_1_Fij_nx222), .CLK (CLK)) ;
    dff CACHE_L0_2_L1_1_Fij_reg_Dout_2 (.Q (CacheFilter_2__1__2), .QB (
        \$dummy [1480]), .D (CACHE_L0_2_L1_1_Fij_nx232), .CLK (CLK)) ;
    dff CACHE_L0_2_L1_1_Fij_reg_Dout_3 (.Q (CacheFilter_2__1__3), .QB (
        \$dummy [1481]), .D (CACHE_L0_2_L1_1_Fij_nx242), .CLK (CLK)) ;
    dff CACHE_L0_2_L1_1_Fij_reg_Dout_4 (.Q (CacheFilter_2__1__4), .QB (
        \$dummy [1482]), .D (CACHE_L0_2_L1_1_Fij_nx252), .CLK (CLK)) ;
    dff CACHE_L0_2_L1_1_Fij_reg_Dout_5 (.Q (CacheFilter_2__1__5), .QB (
        \$dummy [1483]), .D (CACHE_L0_2_L1_1_Fij_nx262), .CLK (CLK)) ;
    dff CACHE_L0_2_L1_1_Fij_reg_Dout_6 (.Q (CacheFilter_2__1__6), .QB (
        \$dummy [1484]), .D (CACHE_L0_2_L1_1_Fij_nx272), .CLK (CLK)) ;
    dff CACHE_L0_2_L1_1_Fij_reg_Dout_7 (.Q (CacheFilter_2__1__7), .QB (
        \$dummy [1485]), .D (CACHE_L0_2_L1_1_Fij_nx282), .CLK (CLK)) ;
    buf02 CACHE_L0_2_L1_1_Fij_ix330 (.Y (CACHE_L0_2_L1_1_Fij_nx331), .A (
          CACHE_EN_dup_1293)) ;
    buf02 CACHE_L0_2_L1_1_Fij_ix332 (.Y (CACHE_L0_2_L1_1_Fij_nx333), .A (
          CACHE_EN_dup_1293)) ;
    dff CACHE_L0_2_L1_1_Wij_reg_Dout_0 (.Q (CacheWindow_2__1__0), .QB (
        \$dummy [1486]), .D (CACHE_L0_2_L1_1_Wij_nx212), .CLK (CLK)) ;
    nor02_2x CACHE_L0_2_L1_1_Wij_ix297 (.Y (CACHE_L0_2_L1_1_Wij_nx296), .A0 (
             nx8401), .A1 (CACHE_L0_2_L1_1_Wij_nx331)) ;
    dff CACHE_L0_2_L1_1_Wij_reg_Dout_1 (.Q (CacheWindow_2__1__1), .QB (
        \$dummy [1487]), .D (CACHE_L0_2_L1_1_Wij_nx222), .CLK (CLK)) ;
    dff CACHE_L0_2_L1_1_Wij_reg_Dout_2 (.Q (CacheWindow_2__1__2), .QB (
        \$dummy [1488]), .D (CACHE_L0_2_L1_1_Wij_nx232), .CLK (CLK)) ;
    dff CACHE_L0_2_L1_1_Wij_reg_Dout_3 (.Q (CacheWindow_2__1__3), .QB (
        \$dummy [1489]), .D (CACHE_L0_2_L1_1_Wij_nx242), .CLK (CLK)) ;
    dff CACHE_L0_2_L1_1_Wij_reg_Dout_4 (.Q (CacheWindow_2__1__4), .QB (
        \$dummy [1490]), .D (CACHE_L0_2_L1_1_Wij_nx252), .CLK (CLK)) ;
    dff CACHE_L0_2_L1_1_Wij_reg_Dout_5 (.Q (CacheWindow_2__1__5), .QB (
        \$dummy [1491]), .D (CACHE_L0_2_L1_1_Wij_nx262), .CLK (CLK)) ;
    dff CACHE_L0_2_L1_1_Wij_reg_Dout_6 (.Q (CacheWindow_2__1__6), .QB (
        \$dummy [1492]), .D (CACHE_L0_2_L1_1_Wij_nx272), .CLK (CLK)) ;
    dff CACHE_L0_2_L1_1_Wij_reg_Dout_7 (.Q (CacheWindow_2__1__7), .QB (
        \$dummy [1493]), .D (CACHE_L0_2_L1_1_Wij_nx282), .CLK (CLK)) ;
    buf02 CACHE_L0_2_L1_1_Wij_ix330 (.Y (CACHE_L0_2_L1_1_Wij_nx331), .A (
          CACHE_EN_dup_1304)) ;
    buf02 CACHE_L0_2_L1_1_Wij_ix332 (.Y (CACHE_L0_2_L1_1_Wij_nx333), .A (
          CACHE_EN_dup_1304)) ;
    dff CACHE_L0_2_L1_2_Fij_reg_Dout_0 (.Q (CacheFilter_2__2__0), .QB (
        \$dummy [1494]), .D (CACHE_L0_2_L1_2_Fij_nx212), .CLK (CLK)) ;
    nor02_2x CACHE_L0_2_L1_2_Fij_ix297 (.Y (CACHE_L0_2_L1_2_Fij_nx296), .A0 (
             nx8405), .A1 (CACHE_L0_2_L1_2_Fij_nx331)) ;
    dff CACHE_L0_2_L1_2_Fij_reg_Dout_1 (.Q (CacheFilter_2__2__1), .QB (
        \$dummy [1495]), .D (CACHE_L0_2_L1_2_Fij_nx222), .CLK (CLK)) ;
    dff CACHE_L0_2_L1_2_Fij_reg_Dout_2 (.Q (CacheFilter_2__2__2), .QB (
        \$dummy [1496]), .D (CACHE_L0_2_L1_2_Fij_nx232), .CLK (CLK)) ;
    dff CACHE_L0_2_L1_2_Fij_reg_Dout_3 (.Q (CacheFilter_2__2__3), .QB (
        \$dummy [1497]), .D (CACHE_L0_2_L1_2_Fij_nx242), .CLK (CLK)) ;
    dff CACHE_L0_2_L1_2_Fij_reg_Dout_4 (.Q (CacheFilter_2__2__4), .QB (
        \$dummy [1498]), .D (CACHE_L0_2_L1_2_Fij_nx252), .CLK (CLK)) ;
    dff CACHE_L0_2_L1_2_Fij_reg_Dout_5 (.Q (CacheFilter_2__2__5), .QB (
        \$dummy [1499]), .D (CACHE_L0_2_L1_2_Fij_nx262), .CLK (CLK)) ;
    dff CACHE_L0_2_L1_2_Fij_reg_Dout_6 (.Q (CacheFilter_2__2__6), .QB (
        \$dummy [1500]), .D (CACHE_L0_2_L1_2_Fij_nx272), .CLK (CLK)) ;
    dff CACHE_L0_2_L1_2_Fij_reg_Dout_7 (.Q (CacheFilter_2__2__7), .QB (
        \$dummy [1501]), .D (CACHE_L0_2_L1_2_Fij_nx282), .CLK (CLK)) ;
    buf02 CACHE_L0_2_L1_2_Fij_ix330 (.Y (CACHE_L0_2_L1_2_Fij_nx331), .A (
          CACHE_EN_dup_1293)) ;
    buf02 CACHE_L0_2_L1_2_Fij_ix332 (.Y (CACHE_L0_2_L1_2_Fij_nx333), .A (
          CACHE_EN_dup_1293)) ;
    dff CACHE_L0_2_L1_2_Wij_reg_Dout_0 (.Q (CacheWindow_2__2__0), .QB (
        \$dummy [1502]), .D (CACHE_L0_2_L1_2_Wij_nx212), .CLK (CLK)) ;
    nor02_2x CACHE_L0_2_L1_2_Wij_ix297 (.Y (CACHE_L0_2_L1_2_Wij_nx296), .A0 (
             nx8405), .A1 (CACHE_L0_2_L1_2_Wij_nx331)) ;
    dff CACHE_L0_2_L1_2_Wij_reg_Dout_1 (.Q (CacheWindow_2__2__1), .QB (
        \$dummy [1503]), .D (CACHE_L0_2_L1_2_Wij_nx222), .CLK (CLK)) ;
    dff CACHE_L0_2_L1_2_Wij_reg_Dout_2 (.Q (CacheWindow_2__2__2), .QB (
        \$dummy [1504]), .D (CACHE_L0_2_L1_2_Wij_nx232), .CLK (CLK)) ;
    dff CACHE_L0_2_L1_2_Wij_reg_Dout_3 (.Q (CacheWindow_2__2__3), .QB (
        \$dummy [1505]), .D (CACHE_L0_2_L1_2_Wij_nx242), .CLK (CLK)) ;
    dff CACHE_L0_2_L1_2_Wij_reg_Dout_4 (.Q (CacheWindow_2__2__4), .QB (
        \$dummy [1506]), .D (CACHE_L0_2_L1_2_Wij_nx252), .CLK (CLK)) ;
    dff CACHE_L0_2_L1_2_Wij_reg_Dout_5 (.Q (CacheWindow_2__2__5), .QB (
        \$dummy [1507]), .D (CACHE_L0_2_L1_2_Wij_nx262), .CLK (CLK)) ;
    dff CACHE_L0_2_L1_2_Wij_reg_Dout_6 (.Q (CacheWindow_2__2__6), .QB (
        \$dummy [1508]), .D (CACHE_L0_2_L1_2_Wij_nx272), .CLK (CLK)) ;
    dff CACHE_L0_2_L1_2_Wij_reg_Dout_7 (.Q (CacheWindow_2__2__7), .QB (
        \$dummy [1509]), .D (CACHE_L0_2_L1_2_Wij_nx282), .CLK (CLK)) ;
    buf02 CACHE_L0_2_L1_2_Wij_ix330 (.Y (CACHE_L0_2_L1_2_Wij_nx331), .A (
          CACHE_EN_dup_1304)) ;
    buf02 CACHE_L0_2_L1_2_Wij_ix332 (.Y (CACHE_L0_2_L1_2_Wij_nx333), .A (
          CACHE_EN_dup_1304)) ;
    dff CACHE_L0_2_L1_3_Fij_reg_Dout_0 (.Q (CacheFilter_2__3__0), .QB (
        \$dummy [1510]), .D (CACHE_L0_2_L1_3_Fij_nx212), .CLK (CLK)) ;
    nor02_2x CACHE_L0_2_L1_3_Fij_ix297 (.Y (CACHE_L0_2_L1_3_Fij_nx296), .A0 (
             nx8409), .A1 (CACHE_L0_2_L1_3_Fij_nx331)) ;
    dff CACHE_L0_2_L1_3_Fij_reg_Dout_1 (.Q (CacheFilter_2__3__1), .QB (
        \$dummy [1511]), .D (CACHE_L0_2_L1_3_Fij_nx222), .CLK (CLK)) ;
    dff CACHE_L0_2_L1_3_Fij_reg_Dout_2 (.Q (CacheFilter_2__3__2), .QB (
        \$dummy [1512]), .D (CACHE_L0_2_L1_3_Fij_nx232), .CLK (CLK)) ;
    dff CACHE_L0_2_L1_3_Fij_reg_Dout_3 (.Q (CacheFilter_2__3__3), .QB (
        \$dummy [1513]), .D (CACHE_L0_2_L1_3_Fij_nx242), .CLK (CLK)) ;
    dff CACHE_L0_2_L1_3_Fij_reg_Dout_4 (.Q (CacheFilter_2__3__4), .QB (
        \$dummy [1514]), .D (CACHE_L0_2_L1_3_Fij_nx252), .CLK (CLK)) ;
    dff CACHE_L0_2_L1_3_Fij_reg_Dout_5 (.Q (CacheFilter_2__3__5), .QB (
        \$dummy [1515]), .D (CACHE_L0_2_L1_3_Fij_nx262), .CLK (CLK)) ;
    dff CACHE_L0_2_L1_3_Fij_reg_Dout_6 (.Q (CacheFilter_2__3__6), .QB (
        \$dummy [1516]), .D (CACHE_L0_2_L1_3_Fij_nx272), .CLK (CLK)) ;
    dff CACHE_L0_2_L1_3_Fij_reg_Dout_7 (.Q (CacheFilter_2__3__7), .QB (
        \$dummy [1517]), .D (CACHE_L0_2_L1_3_Fij_nx282), .CLK (CLK)) ;
    buf02 CACHE_L0_2_L1_3_Fij_ix330 (.Y (CACHE_L0_2_L1_3_Fij_nx331), .A (
          CACHE_EN_dup_1359)) ;
    buf02 CACHE_L0_2_L1_3_Fij_ix332 (.Y (CACHE_L0_2_L1_3_Fij_nx333), .A (
          CACHE_EN_dup_1359)) ;
    dff CACHE_L0_2_L1_3_Wij_reg_Dout_0 (.Q (CacheWindow_2__3__0), .QB (
        \$dummy [1518]), .D (CACHE_L0_2_L1_3_Wij_nx212), .CLK (CLK)) ;
    nor02_2x CACHE_L0_2_L1_3_Wij_ix297 (.Y (CACHE_L0_2_L1_3_Wij_nx296), .A0 (
             nx8409), .A1 (CACHE_L0_2_L1_3_Wij_nx331)) ;
    dff CACHE_L0_2_L1_3_Wij_reg_Dout_1 (.Q (CacheWindow_2__3__1), .QB (
        \$dummy [1519]), .D (CACHE_L0_2_L1_3_Wij_nx222), .CLK (CLK)) ;
    dff CACHE_L0_2_L1_3_Wij_reg_Dout_2 (.Q (CacheWindow_2__3__2), .QB (
        \$dummy [1520]), .D (CACHE_L0_2_L1_3_Wij_nx232), .CLK (CLK)) ;
    dff CACHE_L0_2_L1_3_Wij_reg_Dout_3 (.Q (CacheWindow_2__3__3), .QB (
        \$dummy [1521]), .D (CACHE_L0_2_L1_3_Wij_nx242), .CLK (CLK)) ;
    dff CACHE_L0_2_L1_3_Wij_reg_Dout_4 (.Q (CacheWindow_2__3__4), .QB (
        \$dummy [1522]), .D (CACHE_L0_2_L1_3_Wij_nx252), .CLK (CLK)) ;
    dff CACHE_L0_2_L1_3_Wij_reg_Dout_5 (.Q (CacheWindow_2__3__5), .QB (
        \$dummy [1523]), .D (CACHE_L0_2_L1_3_Wij_nx262), .CLK (CLK)) ;
    dff CACHE_L0_2_L1_3_Wij_reg_Dout_6 (.Q (CacheWindow_2__3__6), .QB (
        \$dummy [1524]), .D (CACHE_L0_2_L1_3_Wij_nx272), .CLK (CLK)) ;
    dff CACHE_L0_2_L1_3_Wij_reg_Dout_7 (.Q (CacheWindow_2__3__7), .QB (
        \$dummy [1525]), .D (CACHE_L0_2_L1_3_Wij_nx282), .CLK (CLK)) ;
    buf02 CACHE_L0_2_L1_3_Wij_ix330 (.Y (CACHE_L0_2_L1_3_Wij_nx331), .A (
          CACHE_EN_dup_1370)) ;
    buf02 CACHE_L0_2_L1_3_Wij_ix332 (.Y (CACHE_L0_2_L1_3_Wij_nx333), .A (
          CACHE_EN_dup_1370)) ;
    dff CACHE_L0_2_L1_4_Fij_reg_Dout_0 (.Q (CacheFilter_2__4__0), .QB (
        \$dummy [1526]), .D (CACHE_L0_2_L1_4_Fij_nx212), .CLK (CLK)) ;
    nor02_2x CACHE_L0_2_L1_4_Fij_ix297 (.Y (CACHE_L0_2_L1_4_Fij_nx296), .A0 (
             nx8413), .A1 (CACHE_L0_2_L1_4_Fij_nx331)) ;
    dff CACHE_L0_2_L1_4_Fij_reg_Dout_1 (.Q (CacheFilter_2__4__1), .QB (
        \$dummy [1527]), .D (CACHE_L0_2_L1_4_Fij_nx222), .CLK (CLK)) ;
    dff CACHE_L0_2_L1_4_Fij_reg_Dout_2 (.Q (CacheFilter_2__4__2), .QB (
        \$dummy [1528]), .D (CACHE_L0_2_L1_4_Fij_nx232), .CLK (CLK)) ;
    dff CACHE_L0_2_L1_4_Fij_reg_Dout_3 (.Q (CacheFilter_2__4__3), .QB (
        \$dummy [1529]), .D (CACHE_L0_2_L1_4_Fij_nx242), .CLK (CLK)) ;
    dff CACHE_L0_2_L1_4_Fij_reg_Dout_4 (.Q (CacheFilter_2__4__4), .QB (
        \$dummy [1530]), .D (CACHE_L0_2_L1_4_Fij_nx252), .CLK (CLK)) ;
    dff CACHE_L0_2_L1_4_Fij_reg_Dout_5 (.Q (CacheFilter_2__4__5), .QB (
        \$dummy [1531]), .D (CACHE_L0_2_L1_4_Fij_nx262), .CLK (CLK)) ;
    dff CACHE_L0_2_L1_4_Fij_reg_Dout_6 (.Q (CacheFilter_2__4__6), .QB (
        \$dummy [1532]), .D (CACHE_L0_2_L1_4_Fij_nx272), .CLK (CLK)) ;
    dff CACHE_L0_2_L1_4_Fij_reg_Dout_7 (.Q (CacheFilter_2__4__7), .QB (
        \$dummy [1533]), .D (CACHE_L0_2_L1_4_Fij_nx282), .CLK (CLK)) ;
    buf02 CACHE_L0_2_L1_4_Fij_ix330 (.Y (CACHE_L0_2_L1_4_Fij_nx331), .A (
          CACHE_EN_dup_1359)) ;
    buf02 CACHE_L0_2_L1_4_Fij_ix332 (.Y (CACHE_L0_2_L1_4_Fij_nx333), .A (
          CACHE_EN_dup_1359)) ;
    dff CACHE_L0_2_L1_4_Wij_reg_Dout_0 (.Q (CacheWindow_2__4__0), .QB (
        \$dummy [1534]), .D (CACHE_L0_2_L1_4_Wij_nx212), .CLK (CLK)) ;
    nor02_2x CACHE_L0_2_L1_4_Wij_ix297 (.Y (CACHE_L0_2_L1_4_Wij_nx296), .A0 (
             nx8413), .A1 (CACHE_L0_2_L1_4_Wij_nx331)) ;
    dff CACHE_L0_2_L1_4_Wij_reg_Dout_1 (.Q (CacheWindow_2__4__1), .QB (
        \$dummy [1535]), .D (CACHE_L0_2_L1_4_Wij_nx222), .CLK (CLK)) ;
    dff CACHE_L0_2_L1_4_Wij_reg_Dout_2 (.Q (CacheWindow_2__4__2), .QB (
        \$dummy [1536]), .D (CACHE_L0_2_L1_4_Wij_nx232), .CLK (CLK)) ;
    dff CACHE_L0_2_L1_4_Wij_reg_Dout_3 (.Q (CacheWindow_2__4__3), .QB (
        \$dummy [1537]), .D (CACHE_L0_2_L1_4_Wij_nx242), .CLK (CLK)) ;
    dff CACHE_L0_2_L1_4_Wij_reg_Dout_4 (.Q (CacheWindow_2__4__4), .QB (
        \$dummy [1538]), .D (CACHE_L0_2_L1_4_Wij_nx252), .CLK (CLK)) ;
    dff CACHE_L0_2_L1_4_Wij_reg_Dout_5 (.Q (CacheWindow_2__4__5), .QB (
        \$dummy [1539]), .D (CACHE_L0_2_L1_4_Wij_nx262), .CLK (CLK)) ;
    dff CACHE_L0_2_L1_4_Wij_reg_Dout_6 (.Q (CacheWindow_2__4__6), .QB (
        \$dummy [1540]), .D (CACHE_L0_2_L1_4_Wij_nx272), .CLK (CLK)) ;
    dff CACHE_L0_2_L1_4_Wij_reg_Dout_7 (.Q (CacheWindow_2__4__7), .QB (
        \$dummy [1541]), .D (CACHE_L0_2_L1_4_Wij_nx282), .CLK (CLK)) ;
    buf02 CACHE_L0_2_L1_4_Wij_ix330 (.Y (CACHE_L0_2_L1_4_Wij_nx331), .A (
          CACHE_EN_dup_1370)) ;
    buf02 CACHE_L0_2_L1_4_Wij_ix332 (.Y (CACHE_L0_2_L1_4_Wij_nx333), .A (
          CACHE_EN_dup_1370)) ;
    dff CACHE_L0_3_L1_0_Fij_reg_Dout_0 (.Q (CacheFilter_3__0__0), .QB (
        \$dummy [1542]), .D (CACHE_L0_3_L1_0_Fij_nx212), .CLK (CLK)) ;
    nor02_2x CACHE_L0_3_L1_0_Fij_ix297 (.Y (CACHE_L0_3_L1_0_Fij_nx296), .A0 (
             nx8417), .A1 (CACHE_L0_3_L1_0_Fij_nx331)) ;
    dff CACHE_L0_3_L1_0_Fij_reg_Dout_1 (.Q (CacheFilter_3__0__1), .QB (
        \$dummy [1543]), .D (CACHE_L0_3_L1_0_Fij_nx222), .CLK (CLK)) ;
    dff CACHE_L0_3_L1_0_Fij_reg_Dout_2 (.Q (CacheFilter_3__0__2), .QB (
        \$dummy [1544]), .D (CACHE_L0_3_L1_0_Fij_nx232), .CLK (CLK)) ;
    dff CACHE_L0_3_L1_0_Fij_reg_Dout_3 (.Q (CacheFilter_3__0__3), .QB (
        \$dummy [1545]), .D (CACHE_L0_3_L1_0_Fij_nx242), .CLK (CLK)) ;
    dff CACHE_L0_3_L1_0_Fij_reg_Dout_4 (.Q (CacheFilter_3__0__4), .QB (
        \$dummy [1546]), .D (CACHE_L0_3_L1_0_Fij_nx252), .CLK (CLK)) ;
    dff CACHE_L0_3_L1_0_Fij_reg_Dout_5 (.Q (CacheFilter_3__0__5), .QB (
        \$dummy [1547]), .D (CACHE_L0_3_L1_0_Fij_nx262), .CLK (CLK)) ;
    dff CACHE_L0_3_L1_0_Fij_reg_Dout_6 (.Q (CacheFilter_3__0__6), .QB (
        \$dummy [1548]), .D (CACHE_L0_3_L1_0_Fij_nx272), .CLK (CLK)) ;
    dff CACHE_L0_3_L1_0_Fij_reg_Dout_7 (.Q (CacheFilter_3__0__7), .QB (
        \$dummy [1549]), .D (CACHE_L0_3_L1_0_Fij_nx282), .CLK (CLK)) ;
    buf02 CACHE_L0_3_L1_0_Fij_ix330 (.Y (CACHE_L0_3_L1_0_Fij_nx331), .A (
          CACHE_EN_dup_1403)) ;
    buf02 CACHE_L0_3_L1_0_Fij_ix332 (.Y (CACHE_L0_3_L1_0_Fij_nx333), .A (
          CACHE_EN_dup_1403)) ;
    dff CACHE_L0_3_L1_0_Wij_reg_Dout_0 (.Q (CacheWindow_3__0__0), .QB (
        \$dummy [1550]), .D (CACHE_L0_3_L1_0_Wij_nx212), .CLK (CLK)) ;
    nor02_2x CACHE_L0_3_L1_0_Wij_ix297 (.Y (CACHE_L0_3_L1_0_Wij_nx296), .A0 (
             nx8417), .A1 (CACHE_L0_3_L1_0_Wij_nx331)) ;
    dff CACHE_L0_3_L1_0_Wij_reg_Dout_1 (.Q (CacheWindow_3__0__1), .QB (
        \$dummy [1551]), .D (CACHE_L0_3_L1_0_Wij_nx222), .CLK (CLK)) ;
    dff CACHE_L0_3_L1_0_Wij_reg_Dout_2 (.Q (CacheWindow_3__0__2), .QB (
        \$dummy [1552]), .D (CACHE_L0_3_L1_0_Wij_nx232), .CLK (CLK)) ;
    dff CACHE_L0_3_L1_0_Wij_reg_Dout_3 (.Q (CacheWindow_3__0__3), .QB (
        \$dummy [1553]), .D (CACHE_L0_3_L1_0_Wij_nx242), .CLK (CLK)) ;
    dff CACHE_L0_3_L1_0_Wij_reg_Dout_4 (.Q (CacheWindow_3__0__4), .QB (
        \$dummy [1554]), .D (CACHE_L0_3_L1_0_Wij_nx252), .CLK (CLK)) ;
    dff CACHE_L0_3_L1_0_Wij_reg_Dout_5 (.Q (CacheWindow_3__0__5), .QB (
        \$dummy [1555]), .D (CACHE_L0_3_L1_0_Wij_nx262), .CLK (CLK)) ;
    dff CACHE_L0_3_L1_0_Wij_reg_Dout_6 (.Q (CacheWindow_3__0__6), .QB (
        \$dummy [1556]), .D (CACHE_L0_3_L1_0_Wij_nx272), .CLK (CLK)) ;
    dff CACHE_L0_3_L1_0_Wij_reg_Dout_7 (.Q (CacheWindow_3__0__7), .QB (
        \$dummy [1557]), .D (CACHE_L0_3_L1_0_Wij_nx282), .CLK (CLK)) ;
    buf02 CACHE_L0_3_L1_0_Wij_ix330 (.Y (CACHE_L0_3_L1_0_Wij_nx331), .A (
          CACHE_EN_dup_1414)) ;
    buf02 CACHE_L0_3_L1_0_Wij_ix332 (.Y (CACHE_L0_3_L1_0_Wij_nx333), .A (
          CACHE_EN_dup_1414)) ;
    dff CACHE_L0_3_L1_1_Fij_reg_Dout_0 (.Q (CacheFilter_3__1__0), .QB (
        \$dummy [1558]), .D (CACHE_L0_3_L1_1_Fij_nx212), .CLK (CLK)) ;
    nor02_2x CACHE_L0_3_L1_1_Fij_ix297 (.Y (CACHE_L0_3_L1_1_Fij_nx296), .A0 (
             nx8421), .A1 (CACHE_L0_3_L1_1_Fij_nx331)) ;
    dff CACHE_L0_3_L1_1_Fij_reg_Dout_1 (.Q (CacheFilter_3__1__1), .QB (
        \$dummy [1559]), .D (CACHE_L0_3_L1_1_Fij_nx222), .CLK (CLK)) ;
    dff CACHE_L0_3_L1_1_Fij_reg_Dout_2 (.Q (CacheFilter_3__1__2), .QB (
        \$dummy [1560]), .D (CACHE_L0_3_L1_1_Fij_nx232), .CLK (CLK)) ;
    dff CACHE_L0_3_L1_1_Fij_reg_Dout_3 (.Q (CacheFilter_3__1__3), .QB (
        \$dummy [1561]), .D (CACHE_L0_3_L1_1_Fij_nx242), .CLK (CLK)) ;
    dff CACHE_L0_3_L1_1_Fij_reg_Dout_4 (.Q (CacheFilter_3__1__4), .QB (
        \$dummy [1562]), .D (CACHE_L0_3_L1_1_Fij_nx252), .CLK (CLK)) ;
    dff CACHE_L0_3_L1_1_Fij_reg_Dout_5 (.Q (CacheFilter_3__1__5), .QB (
        \$dummy [1563]), .D (CACHE_L0_3_L1_1_Fij_nx262), .CLK (CLK)) ;
    dff CACHE_L0_3_L1_1_Fij_reg_Dout_6 (.Q (CacheFilter_3__1__6), .QB (
        \$dummy [1564]), .D (CACHE_L0_3_L1_1_Fij_nx272), .CLK (CLK)) ;
    dff CACHE_L0_3_L1_1_Fij_reg_Dout_7 (.Q (CacheFilter_3__1__7), .QB (
        \$dummy [1565]), .D (CACHE_L0_3_L1_1_Fij_nx282), .CLK (CLK)) ;
    buf02 CACHE_L0_3_L1_1_Fij_ix330 (.Y (CACHE_L0_3_L1_1_Fij_nx331), .A (
          CACHE_EN_dup_1403)) ;
    buf02 CACHE_L0_3_L1_1_Fij_ix332 (.Y (CACHE_L0_3_L1_1_Fij_nx333), .A (
          CACHE_EN_dup_1403)) ;
    dff CACHE_L0_3_L1_1_Wij_reg_Dout_0 (.Q (CacheWindow_3__1__0), .QB (
        \$dummy [1566]), .D (CACHE_L0_3_L1_1_Wij_nx212), .CLK (CLK)) ;
    nor02_2x CACHE_L0_3_L1_1_Wij_ix297 (.Y (CACHE_L0_3_L1_1_Wij_nx296), .A0 (
             nx8421), .A1 (CACHE_L0_3_L1_1_Wij_nx331)) ;
    dff CACHE_L0_3_L1_1_Wij_reg_Dout_1 (.Q (CacheWindow_3__1__1), .QB (
        \$dummy [1567]), .D (CACHE_L0_3_L1_1_Wij_nx222), .CLK (CLK)) ;
    dff CACHE_L0_3_L1_1_Wij_reg_Dout_2 (.Q (CacheWindow_3__1__2), .QB (
        \$dummy [1568]), .D (CACHE_L0_3_L1_1_Wij_nx232), .CLK (CLK)) ;
    dff CACHE_L0_3_L1_1_Wij_reg_Dout_3 (.Q (CacheWindow_3__1__3), .QB (
        \$dummy [1569]), .D (CACHE_L0_3_L1_1_Wij_nx242), .CLK (CLK)) ;
    dff CACHE_L0_3_L1_1_Wij_reg_Dout_4 (.Q (CacheWindow_3__1__4), .QB (
        \$dummy [1570]), .D (CACHE_L0_3_L1_1_Wij_nx252), .CLK (CLK)) ;
    dff CACHE_L0_3_L1_1_Wij_reg_Dout_5 (.Q (CacheWindow_3__1__5), .QB (
        \$dummy [1571]), .D (CACHE_L0_3_L1_1_Wij_nx262), .CLK (CLK)) ;
    dff CACHE_L0_3_L1_1_Wij_reg_Dout_6 (.Q (CacheWindow_3__1__6), .QB (
        \$dummy [1572]), .D (CACHE_L0_3_L1_1_Wij_nx272), .CLK (CLK)) ;
    dff CACHE_L0_3_L1_1_Wij_reg_Dout_7 (.Q (CacheWindow_3__1__7), .QB (
        \$dummy [1573]), .D (CACHE_L0_3_L1_1_Wij_nx282), .CLK (CLK)) ;
    buf02 CACHE_L0_3_L1_1_Wij_ix330 (.Y (CACHE_L0_3_L1_1_Wij_nx331), .A (
          CACHE_EN_dup_1414)) ;
    buf02 CACHE_L0_3_L1_1_Wij_ix332 (.Y (CACHE_L0_3_L1_1_Wij_nx333), .A (
          CACHE_EN_dup_1414)) ;
    dff CACHE_L0_3_L1_2_Fij_reg_Dout_0 (.Q (CacheFilter_3__2__0), .QB (
        \$dummy [1574]), .D (CACHE_L0_3_L1_2_Fij_nx212), .CLK (CLK)) ;
    nor02_2x CACHE_L0_3_L1_2_Fij_ix297 (.Y (CACHE_L0_3_L1_2_Fij_nx296), .A0 (
             nx8425), .A1 (CACHE_L0_3_L1_2_Fij_nx331)) ;
    dff CACHE_L0_3_L1_2_Fij_reg_Dout_1 (.Q (CacheFilter_3__2__1), .QB (
        \$dummy [1575]), .D (CACHE_L0_3_L1_2_Fij_nx222), .CLK (CLK)) ;
    dff CACHE_L0_3_L1_2_Fij_reg_Dout_2 (.Q (CacheFilter_3__2__2), .QB (
        \$dummy [1576]), .D (CACHE_L0_3_L1_2_Fij_nx232), .CLK (CLK)) ;
    dff CACHE_L0_3_L1_2_Fij_reg_Dout_3 (.Q (CacheFilter_3__2__3), .QB (
        \$dummy [1577]), .D (CACHE_L0_3_L1_2_Fij_nx242), .CLK (CLK)) ;
    dff CACHE_L0_3_L1_2_Fij_reg_Dout_4 (.Q (CacheFilter_3__2__4), .QB (
        \$dummy [1578]), .D (CACHE_L0_3_L1_2_Fij_nx252), .CLK (CLK)) ;
    dff CACHE_L0_3_L1_2_Fij_reg_Dout_5 (.Q (CacheFilter_3__2__5), .QB (
        \$dummy [1579]), .D (CACHE_L0_3_L1_2_Fij_nx262), .CLK (CLK)) ;
    dff CACHE_L0_3_L1_2_Fij_reg_Dout_6 (.Q (CacheFilter_3__2__6), .QB (
        \$dummy [1580]), .D (CACHE_L0_3_L1_2_Fij_nx272), .CLK (CLK)) ;
    dff CACHE_L0_3_L1_2_Fij_reg_Dout_7 (.Q (CacheFilter_3__2__7), .QB (
        \$dummy [1581]), .D (CACHE_L0_3_L1_2_Fij_nx282), .CLK (CLK)) ;
    buf02 CACHE_L0_3_L1_2_Fij_ix330 (.Y (CACHE_L0_3_L1_2_Fij_nx331), .A (
          CACHE_EN_dup_1403)) ;
    buf02 CACHE_L0_3_L1_2_Fij_ix332 (.Y (CACHE_L0_3_L1_2_Fij_nx333), .A (
          CACHE_EN_dup_1403)) ;
    dff CACHE_L0_3_L1_2_Wij_reg_Dout_0 (.Q (CacheWindow_3__2__0), .QB (
        \$dummy [1582]), .D (CACHE_L0_3_L1_2_Wij_nx212), .CLK (CLK)) ;
    nor02_2x CACHE_L0_3_L1_2_Wij_ix297 (.Y (CACHE_L0_3_L1_2_Wij_nx296), .A0 (
             nx8425), .A1 (CACHE_L0_3_L1_2_Wij_nx331)) ;
    dff CACHE_L0_3_L1_2_Wij_reg_Dout_1 (.Q (CacheWindow_3__2__1), .QB (
        \$dummy [1583]), .D (CACHE_L0_3_L1_2_Wij_nx222), .CLK (CLK)) ;
    dff CACHE_L0_3_L1_2_Wij_reg_Dout_2 (.Q (CacheWindow_3__2__2), .QB (
        \$dummy [1584]), .D (CACHE_L0_3_L1_2_Wij_nx232), .CLK (CLK)) ;
    dff CACHE_L0_3_L1_2_Wij_reg_Dout_3 (.Q (CacheWindow_3__2__3), .QB (
        \$dummy [1585]), .D (CACHE_L0_3_L1_2_Wij_nx242), .CLK (CLK)) ;
    dff CACHE_L0_3_L1_2_Wij_reg_Dout_4 (.Q (CacheWindow_3__2__4), .QB (
        \$dummy [1586]), .D (CACHE_L0_3_L1_2_Wij_nx252), .CLK (CLK)) ;
    dff CACHE_L0_3_L1_2_Wij_reg_Dout_5 (.Q (CacheWindow_3__2__5), .QB (
        \$dummy [1587]), .D (CACHE_L0_3_L1_2_Wij_nx262), .CLK (CLK)) ;
    dff CACHE_L0_3_L1_2_Wij_reg_Dout_6 (.Q (CacheWindow_3__2__6), .QB (
        \$dummy [1588]), .D (CACHE_L0_3_L1_2_Wij_nx272), .CLK (CLK)) ;
    dff CACHE_L0_3_L1_2_Wij_reg_Dout_7 (.Q (CacheWindow_3__2__7), .QB (
        \$dummy [1589]), .D (CACHE_L0_3_L1_2_Wij_nx282), .CLK (CLK)) ;
    buf02 CACHE_L0_3_L1_2_Wij_ix330 (.Y (CACHE_L0_3_L1_2_Wij_nx331), .A (
          CACHE_EN_dup_1414)) ;
    buf02 CACHE_L0_3_L1_2_Wij_ix332 (.Y (CACHE_L0_3_L1_2_Wij_nx333), .A (
          CACHE_EN_dup_1414)) ;
    dff CACHE_L0_3_L1_3_Fij_reg_Dout_0 (.Q (CacheFilter_3__3__0), .QB (
        \$dummy [1590]), .D (CACHE_L0_3_L1_3_Fij_nx212), .CLK (CLK)) ;
    nor02_2x CACHE_L0_3_L1_3_Fij_ix297 (.Y (CACHE_L0_3_L1_3_Fij_nx296), .A0 (
             nx8429), .A1 (CACHE_L0_3_L1_3_Fij_nx331)) ;
    dff CACHE_L0_3_L1_3_Fij_reg_Dout_1 (.Q (CacheFilter_3__3__1), .QB (
        \$dummy [1591]), .D (CACHE_L0_3_L1_3_Fij_nx222), .CLK (CLK)) ;
    dff CACHE_L0_3_L1_3_Fij_reg_Dout_2 (.Q (CacheFilter_3__3__2), .QB (
        \$dummy [1592]), .D (CACHE_L0_3_L1_3_Fij_nx232), .CLK (CLK)) ;
    dff CACHE_L0_3_L1_3_Fij_reg_Dout_3 (.Q (CacheFilter_3__3__3), .QB (
        \$dummy [1593]), .D (CACHE_L0_3_L1_3_Fij_nx242), .CLK (CLK)) ;
    dff CACHE_L0_3_L1_3_Fij_reg_Dout_4 (.Q (CacheFilter_3__3__4), .QB (
        \$dummy [1594]), .D (CACHE_L0_3_L1_3_Fij_nx252), .CLK (CLK)) ;
    dff CACHE_L0_3_L1_3_Fij_reg_Dout_5 (.Q (CacheFilter_3__3__5), .QB (
        \$dummy [1595]), .D (CACHE_L0_3_L1_3_Fij_nx262), .CLK (CLK)) ;
    dff CACHE_L0_3_L1_3_Fij_reg_Dout_6 (.Q (CacheFilter_3__3__6), .QB (
        \$dummy [1596]), .D (CACHE_L0_3_L1_3_Fij_nx272), .CLK (CLK)) ;
    dff CACHE_L0_3_L1_3_Fij_reg_Dout_7 (.Q (CacheFilter_3__3__7), .QB (
        \$dummy [1597]), .D (CACHE_L0_3_L1_3_Fij_nx282), .CLK (CLK)) ;
    buf02 CACHE_L0_3_L1_3_Fij_ix330 (.Y (CACHE_L0_3_L1_3_Fij_nx331), .A (
          CACHE_EN_dup_1359)) ;
    buf02 CACHE_L0_3_L1_3_Fij_ix332 (.Y (CACHE_L0_3_L1_3_Fij_nx333), .A (
          CACHE_EN_dup_1359)) ;
    dff CACHE_L0_3_L1_3_Wij_reg_Dout_0 (.Q (CacheWindow_3__3__0), .QB (
        \$dummy [1598]), .D (CACHE_L0_3_L1_3_Wij_nx212), .CLK (CLK)) ;
    nor02_2x CACHE_L0_3_L1_3_Wij_ix297 (.Y (CACHE_L0_3_L1_3_Wij_nx296), .A0 (
             nx8429), .A1 (CACHE_L0_3_L1_3_Wij_nx331)) ;
    dff CACHE_L0_3_L1_3_Wij_reg_Dout_1 (.Q (CacheWindow_3__3__1), .QB (
        \$dummy [1599]), .D (CACHE_L0_3_L1_3_Wij_nx222), .CLK (CLK)) ;
    dff CACHE_L0_3_L1_3_Wij_reg_Dout_2 (.Q (CacheWindow_3__3__2), .QB (
        \$dummy [1600]), .D (CACHE_L0_3_L1_3_Wij_nx232), .CLK (CLK)) ;
    dff CACHE_L0_3_L1_3_Wij_reg_Dout_3 (.Q (CacheWindow_3__3__3), .QB (
        \$dummy [1601]), .D (CACHE_L0_3_L1_3_Wij_nx242), .CLK (CLK)) ;
    dff CACHE_L0_3_L1_3_Wij_reg_Dout_4 (.Q (CacheWindow_3__3__4), .QB (
        \$dummy [1602]), .D (CACHE_L0_3_L1_3_Wij_nx252), .CLK (CLK)) ;
    dff CACHE_L0_3_L1_3_Wij_reg_Dout_5 (.Q (CacheWindow_3__3__5), .QB (
        \$dummy [1603]), .D (CACHE_L0_3_L1_3_Wij_nx262), .CLK (CLK)) ;
    dff CACHE_L0_3_L1_3_Wij_reg_Dout_6 (.Q (CacheWindow_3__3__6), .QB (
        \$dummy [1604]), .D (CACHE_L0_3_L1_3_Wij_nx272), .CLK (CLK)) ;
    dff CACHE_L0_3_L1_3_Wij_reg_Dout_7 (.Q (CacheWindow_3__3__7), .QB (
        \$dummy [1605]), .D (CACHE_L0_3_L1_3_Wij_nx282), .CLK (CLK)) ;
    buf02 CACHE_L0_3_L1_3_Wij_ix330 (.Y (CACHE_L0_3_L1_3_Wij_nx331), .A (
          CACHE_EN_dup_1370)) ;
    buf02 CACHE_L0_3_L1_3_Wij_ix332 (.Y (CACHE_L0_3_L1_3_Wij_nx333), .A (
          CACHE_EN_dup_1370)) ;
    dff CACHE_L0_3_L1_4_Fij_reg_Dout_0 (.Q (CacheFilter_3__4__0), .QB (
        \$dummy [1606]), .D (CACHE_L0_3_L1_4_Fij_nx212), .CLK (CLK)) ;
    nor02_2x CACHE_L0_3_L1_4_Fij_ix297 (.Y (CACHE_L0_3_L1_4_Fij_nx296), .A0 (
             nx8433), .A1 (CACHE_L0_3_L1_4_Fij_nx331)) ;
    dff CACHE_L0_3_L1_4_Fij_reg_Dout_1 (.Q (CacheFilter_3__4__1), .QB (
        \$dummy [1607]), .D (CACHE_L0_3_L1_4_Fij_nx222), .CLK (CLK)) ;
    dff CACHE_L0_3_L1_4_Fij_reg_Dout_2 (.Q (CacheFilter_3__4__2), .QB (
        \$dummy [1608]), .D (CACHE_L0_3_L1_4_Fij_nx232), .CLK (CLK)) ;
    dff CACHE_L0_3_L1_4_Fij_reg_Dout_3 (.Q (CacheFilter_3__4__3), .QB (
        \$dummy [1609]), .D (CACHE_L0_3_L1_4_Fij_nx242), .CLK (CLK)) ;
    dff CACHE_L0_3_L1_4_Fij_reg_Dout_4 (.Q (CacheFilter_3__4__4), .QB (
        \$dummy [1610]), .D (CACHE_L0_3_L1_4_Fij_nx252), .CLK (CLK)) ;
    dff CACHE_L0_3_L1_4_Fij_reg_Dout_5 (.Q (CacheFilter_3__4__5), .QB (
        \$dummy [1611]), .D (CACHE_L0_3_L1_4_Fij_nx262), .CLK (CLK)) ;
    dff CACHE_L0_3_L1_4_Fij_reg_Dout_6 (.Q (CacheFilter_3__4__6), .QB (
        \$dummy [1612]), .D (CACHE_L0_3_L1_4_Fij_nx272), .CLK (CLK)) ;
    dff CACHE_L0_3_L1_4_Fij_reg_Dout_7 (.Q (CacheFilter_3__4__7), .QB (
        \$dummy [1613]), .D (CACHE_L0_3_L1_4_Fij_nx282), .CLK (CLK)) ;
    buf02 CACHE_L0_3_L1_4_Fij_ix330 (.Y (CACHE_L0_3_L1_4_Fij_nx331), .A (
          CACHE_EN_dup_1491)) ;
    buf02 CACHE_L0_3_L1_4_Fij_ix332 (.Y (CACHE_L0_3_L1_4_Fij_nx333), .A (
          CACHE_EN_dup_1491)) ;
    dff CACHE_L0_3_L1_4_Wij_reg_Dout_0 (.Q (CacheWindow_3__4__0), .QB (
        \$dummy [1614]), .D (CACHE_L0_3_L1_4_Wij_nx212), .CLK (CLK)) ;
    nor02_2x CACHE_L0_3_L1_4_Wij_ix297 (.Y (CACHE_L0_3_L1_4_Wij_nx296), .A0 (
             nx8433), .A1 (CACHE_L0_3_L1_4_Wij_nx331)) ;
    dff CACHE_L0_3_L1_4_Wij_reg_Dout_1 (.Q (CacheWindow_3__4__1), .QB (
        \$dummy [1615]), .D (CACHE_L0_3_L1_4_Wij_nx222), .CLK (CLK)) ;
    dff CACHE_L0_3_L1_4_Wij_reg_Dout_2 (.Q (CacheWindow_3__4__2), .QB (
        \$dummy [1616]), .D (CACHE_L0_3_L1_4_Wij_nx232), .CLK (CLK)) ;
    dff CACHE_L0_3_L1_4_Wij_reg_Dout_3 (.Q (CacheWindow_3__4__3), .QB (
        \$dummy [1617]), .D (CACHE_L0_3_L1_4_Wij_nx242), .CLK (CLK)) ;
    dff CACHE_L0_3_L1_4_Wij_reg_Dout_4 (.Q (CacheWindow_3__4__4), .QB (
        \$dummy [1618]), .D (CACHE_L0_3_L1_4_Wij_nx252), .CLK (CLK)) ;
    dff CACHE_L0_3_L1_4_Wij_reg_Dout_5 (.Q (CacheWindow_3__4__5), .QB (
        \$dummy [1619]), .D (CACHE_L0_3_L1_4_Wij_nx262), .CLK (CLK)) ;
    dff CACHE_L0_3_L1_4_Wij_reg_Dout_6 (.Q (CacheWindow_3__4__6), .QB (
        \$dummy [1620]), .D (CACHE_L0_3_L1_4_Wij_nx272), .CLK (CLK)) ;
    dff CACHE_L0_3_L1_4_Wij_reg_Dout_7 (.Q (CacheWindow_3__4__7), .QB (
        \$dummy [1621]), .D (CACHE_L0_3_L1_4_Wij_nx282), .CLK (CLK)) ;
    buf02 CACHE_L0_3_L1_4_Wij_ix330 (.Y (CACHE_L0_3_L1_4_Wij_nx331), .A (
          CACHE_EN_dup_1502)) ;
    buf02 CACHE_L0_3_L1_4_Wij_ix332 (.Y (CACHE_L0_3_L1_4_Wij_nx333), .A (
          CACHE_EN_dup_1502)) ;
    dff CACHE_L0_4_L1_0_Fij_reg_Dout_0 (.Q (CacheFilter_4__0__0), .QB (
        \$dummy [1622]), .D (CACHE_L0_4_L1_0_Fij_nx212), .CLK (CLK)) ;
    nor02_2x CACHE_L0_4_L1_0_Fij_ix297 (.Y (CACHE_L0_4_L1_0_Fij_nx296), .A0 (
             nx8437), .A1 (CACHE_L0_4_L1_0_Fij_nx331)) ;
    dff CACHE_L0_4_L1_0_Fij_reg_Dout_1 (.Q (CacheFilter_4__0__1), .QB (
        \$dummy [1623]), .D (CACHE_L0_4_L1_0_Fij_nx222), .CLK (CLK)) ;
    dff CACHE_L0_4_L1_0_Fij_reg_Dout_2 (.Q (CacheFilter_4__0__2), .QB (
        \$dummy [1624]), .D (CACHE_L0_4_L1_0_Fij_nx232), .CLK (CLK)) ;
    dff CACHE_L0_4_L1_0_Fij_reg_Dout_3 (.Q (CacheFilter_4__0__3), .QB (
        \$dummy [1625]), .D (CACHE_L0_4_L1_0_Fij_nx242), .CLK (CLK)) ;
    dff CACHE_L0_4_L1_0_Fij_reg_Dout_4 (.Q (CacheFilter_4__0__4), .QB (
        \$dummy [1626]), .D (CACHE_L0_4_L1_0_Fij_nx252), .CLK (CLK)) ;
    dff CACHE_L0_4_L1_0_Fij_reg_Dout_5 (.Q (CacheFilter_4__0__5), .QB (
        \$dummy [1627]), .D (CACHE_L0_4_L1_0_Fij_nx262), .CLK (CLK)) ;
    dff CACHE_L0_4_L1_0_Fij_reg_Dout_6 (.Q (CacheFilter_4__0__6), .QB (
        \$dummy [1628]), .D (CACHE_L0_4_L1_0_Fij_nx272), .CLK (CLK)) ;
    dff CACHE_L0_4_L1_0_Fij_reg_Dout_7 (.Q (CacheFilter_4__0__7), .QB (
        \$dummy [1629]), .D (CACHE_L0_4_L1_0_Fij_nx282), .CLK (CLK)) ;
    buf02 CACHE_L0_4_L1_0_Fij_ix330 (.Y (CACHE_L0_4_L1_0_Fij_nx331), .A (
          CACHE_EN_dup_1513)) ;
    buf02 CACHE_L0_4_L1_0_Fij_ix332 (.Y (CACHE_L0_4_L1_0_Fij_nx333), .A (
          CACHE_EN_dup_1513)) ;
    dff CACHE_L0_4_L1_0_Wij_reg_Dout_0 (.Q (CacheWindow_4__0__0), .QB (
        \$dummy [1630]), .D (CACHE_L0_4_L1_0_Wij_nx212), .CLK (CLK)) ;
    nor02_2x CACHE_L0_4_L1_0_Wij_ix297 (.Y (CACHE_L0_4_L1_0_Wij_nx296), .A0 (
             nx8437), .A1 (CACHE_L0_4_L1_0_Wij_nx331)) ;
    dff CACHE_L0_4_L1_0_Wij_reg_Dout_1 (.Q (CacheWindow_4__0__1), .QB (
        \$dummy [1631]), .D (CACHE_L0_4_L1_0_Wij_nx222), .CLK (CLK)) ;
    dff CACHE_L0_4_L1_0_Wij_reg_Dout_2 (.Q (CacheWindow_4__0__2), .QB (
        \$dummy [1632]), .D (CACHE_L0_4_L1_0_Wij_nx232), .CLK (CLK)) ;
    dff CACHE_L0_4_L1_0_Wij_reg_Dout_3 (.Q (CacheWindow_4__0__3), .QB (
        \$dummy [1633]), .D (CACHE_L0_4_L1_0_Wij_nx242), .CLK (CLK)) ;
    dff CACHE_L0_4_L1_0_Wij_reg_Dout_4 (.Q (CacheWindow_4__0__4), .QB (
        \$dummy [1634]), .D (CACHE_L0_4_L1_0_Wij_nx252), .CLK (CLK)) ;
    dff CACHE_L0_4_L1_0_Wij_reg_Dout_5 (.Q (CacheWindow_4__0__5), .QB (
        \$dummy [1635]), .D (CACHE_L0_4_L1_0_Wij_nx262), .CLK (CLK)) ;
    dff CACHE_L0_4_L1_0_Wij_reg_Dout_6 (.Q (CacheWindow_4__0__6), .QB (
        \$dummy [1636]), .D (CACHE_L0_4_L1_0_Wij_nx272), .CLK (CLK)) ;
    dff CACHE_L0_4_L1_0_Wij_reg_Dout_7 (.Q (CacheWindow_4__0__7), .QB (
        \$dummy [1637]), .D (CACHE_L0_4_L1_0_Wij_nx282), .CLK (CLK)) ;
    buf02 CACHE_L0_4_L1_0_Wij_ix330 (.Y (CACHE_L0_4_L1_0_Wij_nx331), .A (
          CACHE_EN_dup_1524)) ;
    buf02 CACHE_L0_4_L1_0_Wij_ix332 (.Y (CACHE_L0_4_L1_0_Wij_nx333), .A (
          CACHE_EN_dup_1524)) ;
    dff CACHE_L0_4_L1_1_Fij_reg_Dout_0 (.Q (CacheFilter_4__1__0), .QB (
        \$dummy [1638]), .D (CACHE_L0_4_L1_1_Fij_nx212), .CLK (CLK)) ;
    nor02_2x CACHE_L0_4_L1_1_Fij_ix297 (.Y (CACHE_L0_4_L1_1_Fij_nx296), .A0 (
             nx8441), .A1 (CACHE_L0_4_L1_1_Fij_nx331)) ;
    dff CACHE_L0_4_L1_1_Fij_reg_Dout_1 (.Q (CacheFilter_4__1__1), .QB (
        \$dummy [1639]), .D (CACHE_L0_4_L1_1_Fij_nx222), .CLK (CLK)) ;
    dff CACHE_L0_4_L1_1_Fij_reg_Dout_2 (.Q (CacheFilter_4__1__2), .QB (
        \$dummy [1640]), .D (CACHE_L0_4_L1_1_Fij_nx232), .CLK (CLK)) ;
    dff CACHE_L0_4_L1_1_Fij_reg_Dout_3 (.Q (CacheFilter_4__1__3), .QB (
        \$dummy [1641]), .D (CACHE_L0_4_L1_1_Fij_nx242), .CLK (CLK)) ;
    dff CACHE_L0_4_L1_1_Fij_reg_Dout_4 (.Q (CacheFilter_4__1__4), .QB (
        \$dummy [1642]), .D (CACHE_L0_4_L1_1_Fij_nx252), .CLK (CLK)) ;
    dff CACHE_L0_4_L1_1_Fij_reg_Dout_5 (.Q (CacheFilter_4__1__5), .QB (
        \$dummy [1643]), .D (CACHE_L0_4_L1_1_Fij_nx262), .CLK (CLK)) ;
    dff CACHE_L0_4_L1_1_Fij_reg_Dout_6 (.Q (CacheFilter_4__1__6), .QB (
        \$dummy [1644]), .D (CACHE_L0_4_L1_1_Fij_nx272), .CLK (CLK)) ;
    dff CACHE_L0_4_L1_1_Fij_reg_Dout_7 (.Q (CacheFilter_4__1__7), .QB (
        \$dummy [1645]), .D (CACHE_L0_4_L1_1_Fij_nx282), .CLK (CLK)) ;
    buf02 CACHE_L0_4_L1_1_Fij_ix330 (.Y (CACHE_L0_4_L1_1_Fij_nx331), .A (
          CACHE_EN_dup_1513)) ;
    buf02 CACHE_L0_4_L1_1_Fij_ix332 (.Y (CACHE_L0_4_L1_1_Fij_nx333), .A (
          CACHE_EN_dup_1513)) ;
    dff CACHE_L0_4_L1_1_Wij_reg_Dout_0 (.Q (CacheWindow_4__1__0), .QB (
        \$dummy [1646]), .D (CACHE_L0_4_L1_1_Wij_nx212), .CLK (CLK)) ;
    nor02_2x CACHE_L0_4_L1_1_Wij_ix297 (.Y (CACHE_L0_4_L1_1_Wij_nx296), .A0 (
             nx8441), .A1 (CACHE_L0_4_L1_1_Wij_nx331)) ;
    dff CACHE_L0_4_L1_1_Wij_reg_Dout_1 (.Q (CacheWindow_4__1__1), .QB (
        \$dummy [1647]), .D (CACHE_L0_4_L1_1_Wij_nx222), .CLK (CLK)) ;
    dff CACHE_L0_4_L1_1_Wij_reg_Dout_2 (.Q (CacheWindow_4__1__2), .QB (
        \$dummy [1648]), .D (CACHE_L0_4_L1_1_Wij_nx232), .CLK (CLK)) ;
    dff CACHE_L0_4_L1_1_Wij_reg_Dout_3 (.Q (CacheWindow_4__1__3), .QB (
        \$dummy [1649]), .D (CACHE_L0_4_L1_1_Wij_nx242), .CLK (CLK)) ;
    dff CACHE_L0_4_L1_1_Wij_reg_Dout_4 (.Q (CacheWindow_4__1__4), .QB (
        \$dummy [1650]), .D (CACHE_L0_4_L1_1_Wij_nx252), .CLK (CLK)) ;
    dff CACHE_L0_4_L1_1_Wij_reg_Dout_5 (.Q (CacheWindow_4__1__5), .QB (
        \$dummy [1651]), .D (CACHE_L0_4_L1_1_Wij_nx262), .CLK (CLK)) ;
    dff CACHE_L0_4_L1_1_Wij_reg_Dout_6 (.Q (CacheWindow_4__1__6), .QB (
        \$dummy [1652]), .D (CACHE_L0_4_L1_1_Wij_nx272), .CLK (CLK)) ;
    dff CACHE_L0_4_L1_1_Wij_reg_Dout_7 (.Q (CacheWindow_4__1__7), .QB (
        \$dummy [1653]), .D (CACHE_L0_4_L1_1_Wij_nx282), .CLK (CLK)) ;
    buf02 CACHE_L0_4_L1_1_Wij_ix330 (.Y (CACHE_L0_4_L1_1_Wij_nx331), .A (
          CACHE_EN_dup_1524)) ;
    buf02 CACHE_L0_4_L1_1_Wij_ix332 (.Y (CACHE_L0_4_L1_1_Wij_nx333), .A (
          CACHE_EN_dup_1524)) ;
    dff CACHE_L0_4_L1_2_Fij_reg_Dout_0 (.Q (CacheFilter_4__2__0), .QB (
        \$dummy [1654]), .D (CACHE_L0_4_L1_2_Fij_nx212), .CLK (CLK)) ;
    nor02_2x CACHE_L0_4_L1_2_Fij_ix297 (.Y (CACHE_L0_4_L1_2_Fij_nx296), .A0 (
             nx8445), .A1 (CACHE_L0_4_L1_2_Fij_nx331)) ;
    dff CACHE_L0_4_L1_2_Fij_reg_Dout_1 (.Q (CacheFilter_4__2__1), .QB (
        \$dummy [1655]), .D (CACHE_L0_4_L1_2_Fij_nx222), .CLK (CLK)) ;
    dff CACHE_L0_4_L1_2_Fij_reg_Dout_2 (.Q (CacheFilter_4__2__2), .QB (
        \$dummy [1656]), .D (CACHE_L0_4_L1_2_Fij_nx232), .CLK (CLK)) ;
    dff CACHE_L0_4_L1_2_Fij_reg_Dout_3 (.Q (CacheFilter_4__2__3), .QB (
        \$dummy [1657]), .D (CACHE_L0_4_L1_2_Fij_nx242), .CLK (CLK)) ;
    dff CACHE_L0_4_L1_2_Fij_reg_Dout_4 (.Q (CacheFilter_4__2__4), .QB (
        \$dummy [1658]), .D (CACHE_L0_4_L1_2_Fij_nx252), .CLK (CLK)) ;
    dff CACHE_L0_4_L1_2_Fij_reg_Dout_5 (.Q (CacheFilter_4__2__5), .QB (
        \$dummy [1659]), .D (CACHE_L0_4_L1_2_Fij_nx262), .CLK (CLK)) ;
    dff CACHE_L0_4_L1_2_Fij_reg_Dout_6 (.Q (CacheFilter_4__2__6), .QB (
        \$dummy [1660]), .D (CACHE_L0_4_L1_2_Fij_nx272), .CLK (CLK)) ;
    dff CACHE_L0_4_L1_2_Fij_reg_Dout_7 (.Q (CacheFilter_4__2__7), .QB (
        \$dummy [1661]), .D (CACHE_L0_4_L1_2_Fij_nx282), .CLK (CLK)) ;
    buf02 CACHE_L0_4_L1_2_Fij_ix330 (.Y (CACHE_L0_4_L1_2_Fij_nx331), .A (
          CACHE_EN_dup_1513)) ;
    buf02 CACHE_L0_4_L1_2_Fij_ix332 (.Y (CACHE_L0_4_L1_2_Fij_nx333), .A (
          CACHE_EN_dup_1513)) ;
    dff CACHE_L0_4_L1_2_Wij_reg_Dout_0 (.Q (CacheWindow_4__2__0), .QB (
        \$dummy [1662]), .D (CACHE_L0_4_L1_2_Wij_nx212), .CLK (CLK)) ;
    nor02_2x CACHE_L0_4_L1_2_Wij_ix297 (.Y (CACHE_L0_4_L1_2_Wij_nx296), .A0 (
             nx8445), .A1 (CACHE_L0_4_L1_2_Wij_nx331)) ;
    dff CACHE_L0_4_L1_2_Wij_reg_Dout_1 (.Q (CacheWindow_4__2__1), .QB (
        \$dummy [1663]), .D (CACHE_L0_4_L1_2_Wij_nx222), .CLK (CLK)) ;
    dff CACHE_L0_4_L1_2_Wij_reg_Dout_2 (.Q (CacheWindow_4__2__2), .QB (
        \$dummy [1664]), .D (CACHE_L0_4_L1_2_Wij_nx232), .CLK (CLK)) ;
    dff CACHE_L0_4_L1_2_Wij_reg_Dout_3 (.Q (CacheWindow_4__2__3), .QB (
        \$dummy [1665]), .D (CACHE_L0_4_L1_2_Wij_nx242), .CLK (CLK)) ;
    dff CACHE_L0_4_L1_2_Wij_reg_Dout_4 (.Q (CacheWindow_4__2__4), .QB (
        \$dummy [1666]), .D (CACHE_L0_4_L1_2_Wij_nx252), .CLK (CLK)) ;
    dff CACHE_L0_4_L1_2_Wij_reg_Dout_5 (.Q (CacheWindow_4__2__5), .QB (
        \$dummy [1667]), .D (CACHE_L0_4_L1_2_Wij_nx262), .CLK (CLK)) ;
    dff CACHE_L0_4_L1_2_Wij_reg_Dout_6 (.Q (CacheWindow_4__2__6), .QB (
        \$dummy [1668]), .D (CACHE_L0_4_L1_2_Wij_nx272), .CLK (CLK)) ;
    dff CACHE_L0_4_L1_2_Wij_reg_Dout_7 (.Q (CacheWindow_4__2__7), .QB (
        \$dummy [1669]), .D (CACHE_L0_4_L1_2_Wij_nx282), .CLK (CLK)) ;
    buf02 CACHE_L0_4_L1_2_Wij_ix330 (.Y (CACHE_L0_4_L1_2_Wij_nx331), .A (
          CACHE_EN_dup_1524)) ;
    buf02 CACHE_L0_4_L1_2_Wij_ix332 (.Y (CACHE_L0_4_L1_2_Wij_nx333), .A (
          CACHE_EN_dup_1524)) ;
    dff CACHE_L0_4_L1_3_Fij_reg_Dout_0 (.Q (CacheFilter_4__3__0), .QB (
        \$dummy [1670]), .D (CACHE_L0_4_L1_3_Fij_nx212), .CLK (CLK)) ;
    nor02_2x CACHE_L0_4_L1_3_Fij_ix297 (.Y (CACHE_L0_4_L1_3_Fij_nx296), .A0 (
             nx8449), .A1 (CACHE_L0_4_L1_3_Fij_nx331)) ;
    dff CACHE_L0_4_L1_3_Fij_reg_Dout_1 (.Q (CacheFilter_4__3__1), .QB (
        \$dummy [1671]), .D (CACHE_L0_4_L1_3_Fij_nx222), .CLK (CLK)) ;
    dff CACHE_L0_4_L1_3_Fij_reg_Dout_2 (.Q (CacheFilter_4__3__2), .QB (
        \$dummy [1672]), .D (CACHE_L0_4_L1_3_Fij_nx232), .CLK (CLK)) ;
    dff CACHE_L0_4_L1_3_Fij_reg_Dout_3 (.Q (CacheFilter_4__3__3), .QB (
        \$dummy [1673]), .D (CACHE_L0_4_L1_3_Fij_nx242), .CLK (CLK)) ;
    dff CACHE_L0_4_L1_3_Fij_reg_Dout_4 (.Q (CacheFilter_4__3__4), .QB (
        \$dummy [1674]), .D (CACHE_L0_4_L1_3_Fij_nx252), .CLK (CLK)) ;
    dff CACHE_L0_4_L1_3_Fij_reg_Dout_5 (.Q (CacheFilter_4__3__5), .QB (
        \$dummy [1675]), .D (CACHE_L0_4_L1_3_Fij_nx262), .CLK (CLK)) ;
    dff CACHE_L0_4_L1_3_Fij_reg_Dout_6 (.Q (CacheFilter_4__3__6), .QB (
        \$dummy [1676]), .D (CACHE_L0_4_L1_3_Fij_nx272), .CLK (CLK)) ;
    dff CACHE_L0_4_L1_3_Fij_reg_Dout_7 (.Q (CacheFilter_4__3__7), .QB (
        \$dummy [1677]), .D (CACHE_L0_4_L1_3_Fij_nx282), .CLK (CLK)) ;
    buf02 CACHE_L0_4_L1_3_Fij_ix330 (.Y (CACHE_L0_4_L1_3_Fij_nx331), .A (
          CACHE_EN_dup_1491)) ;
    buf02 CACHE_L0_4_L1_3_Fij_ix332 (.Y (CACHE_L0_4_L1_3_Fij_nx333), .A (
          CACHE_EN_dup_1491)) ;
    dff CACHE_L0_4_L1_3_Wij_reg_Dout_0 (.Q (CacheWindow_4__3__0), .QB (
        \$dummy [1678]), .D (CACHE_L0_4_L1_3_Wij_nx212), .CLK (CLK)) ;
    nor02_2x CACHE_L0_4_L1_3_Wij_ix297 (.Y (CACHE_L0_4_L1_3_Wij_nx296), .A0 (
             nx8449), .A1 (CACHE_L0_4_L1_3_Wij_nx331)) ;
    dff CACHE_L0_4_L1_3_Wij_reg_Dout_1 (.Q (CacheWindow_4__3__1), .QB (
        \$dummy [1679]), .D (CACHE_L0_4_L1_3_Wij_nx222), .CLK (CLK)) ;
    dff CACHE_L0_4_L1_3_Wij_reg_Dout_2 (.Q (CacheWindow_4__3__2), .QB (
        \$dummy [1680]), .D (CACHE_L0_4_L1_3_Wij_nx232), .CLK (CLK)) ;
    dff CACHE_L0_4_L1_3_Wij_reg_Dout_3 (.Q (CacheWindow_4__3__3), .QB (
        \$dummy [1681]), .D (CACHE_L0_4_L1_3_Wij_nx242), .CLK (CLK)) ;
    dff CACHE_L0_4_L1_3_Wij_reg_Dout_4 (.Q (CacheWindow_4__3__4), .QB (
        \$dummy [1682]), .D (CACHE_L0_4_L1_3_Wij_nx252), .CLK (CLK)) ;
    dff CACHE_L0_4_L1_3_Wij_reg_Dout_5 (.Q (CacheWindow_4__3__5), .QB (
        \$dummy [1683]), .D (CACHE_L0_4_L1_3_Wij_nx262), .CLK (CLK)) ;
    dff CACHE_L0_4_L1_3_Wij_reg_Dout_6 (.Q (CacheWindow_4__3__6), .QB (
        \$dummy [1684]), .D (CACHE_L0_4_L1_3_Wij_nx272), .CLK (CLK)) ;
    dff CACHE_L0_4_L1_3_Wij_reg_Dout_7 (.Q (CacheWindow_4__3__7), .QB (
        \$dummy [1685]), .D (CACHE_L0_4_L1_3_Wij_nx282), .CLK (CLK)) ;
    buf02 CACHE_L0_4_L1_3_Wij_ix330 (.Y (CACHE_L0_4_L1_3_Wij_nx331), .A (
          CACHE_EN_dup_1502)) ;
    buf02 CACHE_L0_4_L1_3_Wij_ix332 (.Y (CACHE_L0_4_L1_3_Wij_nx333), .A (
          CACHE_EN_dup_1502)) ;
    dff CACHE_L0_4_L1_4_Fij_reg_Dout_0 (.Q (CacheFilter_4__4__0), .QB (
        \$dummy [1686]), .D (CACHE_L0_4_L1_4_Fij_nx212), .CLK (CLK)) ;
    nor02_2x CACHE_L0_4_L1_4_Fij_ix297 (.Y (CACHE_L0_4_L1_4_Fij_nx296), .A0 (
             nx8453), .A1 (CACHE_L0_4_L1_4_Fij_nx331)) ;
    dff CACHE_L0_4_L1_4_Fij_reg_Dout_1 (.Q (CacheFilter_4__4__1), .QB (
        \$dummy [1687]), .D (CACHE_L0_4_L1_4_Fij_nx222), .CLK (CLK)) ;
    dff CACHE_L0_4_L1_4_Fij_reg_Dout_2 (.Q (CacheFilter_4__4__2), .QB (
        \$dummy [1688]), .D (CACHE_L0_4_L1_4_Fij_nx232), .CLK (CLK)) ;
    dff CACHE_L0_4_L1_4_Fij_reg_Dout_3 (.Q (CacheFilter_4__4__3), .QB (
        \$dummy [1689]), .D (CACHE_L0_4_L1_4_Fij_nx242), .CLK (CLK)) ;
    dff CACHE_L0_4_L1_4_Fij_reg_Dout_4 (.Q (CacheFilter_4__4__4), .QB (
        \$dummy [1690]), .D (CACHE_L0_4_L1_4_Fij_nx252), .CLK (CLK)) ;
    dff CACHE_L0_4_L1_4_Fij_reg_Dout_5 (.Q (CacheFilter_4__4__5), .QB (
        \$dummy [1691]), .D (CACHE_L0_4_L1_4_Fij_nx262), .CLK (CLK)) ;
    dff CACHE_L0_4_L1_4_Fij_reg_Dout_6 (.Q (CacheFilter_4__4__6), .QB (
        \$dummy [1692]), .D (CACHE_L0_4_L1_4_Fij_nx272), .CLK (CLK)) ;
    dff CACHE_L0_4_L1_4_Fij_reg_Dout_7 (.Q (CacheFilter_4__4__7), .QB (
        \$dummy [1693]), .D (CACHE_L0_4_L1_4_Fij_nx282), .CLK (CLK)) ;
    buf02 CACHE_L0_4_L1_4_Fij_ix330 (.Y (CACHE_L0_4_L1_4_Fij_nx331), .A (
          CACHE_EN_dup_1491)) ;
    buf02 CACHE_L0_4_L1_4_Fij_ix332 (.Y (CACHE_L0_4_L1_4_Fij_nx333), .A (
          CACHE_EN_dup_1491)) ;
    dff CACHE_L0_4_L1_4_Wij_reg_Dout_0 (.Q (CacheWindow_4__4__0), .QB (
        \$dummy [1694]), .D (CACHE_L0_4_L1_4_Wij_nx212), .CLK (CLK)) ;
    nor02_2x CACHE_L0_4_L1_4_Wij_ix297 (.Y (CACHE_L0_4_L1_4_Wij_nx296), .A0 (
             nx8453), .A1 (CACHE_L0_4_L1_4_Wij_nx331)) ;
    dff CACHE_L0_4_L1_4_Wij_reg_Dout_1 (.Q (CacheWindow_4__4__1), .QB (
        \$dummy [1695]), .D (CACHE_L0_4_L1_4_Wij_nx222), .CLK (CLK)) ;
    dff CACHE_L0_4_L1_4_Wij_reg_Dout_2 (.Q (CacheWindow_4__4__2), .QB (
        \$dummy [1696]), .D (CACHE_L0_4_L1_4_Wij_nx232), .CLK (CLK)) ;
    dff CACHE_L0_4_L1_4_Wij_reg_Dout_3 (.Q (CacheWindow_4__4__3), .QB (
        \$dummy [1697]), .D (CACHE_L0_4_L1_4_Wij_nx242), .CLK (CLK)) ;
    dff CACHE_L0_4_L1_4_Wij_reg_Dout_4 (.Q (CacheWindow_4__4__4), .QB (
        \$dummy [1698]), .D (CACHE_L0_4_L1_4_Wij_nx252), .CLK (CLK)) ;
    dff CACHE_L0_4_L1_4_Wij_reg_Dout_5 (.Q (CacheWindow_4__4__5), .QB (
        \$dummy [1699]), .D (CACHE_L0_4_L1_4_Wij_nx262), .CLK (CLK)) ;
    dff CACHE_L0_4_L1_4_Wij_reg_Dout_6 (.Q (CacheWindow_4__4__6), .QB (
        \$dummy [1700]), .D (CACHE_L0_4_L1_4_Wij_nx272), .CLK (CLK)) ;
    dff CACHE_L0_4_L1_4_Wij_reg_Dout_7 (.Q (CacheWindow_4__4__7), .QB (
        \$dummy [1701]), .D (CACHE_L0_4_L1_4_Wij_nx282), .CLK (CLK)) ;
    buf02 CACHE_L0_4_L1_4_Wij_ix330 (.Y (CACHE_L0_4_L1_4_Wij_nx331), .A (
          CACHE_EN_dup_1502)) ;
    buf02 CACHE_L0_4_L1_4_Wij_ix332 (.Y (CACHE_L0_4_L1_4_Wij_nx333), .A (
          CACHE_EN_dup_1502)) ;
    oai21 CONTROLLER_ix511 (.Y (CONTROLLER_CntEN), .A0 (CONTROLLER_nx502), .A1 (
          nx619), .B0 (nx621)) ;
    inv01 ix618 (.Y (nx619), .A (MemRD)) ;
    inv01 ix620 (.Y (nx621), .A (CONTROLLER_nx791)) ;
    oai22 CONTROLLER_ix459 (.Y (MemAddr[15]), .A0 (CONTROLLER_nx640), .A1 (
          CONTROLLER_nx811), .B0 (CONTROLLER_nx781), .B1 (CONTROLLER_nx815)) ;
    xnor2 CONTROLLER_ix57 (.Y (CONTROLLER_NxtRow_1), .A0 (CONTROLLER_CurRow_1), 
          .A1 (CONTROLLER_NxtRow_0)) ;
    nand02 CONTROLLER_ix623 (.Y (CONTROLLER_nx622), .A0 (CONTROLLER_CurRow_1), .A1 (
           CONTROLLER_CurRow_0)) ;
    nor02_2x CONTROLLER_ix741 (.Y (CONTROLLER_nx740), .A0 (FilterSize), .A1 (
             CONTROLLER_CurRow_0)) ;
    xnor2 CONTROLLER_ix321 (.Y (CONTROLLER_nx320), .A0 (FilterSize), .A1 (
          CONTROLLER_CurRow_1)) ;
    oai32 CONTROLLER_STATE_ix153 (.Y (CONTROLLER_STATE_nx152), .A0 (nx623), .A1 (
          nx7285), .A2 (nx625), .B0 (CACHE_nx1025), .B1 (nx627)) ;
    inv01 ix622 (.Y (nx623), .A (CONTROLLER_NxtState_0)) ;
    inv02 ix624 (.Y (nx625), .A (CONTROLLER_FilterAddr_17)) ;
    inv02 ix626 (.Y (nx627), .A (CONTROLLER_STATE_nx206)) ;
    oai32 CONTROLLER_STATE_ix163 (.Y (CONTROLLER_STATE_nx162), .A0 (nx629), .A1 (
          nx7285), .A2 (nx625), .B0 (CACHE_nx1033), .B1 (nx627)) ;
    inv01 ix628 (.Y (nx629), .A (CONTROLLER_NxtState_1)) ;
    oai32 CONTROLLER_STATE_ix173 (.Y (CONTROLLER_STATE_nx172), .A0 (nx631), .A1 (
          nx7285), .A2 (nx625), .B0 (nx633), .B1 (nx627)) ;
    inv01 ix630 (.Y (nx631), .A (CONTROLLER_NxtState_2)) ;
    inv01 ix632 (.Y (nx633), .A (MemWR)) ;
    oai32 CONTROLLER_STATE_ix183 (.Y (CONTROLLER_STATE_nx182), .A0 (nx635), .A1 (
          nx7285), .A2 (nx625), .B0 (nx637), .B1 (nx627)) ;
    inv01 ix634 (.Y (nx635), .A (CONTROLLER_NxtState_3)) ;
    inv01 ix636 (.Y (nx637), .A (Calculating)) ;
    oai32 CONTROLLER_STATE_ix193 (.Y (CONTROLLER_STATE_nx192), .A0 (nx639), .A1 (
          nx7285), .A2 (nx625), .B0 (nx641), .B1 (nx627)) ;
    inv01 ix638 (.Y (nx639), .A (CONTROLLER_NxtState_4)) ;
    inv01 ix640 (.Y (nx641), .A (Done)) ;
    oai32 CONTROLLER_ROW_ix213 (.Y (CONTROLLER_ROW_nx212), .A0 (
          CONTROLLER_CurRow_0), .A1 (nx7289), .A2 (nx643), .B0 (
          CONTROLLER_NxtRow_0), .B1 (nx8471)) ;
    inv02 ix642 (.Y (nx643), .A (CONTROLLER_ROW_nx335)) ;
    oai32 CONTROLLER_ROW_ix223 (.Y (CONTROLLER_ROW_nx222), .A0 (nx647), .A1 (
          nx7289), .A2 (nx643), .B0 (CONTROLLER_nx709), .B1 (nx8471)) ;
    inv01 ix646 (.Y (nx647), .A (CONTROLLER_NxtRow_1)) ;
    oai32 CONTROLLER_ROW_ix233 (.Y (CONTROLLER_ROW_nx232), .A0 (nx649), .A1 (
          nx7289), .A2 (nx643), .B0 (CONTROLLER_nx756), .B1 (nx8471)) ;
    inv01 ix648 (.Y (nx649), .A (CONTROLLER_NxtRow_2)) ;
    oai32 CONTROLLER_ROW_ix243 (.Y (CONTROLLER_ROW_nx242), .A0 (nx651), .A1 (
          nx7289), .A2 (nx643), .B0 (CONTROLLER_nx727), .B1 (nx8471)) ;
    inv01 ix650 (.Y (nx651), .A (CONTROLLER_NxtRow_3)) ;
    oai32 CONTROLLER_ROW_ix253 (.Y (CONTROLLER_ROW_nx252), .A0 (nx653), .A1 (
          nx7289), .A2 (nx643), .B0 (CONTROLLER_nx581), .B1 (nx8471)) ;
    inv01 ix652 (.Y (nx653), .A (CONTROLLER_NxtRow_4)) ;
    oai32 CONTROLLER_ROW_ix263 (.Y (CONTROLLER_ROW_nx262), .A0 (nx655), .A1 (
          nx7291), .A2 (nx643), .B0 (CONTROLLER_nx778), .B1 (nx8471)) ;
    inv01 ix654 (.Y (nx655), .A (CONTROLLER_NxtRow_5)) ;
    oai32 CONTROLLER_ROW_ix273 (.Y (CONTROLLER_ROW_nx272), .A0 (nx657), .A1 (
          nx7291), .A2 (nx659), .B0 (CONTROLLER_nx575), .B1 (nx8471)) ;
    inv01 ix656 (.Y (nx657), .A (CONTROLLER_NxtRow_6)) ;
    inv01 ix658 (.Y (nx659), .A (CONTROLLER_ROW_nx337)) ;
    oai32 CONTROLLER_ROW_ix283 (.Y (CONTROLLER_ROW_nx282), .A0 (nx661), .A1 (
          nx7291), .A2 (nx659), .B0 (CONTROLLER_nx640), .B1 (nx8473)) ;
    inv01 ix660 (.Y (nx661), .A (CONTROLLER_NxtRow_7)) ;
    oai32 CONTROLLER_COL_ix213 (.Y (CONTROLLER_COL_nx212), .A0 (nx663), .A1 (
          nx7291), .A2 (nx665), .B0 (CONTROLLER_nx679), .B1 (nx8475)) ;
    inv01 ix662 (.Y (nx663), .A (CONTROLLER_NxtCol_0)) ;
    inv02 ix664 (.Y (nx665), .A (CONTROLLER_COL_nx335)) ;
    oai32 CONTROLLER_COL_ix223 (.Y (CONTROLLER_COL_nx222), .A0 (nx669), .A1 (
          nx7291), .A2 (nx665), .B0 (CONTROLLER_nx599), .B1 (nx8475)) ;
    inv01 ix668 (.Y (nx669), .A (CONTROLLER_NxtCol_1)) ;
    oai32 CONTROLLER_COL_ix233 (.Y (CONTROLLER_COL_nx232), .A0 (nx671), .A1 (
          nx7291), .A2 (nx665), .B0 (CONTROLLER_nx699), .B1 (nx8475)) ;
    inv01 ix670 (.Y (nx671), .A (CONTROLLER_NxtCol_2)) ;
    oai32 CONTROLLER_COL_ix243 (.Y (CONTROLLER_COL_nx242), .A0 (nx673), .A1 (
          nx7291), .A2 (nx665), .B0 (CONTROLLER_nx606), .B1 (nx8475)) ;
    inv01 ix672 (.Y (nx673), .A (CONTROLLER_NxtCol_3)) ;
    oai32 CONTROLLER_COL_ix253 (.Y (CONTROLLER_COL_nx252), .A0 (nx675), .A1 (
          nx7293), .A2 (nx665), .B0 (nx677), .B1 (nx8475)) ;
    inv01 ix674 (.Y (nx675), .A (CONTROLLER_NxtCol_4)) ;
    inv01 ix676 (.Y (nx677), .A (CONTROLLER_CurCol_4)) ;
    oai32 CONTROLLER_COL_ix263 (.Y (CONTROLLER_COL_nx262), .A0 (nx679), .A1 (
          nx7293), .A2 (nx665), .B0 (CONTROLLER_nx613), .B1 (nx8475)) ;
    inv01 ix678 (.Y (nx679), .A (CONTROLLER_NxtCol_5)) ;
    oai32 CONTROLLER_COL_ix273 (.Y (CONTROLLER_COL_nx272), .A0 (nx681), .A1 (
          nx7293), .A2 (nx683), .B0 (CONTROLLER_nx565), .B1 (nx8475)) ;
    inv01 ix680 (.Y (nx681), .A (CONTROLLER_NxtCol_6)) ;
    inv01 ix682 (.Y (nx683), .A (CONTROLLER_COL_nx337)) ;
    oai32 CONTROLLER_COL_ix283 (.Y (CONTROLLER_COL_nx282), .A0 (nx685), .A1 (
          nx7293), .A2 (nx683), .B0 (CONTROLLER_nx567), .B1 (nx8477)) ;
    inv01 ix684 (.Y (nx685), .A (CONTROLLER_NxtCol_7)) ;
    nand02 CALCULATOR_ix89 (.Y (CALCULATOR_CounterRST), .A0 (nx7337), .A1 (
           nx7305)) ;
    oai22 CALCULATOR_ix61 (.Y (MemDin[3]), .A0 (nx687), .A1 (nx689), .B0 (nx691)
          , .B1 (Instr)) ;
    inv01 ix686 (.Y (nx687), .A (CALCULATOR_L5Results_1__6)) ;
    inv01 ix688 (.Y (nx689), .A (CALCULATOR_nx22)) ;
    inv01 ix690 (.Y (nx691), .A (CALCULATOR_L5Results_1__3)) ;
    oai22 CALCULATOR_ix69 (.Y (MemDin[4]), .A0 (nx693), .A1 (nx689), .B0 (nx695)
          , .B1 (Instr)) ;
    inv01 ix692 (.Y (nx693), .A (CALCULATOR_L5Results_1__7)) ;
    inv01 ix694 (.Y (nx695), .A (CALCULATOR_L5Results_1__4)) ;
    mux21 CALCULATOR_ACCELERATOR_COUNTER_ix92 (.Y (
          CALCULATOR_ACCELERATOR_COUNTER_nx91), .A0 (nx697), .A1 (
          CALCULATOR_nx993), .S0 (AccFinishCalc)) ;
    inv01 ix696 (.Y (nx697), .A (CALCULATOR_ACCELERATOR_COUNTER_nx6)) ;
    mux21 CALCULATOR_ACCELERATOR_COUNTER_ix102 (.Y (
          CALCULATOR_ACCELERATOR_COUNTER_nx101), .A0 (nx699), .A1 (
          CALCULATOR_nx995), .S0 (AccFinishCalc)) ;
    inv01 ix698 (.Y (nx699), .A (CALCULATOR_ACCELERATOR_COUNTER_nx12)) ;
    mux21 CALCULATOR_ACCELERATOR_COUNTER_ix112 (.Y (
          CALCULATOR_ACCELERATOR_COUNTER_nx111), .A0 (nx701), .A1 (nx703), .S0 (
          AccFinishCalc)) ;
    inv01 ix700 (.Y (nx701), .A (CALCULATOR_ACCELERATOR_COUNTER_nx18)) ;
    inv01 ix702 (.Y (nx703), .A (CALCULATOR_CounterOut_3)) ;
    xnor2 CALCULATOR_ACCELERATOR_COUNTER_ix82 (.Y (
          CALCULATOR_ACCELERATOR_COUNTER_nx81), .A0 (CALCULATOR_CounterOut_0), .A1 (
          AccFinishCalc)) ;
    mux21 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix404 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx403), .A0 (nx705), .A1 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_2), .S0 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx395)) ;
    inv01 ix704 (.Y (nx705), .A (CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx391)) ;
    mux21 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix414 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx413), .A0 (nx707), .A1 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_3), .S0 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx405)) ;
    inv01 ix706 (.Y (nx707), .A (CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx403)) ;
    mux21 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix424 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx423), .A0 (nx709), .A1 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_4), .S0 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx415)) ;
    inv01 ix708 (.Y (nx709), .A (CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx413)) ;
    mux21 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix434 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx433), .A0 (nx711), .A1 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_5), .S0 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx425)) ;
    inv01 ix710 (.Y (nx711), .A (CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx423)) ;
    mux21 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix444 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx443), .A0 (nx713), .A1 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_6), .S0 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx435)) ;
    inv01 ix712 (.Y (nx713), .A (CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx433)) ;
    mux21 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix454 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx453), .A0 (nx715), .A1 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_7), .S0 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx445)) ;
    inv01 ix714 (.Y (nx715), .A (CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx443)) ;
    mux21 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix462 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx461), .A0 (nx717), .A1 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_8), .S0 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx455)) ;
    inv01 ix716 (.Y (nx717), .A (CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx453)) ;
    mux21 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix468 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx467), .A0 (nx719), .A1 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_9), .S0 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx463)) ;
    inv01 ix718 (.Y (nx719), .A (CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx461)) ;
    mux21 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix476 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx475), .A0 (nx721), .A1 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_10), .S0 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx471)) ;
    inv01 ix720 (.Y (nx721), .A (CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx467)) ;
    mux21 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix484 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx483), .A0 (nx723), .A1 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_11), .S0 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx479)) ;
    inv01 ix722 (.Y (nx723), .A (CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx475)) ;
    mux21 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix492 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx491), .A0 (nx725), .A1 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_12), .S0 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx487)) ;
    inv01 ix724 (.Y (nx725), .A (CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx483)) ;
    mux21 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix500 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx499), .A0 (nx727), .A1 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_13), .S0 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx495)) ;
    inv01 ix726 (.Y (nx727), .A (CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx491)) ;
    mux21 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix508 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx507), .A0 (nx729), .A1 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_14), .S0 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx503)) ;
    inv01 ix728 (.Y (nx729), .A (CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx499)) ;
    mux21 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix516 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx515), .A0 (nx731), .A1 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_15), .S0 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx511)) ;
    inv01 ix730 (.Y (nx731), .A (CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx507)) ;
    mux21 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix161 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_1), .A0 (nx733), .A1 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx379), .S0 (nx7317)) ;
    inv01 ix732 (.Y (nx733), .A (CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_1)) ;
    mux21 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix181 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_2), .A0 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx387), .A1 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx389), .S0 (nx7317)) ;
    mux21 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix201 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_3), .A0 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx399), .A1 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx401), .S0 (nx7317)) ;
    mux21 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix221 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_4), .A0 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx409), .A1 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx411), .S0 (nx7317)) ;
    mux21 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix241 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_5), .A0 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx419), .A1 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx421), .S0 (nx7317)) ;
    mux21 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix261 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_6), .A0 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx429), .A1 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx431), .S0 (nx7317)) ;
    mux21 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix281 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_7), .A0 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx439), .A1 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx441), .S0 (nx7317)) ;
    mux21 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix301 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_8), .A0 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx449), .A1 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx451), .S0 (nx7319)) ;
    mux21 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix321 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_9), .A0 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx469), .A1 (nx735), .S0 (nx7319)) ;
    inv01 ix734 (.Y (nx735), .A (CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx316)) ;
    mux21 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix341 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_10), .A0 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx477), .A1 (nx737), .S0 (nx7319)) ;
    inv01 ix736 (.Y (nx737), .A (CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx336)) ;
    mux21 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix361 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_11), .A0 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx485), .A1 (nx739), .S0 (nx7319)) ;
    inv01 ix738 (.Y (nx739), .A (CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx356)) ;
    mux21 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix381 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_12), .A0 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx493), .A1 (nx741), .S0 (nx7319)) ;
    inv01 ix740 (.Y (nx741), .A (CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx376)) ;
    mux21 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix401 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_13), .A0 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx501), .A1 (nx743), .S0 (nx7319)) ;
    inv01 ix742 (.Y (nx743), .A (CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx396)) ;
    mux21 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix421 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_14), .A0 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx509), .A1 (nx745), .S0 (nx7319)) ;
    inv01 ix744 (.Y (nx745), .A (CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx416)) ;
    mux21 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix441 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_15), .A0 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx517), .A1 (nx747), .S0 (nx7321)) ;
    inv01 ix746 (.Y (nx747), .A (CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx436)) ;
    mux21 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_ix461 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_16), .A0 (nx749), .A1 (
          nx751), .S0 (nx7321)) ;
    inv01 ix748 (.Y (nx749), .A (CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothP_16)) ;
    inv01 ix750 (.Y (nx751), .A (CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx456)) ;
    nor02_2x CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix81 (.Y (
             CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx80), .A0 (Instr), .A1 (
             nx7305)) ;
    nor02_2x CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix319 (.Y (
             CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642), .A0 (
             CALCULATOR_Start_dup_1144), .A1 (
             CALCULATOR_CalculatingBooth_dup_1146)) ;
    nor02_2x CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix85 (.Y (
             CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_0), .A0 (
             nx7331), .A1 (nx753)) ;
    inv01 ix752 (.Y (nx753), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_1)) ;
    mux21 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix125 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_1), .A0 (
          nx755), .A1 (nx757), .S0 (nx7331)) ;
    inv01 ix754 (.Y (nx755), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_2)) ;
    inv01 ix756 (.Y (nx757), .A (CacheWindow_0__0__0)) ;
    mux21 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix133 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_2), .A0 (
          nx759), .A1 (nx761), .S0 (nx7331)) ;
    inv01 ix758 (.Y (nx759), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_3)) ;
    inv01 ix760 (.Y (nx761), .A (CacheWindow_0__0__1)) ;
    mux21 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix141 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_3), .A0 (
          nx763), .A1 (nx765), .S0 (nx7331)) ;
    inv01 ix762 (.Y (nx763), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_4)) ;
    inv01 ix764 (.Y (nx765), .A (CacheWindow_0__0__2)) ;
    mux21 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix149 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_4), .A0 (
          nx767), .A1 (nx769), .S0 (nx7331)) ;
    inv01 ix766 (.Y (nx767), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_5)) ;
    inv01 ix768 (.Y (nx769), .A (CacheWindow_0__0__3)) ;
    mux21 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix157 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_5), .A0 (
          nx771), .A1 (nx773), .S0 (nx7331)) ;
    inv01 ix770 (.Y (nx771), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_6)) ;
    inv01 ix772 (.Y (nx773), .A (CacheWindow_0__0__4)) ;
    mux21 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix165 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_6), .A0 (
          nx775), .A1 (nx777), .S0 (nx7331)) ;
    inv01 ix774 (.Y (nx775), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_7)) ;
    inv01 ix776 (.Y (nx777), .A (CacheWindow_0__0__5)) ;
    mux21 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix173 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_7), .A0 (
          nx779), .A1 (nx781), .S0 (nx7333)) ;
    inv01 ix778 (.Y (nx779), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_8)) ;
    inv01 ix780 (.Y (nx781), .A (CacheWindow_0__0__6)) ;
    mux21 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix181 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_8), .A0 (
          nx783), .A1 (nx785), .S0 (nx7333)) ;
    inv01 ix782 (.Y (nx783), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_9)) ;
    inv01 ix784 (.Y (nx785), .A (CacheWindow_0__0__7)) ;
    nor02_2x CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix89 (.Y (
             CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_9), .A0 (
             nx7333), .A1 (nx787)) ;
    inv01 ix786 (.Y (nx787), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_10)) ;
    nor02_2x CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix93 (.Y (
             CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_10), .A0 (
             nx7333), .A1 (nx789)) ;
    inv01 ix788 (.Y (nx789), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_11)) ;
    nor02_2x CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix97 (.Y (
             CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_11), .A0 (
             nx7333), .A1 (nx791)) ;
    inv01 ix790 (.Y (nx791), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_12)) ;
    nor02_2x CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix101 (.Y (
             CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_12), .A0 (
             nx7333), .A1 (nx793)) ;
    inv01 ix792 (.Y (nx793), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_13)) ;
    nor02_2x CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix105 (.Y (
             CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_13), .A0 (
             nx7333), .A1 (nx795)) ;
    inv01 ix794 (.Y (nx795), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_14)) ;
    nor02_2x CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix109 (.Y (
             CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_14), .A0 (
             nx7335), .A1 (nx797)) ;
    inv01 ix796 (.Y (nx797), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_15)) ;
    nor02_2x CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix113 (.Y (
             CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_15), .A0 (
             nx7335), .A1 (nx799)) ;
    inv01 ix798 (.Y (nx799), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_16)) ;
    nor02_2x CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix117 (.Y (
             CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_16), .A0 (
             nx7335), .A1 (nx799)) ;
    mux21 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix189 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothOperand_0), .A0 (nx801), .A1 (
          nx803), .S0 (nx7323)) ;
    inv01 ix800 (.Y (nx801), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_0)) ;
    inv01 ix802 (.Y (nx803), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_0)) ;
    mux21 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix197 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothOperand_1), .A0 (nx805), .A1 (
          nx807), .S0 (nx7323)) ;
    inv01 ix804 (.Y (nx805), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_1)) ;
    inv01 ix806 (.Y (nx807), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_1)) ;
    mux21 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix205 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothOperand_2), .A0 (nx809), .A1 (
          nx811), .S0 (nx7323)) ;
    inv01 ix808 (.Y (nx809), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_2)) ;
    inv01 ix810 (.Y (nx811), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_2)) ;
    mux21 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix213 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothOperand_3), .A0 (nx813), .A1 (
          nx815), .S0 (nx7323)) ;
    inv01 ix812 (.Y (nx813), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_3)) ;
    inv01 ix814 (.Y (nx815), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_3)) ;
    mux21 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix221 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothOperand_4), .A0 (nx817), .A1 (
          nx819), .S0 (nx7323)) ;
    inv01 ix816 (.Y (nx817), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_4)) ;
    inv01 ix818 (.Y (nx819), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_4)) ;
    mux21 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix229 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothOperand_5), .A0 (nx821), .A1 (
          nx823), .S0 (nx7325)) ;
    inv01 ix820 (.Y (nx821), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_5)) ;
    inv01 ix822 (.Y (nx823), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_5)) ;
    mux21 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix237 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothOperand_6), .A0 (nx825), .A1 (
          nx827), .S0 (nx7325)) ;
    inv01 ix824 (.Y (nx825), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_6)) ;
    inv01 ix826 (.Y (nx827), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_6)) ;
    mux21 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix245 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothOperand_7), .A0 (nx829), .A1 (
          nx831), .S0 (nx7325)) ;
    inv01 ix828 (.Y (nx829), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_7)) ;
    inv01 ix830 (.Y (nx831), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_7)) ;
    mux21 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix253 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothOperand_8), .A0 (nx833), .A1 (
          nx835), .S0 (nx7325)) ;
    inv01 ix832 (.Y (nx833), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_8)) ;
    inv01 ix834 (.Y (nx835), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_8)) ;
    mux21 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix261 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothOperand_9), .A0 (nx837), .A1 (
          nx839), .S0 (nx7325)) ;
    inv01 ix836 (.Y (nx837), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_9)) ;
    inv01 ix838 (.Y (nx839), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_9)) ;
    mux21 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix269 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothOperand_10), .A0 (nx841), .A1 (
          nx843), .S0 (nx7325)) ;
    inv01 ix840 (.Y (nx841), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_10)) ;
    inv01 ix842 (.Y (nx843), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_10)) ;
    mux21 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix277 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothOperand_11), .A0 (nx845), .A1 (
          nx847), .S0 (nx7325)) ;
    inv01 ix844 (.Y (nx845), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_11)) ;
    inv01 ix846 (.Y (nx847), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_11)) ;
    mux21 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix285 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothOperand_12), .A0 (nx849), .A1 (
          nx851), .S0 (nx7327)) ;
    inv01 ix848 (.Y (nx849), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_12)) ;
    inv01 ix850 (.Y (nx851), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_12)) ;
    mux21 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix293 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothOperand_13), .A0 (nx853), .A1 (
          nx855), .S0 (nx7327)) ;
    inv01 ix852 (.Y (nx853), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_13)) ;
    inv01 ix854 (.Y (nx855), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_13)) ;
    mux21 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix301 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothOperand_14), .A0 (nx857), .A1 (
          nx859), .S0 (nx7327)) ;
    inv01 ix856 (.Y (nx857), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_14)) ;
    inv01 ix858 (.Y (nx859), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_14)) ;
    mux21 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix309 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothOperand_15), .A0 (nx861), .A1 (
          nx863), .S0 (nx7327)) ;
    inv01 ix860 (.Y (nx861), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_15)) ;
    inv01 ix862 (.Y (nx863), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_15)) ;
    mux21 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix317 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BoothOperand_16), .A0 (nx865), .A1 (
          nx867), .S0 (nx7327)) ;
    inv01 ix864 (.Y (nx865), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_16)) ;
    inv01 ix866 (.Y (nx867), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_16)) ;
    xnor2 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix321 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_AddPToBoothOperand), .A0 (nx7327), .A1 (
          nx733)) ;
    oai32 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix393 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .A0 (
          nx8479), .A1 (RST), .A2 (nx7379), .B0 (nx803), .B1 (nx871)) ;
    oai32 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix403 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .A0 (
          nx8479), .A1 (RST), .A2 (nx7379), .B0 (nx807), .B1 (nx871)) ;
    oai32 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix413 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .A0 (
          nx8479), .A1 (RST), .A2 (nx7379), .B0 (nx811), .B1 (nx871)) ;
    oai32 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix423 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .A0 (
          nx8479), .A1 (RST), .A2 (nx7379), .B0 (nx815), .B1 (nx871)) ;
    oai32 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix433 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .A0 (
          nx8479), .A1 (RST), .A2 (nx7379), .B0 (nx819), .B1 (nx871)) ;
    oai32 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix443 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .A0 (
          nx8479), .A1 (RST), .A2 (nx7379), .B0 (nx823), .B1 (nx871)) ;
    oai32 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix453 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .A0 (
          nx8479), .A1 (RST), .A2 (nx7381), .B0 (nx827), .B1 (nx871)) ;
    oai32 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix463 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .A0 (
          nx8481), .A1 (RST), .A2 (nx7381), .B0 (nx831), .B1 (nx873)) ;
    oai32 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix473 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .A0 (
          nx8481), .A1 (RST), .A2 (nx7381), .B0 (nx835), .B1 (nx873)) ;
    oai32 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix483 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .A0 (
          nx875), .A1 (RST), .A2 (nx7381), .B0 (nx839), .B1 (nx873)) ;
    inv01 ix874 (.Y (nx875), .A (CacheFilter_0__0__0)) ;
    oai32 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix493 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .A0 (
          nx877), .A1 (RST), .A2 (nx7381), .B0 (nx843), .B1 (nx873)) ;
    inv01 ix876 (.Y (nx877), .A (CacheFilter_0__0__1)) ;
    oai32 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix503 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .A0 (
          nx879), .A1 (RST), .A2 (nx7381), .B0 (nx847), .B1 (nx873)) ;
    inv01 ix878 (.Y (nx879), .A (CacheFilter_0__0__2)) ;
    oai32 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix513 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .A0 (
          nx881), .A1 (RST), .A2 (nx7381), .B0 (nx851), .B1 (nx873)) ;
    inv01 ix880 (.Y (nx881), .A (CacheFilter_0__0__3)) ;
    oai32 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix523 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .A0 (
          nx883), .A1 (RST), .A2 (nx7383), .B0 (nx855), .B1 (nx873)) ;
    inv01 ix882 (.Y (nx883), .A (CacheFilter_0__0__4)) ;
    oai32 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix533 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .A0 (
          nx885), .A1 (RST), .A2 (nx7383), .B0 (nx859), .B1 (nx887)) ;
    inv01 ix884 (.Y (nx885), .A (CacheFilter_0__0__5)) ;
    inv01 ix886 (.Y (nx887), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566)) ;
    oai32 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix543 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .A0 (
          nx889), .A1 (RST), .A2 (nx7383), .B0 (nx863), .B1 (nx887)) ;
    inv01 ix888 (.Y (nx889), .A (CacheFilter_0__0__6)) ;
    oai32 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix553 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .A0 (
          nx891), .A1 (RST), .A2 (nx7383), .B0 (nx867), .B1 (nx887)) ;
    inv01 ix890 (.Y (nx891), .A (CacheFilter_0__0__7)) ;
    nand02_2x CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix633 (.Y (
              nx871), .A0 (nx7337), .A1 (nx7383)) ;
    nand02_2x CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix635 (.Y (
              nx873), .A0 (nx7337), .A1 (nx7383)) ;
    oai32 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix393 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .A0 (
          nx8481), .A1 (RST), .A2 (nx7385), .B0 (nx801), .B1 (nx893)) ;
    oai32 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix403 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .A0 (
          nx8481), .A1 (RST), .A2 (nx7385), .B0 (nx805), .B1 (nx893)) ;
    oai32 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix413 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .A0 (
          nx8481), .A1 (RST), .A2 (nx7385), .B0 (nx809), .B1 (nx893)) ;
    oai32 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix423 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .A0 (
          nx8481), .A1 (RST), .A2 (nx7385), .B0 (nx813), .B1 (nx893)) ;
    oai32 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix433 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .A0 (
          nx8481), .A1 (RST), .A2 (nx7385), .B0 (nx817), .B1 (nx893)) ;
    oai32 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix443 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .A0 (
          nx8483), .A1 (RST), .A2 (nx7385), .B0 (nx821), .B1 (nx893)) ;
    oai32 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix453 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .A0 (
          nx8483), .A1 (RST), .A2 (nx7387), .B0 (nx825), .B1 (nx893)) ;
    oai32 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix463 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .A0 (
          nx8483), .A1 (RST), .A2 (nx7387), .B0 (nx829), .B1 (nx895)) ;
    oai32 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix473 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .A0 (
          nx8483), .A1 (RST), .A2 (nx7387), .B0 (nx833), .B1 (nx895)) ;
    oai32 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix483 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .A0 (
          nx875), .A1 (RST), .A2 (nx7387), .B0 (nx837), .B1 (nx895)) ;
    oai32 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix493 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .A0 (
          nx897), .A1 (RST), .A2 (nx7387), .B0 (nx841), .B1 (nx895)) ;
    inv01 ix896 (.Y (nx897), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_10)) ;
    oai32 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix503 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .A0 (
          nx899), .A1 (RST), .A2 (nx7387), .B0 (nx845), .B1 (nx895)) ;
    inv01 ix898 (.Y (nx899), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_11)) ;
    oai32 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix513 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .A0 (
          nx901), .A1 (RST), .A2 (nx7387), .B0 (nx849), .B1 (nx895)) ;
    inv01 ix900 (.Y (nx901), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_12)) ;
    oai32 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix523 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .A0 (
          nx903), .A1 (RST), .A2 (nx7389), .B0 (nx853), .B1 (nx895)) ;
    inv01 ix902 (.Y (nx903), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_13)) ;
    oai32 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix533 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .A0 (
          nx905), .A1 (RST), .A2 (nx7389), .B0 (nx857), .B1 (nx907)) ;
    inv01 ix904 (.Y (nx905), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_14)) ;
    inv01 ix906 (.Y (nx907), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566)) ;
    oai32 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix543 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .A0 (
          nx909), .A1 (RST), .A2 (nx7389), .B0 (nx861), .B1 (nx907)) ;
    inv01 ix908 (.Y (nx909), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_15)) ;
    oai32 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix553 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .A0 (
          nx911), .A1 (RST), .A2 (nx7389), .B0 (nx865), .B1 (nx907)) ;
    inv01 ix910 (.Y (nx911), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_16)) ;
    nand02_2x CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix633 (.Y (
              nx893), .A0 (nx7337), .A1 (nx7389)) ;
    nand02_2x CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix635 (.Y (
              nx895), .A0 (nx7337), .A1 (nx7389)) ;
    oai32 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix393 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .A0 (
          nx913), .A1 (RST), .A2 (nx7391), .B0 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx384), .B1 (nx915)) ;
    inv01 ix912 (.Y (nx913), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_0)) ;
    oai32 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix403 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .A0 (
          nx917), .A1 (RST), .A2 (nx7391), .B0 (nx733), .B1 (nx915)) ;
    inv01 ix916 (.Y (nx917), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_1)) ;
    oai32 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix413 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .A0 (
          nx919), .A1 (RST), .A2 (nx7391), .B0 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx387), .B1 (nx915)) ;
    inv01 ix918 (.Y (nx919), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_2)) ;
    oai32 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix423 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .A0 (
          nx921), .A1 (RST), .A2 (nx7391), .B0 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx399), .B1 (nx915)) ;
    inv01 ix920 (.Y (nx921), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_3)) ;
    oai32 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix433 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .A0 (
          nx923), .A1 (RST), .A2 (nx7391), .B0 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx409), .B1 (nx915)) ;
    inv01 ix922 (.Y (nx923), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_4)) ;
    oai32 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix443 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .A0 (
          nx925), .A1 (RST), .A2 (nx7391), .B0 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx419), .B1 (nx915)) ;
    inv01 ix924 (.Y (nx925), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_5)) ;
    oai32 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix453 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .A0 (
          nx927), .A1 (RST), .A2 (nx7391), .B0 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx429), .B1 (nx915)) ;
    inv01 ix926 (.Y (nx927), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_6)) ;
    oai32 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix463 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .A0 (
          nx929), .A1 (RST), .A2 (nx7393), .B0 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx439), .B1 (nx931)) ;
    inv01 ix928 (.Y (nx929), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_7)) ;
    oai32 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix473 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .A0 (
          nx933), .A1 (RST), .A2 (nx7393), .B0 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx449), .B1 (nx931)) ;
    inv01 ix932 (.Y (nx933), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_8)) ;
    oai32 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix483 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .A0 (
          nx935), .A1 (RST), .A2 (nx7393), .B0 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx469), .B1 (nx931)) ;
    inv01 ix934 (.Y (nx935), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_9)) ;
    oai32 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix493 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .A0 (
          nx937), .A1 (RST), .A2 (nx7393), .B0 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx477), .B1 (nx931)) ;
    inv01 ix936 (.Y (nx937), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_10)) ;
    oai32 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix503 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .A0 (
          nx939), .A1 (RST), .A2 (nx7393), .B0 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx485), .B1 (nx931)) ;
    inv01 ix938 (.Y (nx939), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_11)) ;
    oai32 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix513 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .A0 (
          nx941), .A1 (RST), .A2 (nx7393), .B0 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx493), .B1 (nx931)) ;
    inv01 ix940 (.Y (nx941), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_12)) ;
    oai32 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix523 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .A0 (
          nx943), .A1 (RST), .A2 (nx7393), .B0 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx501), .B1 (nx931)) ;
    inv01 ix942 (.Y (nx943), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_13)) ;
    oai32 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix533 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .A0 (
          nx945), .A1 (RST), .A2 (nx7395), .B0 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx509), .B1 (nx947)) ;
    inv01 ix944 (.Y (nx945), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_14)) ;
    inv01 ix946 (.Y (nx947), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566)) ;
    oai32 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix543 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .A0 (
          nx949), .A1 (RST), .A2 (nx7395), .B0 (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_nx517), .B1 (nx947)) ;
    inv01 ix948 (.Y (nx949), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_15)) ;
    oai32 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix553 (.Y (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .A0 (
          nx951), .A1 (RST), .A2 (nx7395), .B0 (nx749), .B1 (nx947)) ;
    inv01 ix950 (.Y (nx951), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_16)) ;
    nand02_2x CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix633 (.Y (
              nx915), .A0 (nx7337), .A1 (nx7395)) ;
    nand02_2x CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix635 (.Y (
              nx931), .A0 (nx7337), .A1 (nx7395)) ;
    mux21 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix404 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx403), .A0 (nx953), .A1 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_2), .S0 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx395)) ;
    inv01 ix952 (.Y (nx953), .A (CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx391)) ;
    mux21 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix414 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx413), .A0 (nx955), .A1 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_3), .S0 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx405)) ;
    inv01 ix954 (.Y (nx955), .A (CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx403)) ;
    mux21 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix424 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx423), .A0 (nx957), .A1 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_4), .S0 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx415)) ;
    inv01 ix956 (.Y (nx957), .A (CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx413)) ;
    mux21 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix434 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx433), .A0 (nx959), .A1 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_5), .S0 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx425)) ;
    inv01 ix958 (.Y (nx959), .A (CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx423)) ;
    mux21 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix444 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx443), .A0 (nx961), .A1 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_6), .S0 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx435)) ;
    inv01 ix960 (.Y (nx961), .A (CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx433)) ;
    mux21 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix454 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx453), .A0 (nx963), .A1 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_7), .S0 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx445)) ;
    inv01 ix962 (.Y (nx963), .A (CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx443)) ;
    mux21 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix462 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx461), .A0 (nx965), .A1 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_8), .S0 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx455)) ;
    inv01 ix964 (.Y (nx965), .A (CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx453)) ;
    mux21 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix468 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx467), .A0 (nx967), .A1 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_9), .S0 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx463)) ;
    inv01 ix966 (.Y (nx967), .A (CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx461)) ;
    mux21 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix476 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx475), .A0 (nx969), .A1 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_10), .S0 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx471)) ;
    inv01 ix968 (.Y (nx969), .A (CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx467)) ;
    mux21 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix484 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx483), .A0 (nx971), .A1 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_11), .S0 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx479)) ;
    inv01 ix970 (.Y (nx971), .A (CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx475)) ;
    mux21 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix492 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx491), .A0 (nx973), .A1 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_12), .S0 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx487)) ;
    inv01 ix972 (.Y (nx973), .A (CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx483)) ;
    mux21 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix500 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx499), .A0 (nx975), .A1 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_13), .S0 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx495)) ;
    inv01 ix974 (.Y (nx975), .A (CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx491)) ;
    mux21 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix508 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx507), .A0 (nx977), .A1 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_14), .S0 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx503)) ;
    inv01 ix976 (.Y (nx977), .A (CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx499)) ;
    mux21 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix516 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx515), .A0 (nx979), .A1 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_15), .S0 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx511)) ;
    inv01 ix978 (.Y (nx979), .A (CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx507)) ;
    mux21 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix161 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_1), .A0 (nx981), .A1 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx379), .S0 (nx7399)) ;
    inv01 ix980 (.Y (nx981), .A (CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_1)) ;
    mux21 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix181 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_2), .A0 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx387), .A1 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx389), .S0 (nx7399)) ;
    mux21 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix201 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_3), .A0 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx399), .A1 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx401), .S0 (nx7399)) ;
    mux21 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix221 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_4), .A0 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx409), .A1 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx411), .S0 (nx7399)) ;
    mux21 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix241 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_5), .A0 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx419), .A1 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx421), .S0 (nx7399)) ;
    mux21 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix261 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_6), .A0 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx429), .A1 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx431), .S0 (nx7399)) ;
    mux21 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix281 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_7), .A0 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx439), .A1 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx441), .S0 (nx7399)) ;
    mux21 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix301 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_8), .A0 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx449), .A1 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx451), .S0 (nx7401)) ;
    mux21 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix321 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_9), .A0 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx469), .A1 (nx983), .S0 (nx7401)) ;
    inv01 ix982 (.Y (nx983), .A (CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx316)) ;
    mux21 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix341 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_10), .A0 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx477), .A1 (nx985), .S0 (nx7401)) ;
    inv01 ix984 (.Y (nx985), .A (CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx336)) ;
    mux21 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix361 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_11), .A0 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx485), .A1 (nx987), .S0 (nx7401)) ;
    inv01 ix986 (.Y (nx987), .A (CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx356)) ;
    mux21 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix381 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_12), .A0 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx493), .A1 (nx989), .S0 (nx7401)) ;
    inv01 ix988 (.Y (nx989), .A (CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx376)) ;
    mux21 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix401 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_13), .A0 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx501), .A1 (nx991), .S0 (nx7401)) ;
    inv01 ix990 (.Y (nx991), .A (CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx396)) ;
    mux21 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix421 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_14), .A0 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx509), .A1 (nx993), .S0 (nx7401)) ;
    inv01 ix992 (.Y (nx993), .A (CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx416)) ;
    mux21 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix441 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_15), .A0 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx517), .A1 (nx995), .S0 (nx7403)) ;
    inv01 ix994 (.Y (nx995), .A (CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx436)) ;
    mux21 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_ix461 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_16), .A0 (nx997), .A1 (
          nx999), .S0 (nx7403)) ;
    inv01 ix996 (.Y (nx997), .A (CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothP_16)) ;
    inv01 ix998 (.Y (nx999), .A (CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx456)) ;
    nor02_2x CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix81 (.Y (
             CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx80), .A0 (Instr), .A1 (
             nx7305)) ;
    nor02_2x CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix319 (.Y (
             CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642), .A0 (
             CALCULATOR_Start_dup_1149), .A1 (
             CALCULATOR_CalculatingBooth_dup_1146)) ;
    nor02_2x CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix85 (.Y (
             CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_0), .A0 (
             nx7413), .A1 (nx1001)) ;
    inv01 ix1000 (.Y (nx1001), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_1)) ;
    mux21 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix125 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_1), .A0 (
          nx1003), .A1 (nx1005), .S0 (nx7413)) ;
    inv01 ix1002 (.Y (nx1003), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_2)) ;
    inv01 ix1004 (.Y (nx1005), .A (CacheWindow_0__1__0)) ;
    mux21 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix133 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_2), .A0 (
          nx1007), .A1 (nx1009), .S0 (nx7413)) ;
    inv01 ix1006 (.Y (nx1007), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_3)) ;
    inv01 ix1008 (.Y (nx1009), .A (CacheWindow_0__1__1)) ;
    mux21 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix141 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_3), .A0 (
          nx1011), .A1 (nx1013), .S0 (nx7413)) ;
    inv01 ix1010 (.Y (nx1011), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_4)) ;
    inv01 ix1012 (.Y (nx1013), .A (CacheWindow_0__1__2)) ;
    mux21 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix149 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_4), .A0 (
          nx1015), .A1 (nx1017), .S0 (nx7413)) ;
    inv01 ix1014 (.Y (nx1015), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_5)) ;
    inv01 ix1016 (.Y (nx1017), .A (CacheWindow_0__1__3)) ;
    mux21 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix157 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_5), .A0 (
          nx1019), .A1 (nx1021), .S0 (nx7413)) ;
    inv01 ix1018 (.Y (nx1019), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_6)) ;
    inv01 ix1020 (.Y (nx1021), .A (CacheWindow_0__1__4)) ;
    mux21 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix165 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_6), .A0 (
          nx1023), .A1 (nx1025), .S0 (nx7413)) ;
    inv01 ix1022 (.Y (nx1023), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_7)) ;
    inv01 ix1024 (.Y (nx1025), .A (CacheWindow_0__1__5)) ;
    mux21 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix173 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_7), .A0 (
          nx1027), .A1 (nx1029), .S0 (nx7415)) ;
    inv01 ix1026 (.Y (nx1027), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_8)) ;
    inv01 ix1028 (.Y (nx1029), .A (CacheWindow_0__1__6)) ;
    mux21 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix181 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_8), .A0 (
          nx1031), .A1 (nx1033), .S0 (nx7415)) ;
    inv01 ix1030 (.Y (nx1031), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_9)) ;
    inv01 ix1032 (.Y (nx1033), .A (CacheWindow_0__1__7)) ;
    nor02_2x CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix89 (.Y (
             CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_9), .A0 (
             nx7415), .A1 (nx1035)) ;
    inv01 ix1034 (.Y (nx1035), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_10)) ;
    nor02_2x CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix93 (.Y (
             CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_10), .A0 (
             nx7415), .A1 (nx1037)) ;
    inv01 ix1036 (.Y (nx1037), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_11)) ;
    nor02_2x CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix97 (.Y (
             CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_11), .A0 (
             nx7415), .A1 (nx1039)) ;
    inv01 ix1038 (.Y (nx1039), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_12)) ;
    nor02_2x CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix101 (.Y (
             CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_12), .A0 (
             nx7415), .A1 (nx1041)) ;
    inv01 ix1040 (.Y (nx1041), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_13)) ;
    nor02_2x CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix105 (.Y (
             CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_13), .A0 (
             nx7415), .A1 (nx1043)) ;
    inv01 ix1042 (.Y (nx1043), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_14)) ;
    nor02_2x CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix109 (.Y (
             CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_14), .A0 (
             nx7417), .A1 (nx1045)) ;
    inv01 ix1044 (.Y (nx1045), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_15)) ;
    nor02_2x CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix113 (.Y (
             CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_15), .A0 (
             nx7417), .A1 (nx1047)) ;
    inv01 ix1046 (.Y (nx1047), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_16)) ;
    nor02_2x CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix117 (.Y (
             CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_16), .A0 (
             nx7417), .A1 (nx1047)) ;
    mux21 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix189 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothOperand_0), .A0 (nx1049), .A1 (
          nx1051), .S0 (nx7405)) ;
    inv01 ix1048 (.Y (nx1049), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_0)) ;
    inv01 ix1050 (.Y (nx1051), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_0)) ;
    mux21 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix197 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothOperand_1), .A0 (nx1053), .A1 (
          nx1055), .S0 (nx7405)) ;
    inv01 ix1052 (.Y (nx1053), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_1)) ;
    inv01 ix1054 (.Y (nx1055), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_1)) ;
    mux21 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix205 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothOperand_2), .A0 (nx1057), .A1 (
          nx1059), .S0 (nx7405)) ;
    inv01 ix1056 (.Y (nx1057), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_2)) ;
    inv01 ix1058 (.Y (nx1059), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_2)) ;
    mux21 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix213 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothOperand_3), .A0 (nx1061), .A1 (
          nx1063), .S0 (nx7405)) ;
    inv01 ix1060 (.Y (nx1061), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_3)) ;
    inv01 ix1062 (.Y (nx1063), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_3)) ;
    mux21 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix221 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothOperand_4), .A0 (nx1065), .A1 (
          nx1067), .S0 (nx7405)) ;
    inv01 ix1064 (.Y (nx1065), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_4)) ;
    inv01 ix1066 (.Y (nx1067), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_4)) ;
    mux21 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix229 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothOperand_5), .A0 (nx1069), .A1 (
          nx1071), .S0 (nx7407)) ;
    inv01 ix1068 (.Y (nx1069), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_5)) ;
    inv01 ix1070 (.Y (nx1071), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_5)) ;
    mux21 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix237 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothOperand_6), .A0 (nx1073), .A1 (
          nx1075), .S0 (nx7407)) ;
    inv01 ix1072 (.Y (nx1073), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_6)) ;
    inv01 ix1074 (.Y (nx1075), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_6)) ;
    mux21 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix245 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothOperand_7), .A0 (nx1077), .A1 (
          nx1079), .S0 (nx7407)) ;
    inv01 ix1076 (.Y (nx1077), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_7)) ;
    inv01 ix1078 (.Y (nx1079), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_7)) ;
    mux21 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix253 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothOperand_8), .A0 (nx1081), .A1 (
          nx1083), .S0 (nx7407)) ;
    inv01 ix1080 (.Y (nx1081), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_8)) ;
    inv01 ix1082 (.Y (nx1083), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_8)) ;
    mux21 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix261 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothOperand_9), .A0 (nx1085), .A1 (
          nx1087), .S0 (nx7407)) ;
    inv01 ix1084 (.Y (nx1085), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_9)) ;
    inv01 ix1086 (.Y (nx1087), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_9)) ;
    mux21 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix269 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothOperand_10), .A0 (nx1089), .A1 (
          nx1091), .S0 (nx7407)) ;
    inv01 ix1088 (.Y (nx1089), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_10)) ;
    inv01 ix1090 (.Y (nx1091), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_10)) ;
    mux21 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix277 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothOperand_11), .A0 (nx1093), .A1 (
          nx1095), .S0 (nx7407)) ;
    inv01 ix1092 (.Y (nx1093), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_11)) ;
    inv01 ix1094 (.Y (nx1095), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_11)) ;
    mux21 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix285 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothOperand_12), .A0 (nx1097), .A1 (
          nx1099), .S0 (nx7409)) ;
    inv01 ix1096 (.Y (nx1097), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_12)) ;
    inv01 ix1098 (.Y (nx1099), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_12)) ;
    mux21 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix293 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothOperand_13), .A0 (nx1101), .A1 (
          nx1103), .S0 (nx7409)) ;
    inv01 ix1100 (.Y (nx1101), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_13)) ;
    inv01 ix1102 (.Y (nx1103), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_13)) ;
    mux21 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix301 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothOperand_14), .A0 (nx1105), .A1 (
          nx1107), .S0 (nx7409)) ;
    inv01 ix1104 (.Y (nx1105), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_14)) ;
    inv01 ix1106 (.Y (nx1107), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_14)) ;
    mux21 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix309 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothOperand_15), .A0 (nx1109), .A1 (
          nx1111), .S0 (nx7409)) ;
    inv01 ix1108 (.Y (nx1109), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_15)) ;
    inv01 ix1110 (.Y (nx1111), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_15)) ;
    mux21 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix317 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BoothOperand_16), .A0 (nx1113), .A1 (
          nx1115), .S0 (nx7409)) ;
    inv01 ix1112 (.Y (nx1113), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_16)) ;
    inv01 ix1114 (.Y (nx1115), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_16)) ;
    xnor2 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix321 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_AddPToBoothOperand), .A0 (nx7409), .A1 (
          nx981)) ;
    oai32 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix393 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .A0 (
          nx8485), .A1 (RST), .A2 (nx7419), .B0 (nx1051), .B1 (nx1119)) ;
    oai32 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix403 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .A0 (
          nx8485), .A1 (RST), .A2 (nx7419), .B0 (nx1055), .B1 (nx1119)) ;
    oai32 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix413 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .A0 (
          nx8485), .A1 (RST), .A2 (nx7419), .B0 (nx1059), .B1 (nx1119)) ;
    oai32 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix423 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .A0 (
          nx8485), .A1 (RST), .A2 (nx7419), .B0 (nx1063), .B1 (nx1119)) ;
    oai32 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix433 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .A0 (
          nx8485), .A1 (RST), .A2 (nx7419), .B0 (nx1067), .B1 (nx1119)) ;
    oai32 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix443 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .A0 (
          nx8485), .A1 (RST), .A2 (nx7419), .B0 (nx1071), .B1 (nx1119)) ;
    oai32 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix453 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .A0 (
          nx8485), .A1 (RST), .A2 (nx7421), .B0 (nx1075), .B1 (nx1119)) ;
    oai32 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix463 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .A0 (
          nx8487), .A1 (RST), .A2 (nx7421), .B0 (nx1079), .B1 (nx1121)) ;
    oai32 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix473 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .A0 (
          nx8487), .A1 (RST), .A2 (nx7421), .B0 (nx1083), .B1 (nx1121)) ;
    oai32 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix483 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .A0 (
          nx1123), .A1 (RST), .A2 (nx7421), .B0 (nx1087), .B1 (nx1121)) ;
    inv01 ix1122 (.Y (nx1123), .A (CacheFilter_0__1__0)) ;
    oai32 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix493 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .A0 (
          nx1125), .A1 (RST), .A2 (nx7421), .B0 (nx1091), .B1 (nx1121)) ;
    inv01 ix1124 (.Y (nx1125), .A (CacheFilter_0__1__1)) ;
    oai32 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix503 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .A0 (
          nx1127), .A1 (RST), .A2 (nx7421), .B0 (nx1095), .B1 (nx1121)) ;
    inv01 ix1126 (.Y (nx1127), .A (CacheFilter_0__1__2)) ;
    oai32 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix513 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .A0 (
          nx1129), .A1 (RST), .A2 (nx7421), .B0 (nx1099), .B1 (nx1121)) ;
    inv01 ix1128 (.Y (nx1129), .A (CacheFilter_0__1__3)) ;
    oai32 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix523 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .A0 (
          nx1131), .A1 (RST), .A2 (nx7423), .B0 (nx1103), .B1 (nx1121)) ;
    inv01 ix1130 (.Y (nx1131), .A (CacheFilter_0__1__4)) ;
    oai32 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix533 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .A0 (
          nx1133), .A1 (RST), .A2 (nx7423), .B0 (nx1107), .B1 (nx1135)) ;
    inv01 ix1132 (.Y (nx1133), .A (CacheFilter_0__1__5)) ;
    inv01 ix1134 (.Y (nx1135), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566)) ;
    oai32 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix543 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .A0 (
          nx1137), .A1 (RST), .A2 (nx7423), .B0 (nx1111), .B1 (nx1135)) ;
    inv01 ix1136 (.Y (nx1137), .A (CacheFilter_0__1__6)) ;
    oai32 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix553 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .A0 (
          nx1139), .A1 (RST), .A2 (nx7423), .B0 (nx1115), .B1 (nx1135)) ;
    inv01 ix1138 (.Y (nx1139), .A (CacheFilter_0__1__7)) ;
    nand02_2x CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix633 (.Y (
              nx1119), .A0 (nx7339), .A1 (nx7423)) ;
    nand02_2x CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix635 (.Y (
              nx1121), .A0 (nx7339), .A1 (nx7423)) ;
    oai32 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix393 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .A0 (
          nx8487), .A1 (RST), .A2 (nx7425), .B0 (nx1049), .B1 (nx1141)) ;
    oai32 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix403 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .A0 (
          nx8487), .A1 (RST), .A2 (nx7425), .B0 (nx1053), .B1 (nx1141)) ;
    oai32 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix413 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .A0 (
          nx8487), .A1 (RST), .A2 (nx7425), .B0 (nx1057), .B1 (nx1141)) ;
    oai32 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix423 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .A0 (
          nx8487), .A1 (RST), .A2 (nx7425), .B0 (nx1061), .B1 (nx1141)) ;
    oai32 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix433 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .A0 (
          nx8487), .A1 (RST), .A2 (nx7425), .B0 (nx1065), .B1 (nx1141)) ;
    oai32 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix443 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .A0 (
          nx8489), .A1 (RST), .A2 (nx7425), .B0 (nx1069), .B1 (nx1141)) ;
    oai32 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix453 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .A0 (
          nx8489), .A1 (RST), .A2 (nx7427), .B0 (nx1073), .B1 (nx1141)) ;
    oai32 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix463 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .A0 (
          nx8489), .A1 (RST), .A2 (nx7427), .B0 (nx1077), .B1 (nx1143)) ;
    oai32 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix473 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .A0 (
          nx8489), .A1 (RST), .A2 (nx7427), .B0 (nx1081), .B1 (nx1143)) ;
    oai32 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix483 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .A0 (
          nx1123), .A1 (RST), .A2 (nx7427), .B0 (nx1085), .B1 (nx1143)) ;
    oai32 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix493 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .A0 (
          nx1145), .A1 (RST), .A2 (nx7427), .B0 (nx1089), .B1 (nx1143)) ;
    inv01 ix1144 (.Y (nx1145), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_10)) ;
    oai32 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix503 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .A0 (
          nx1147), .A1 (RST), .A2 (nx7427), .B0 (nx1093), .B1 (nx1143)) ;
    inv01 ix1146 (.Y (nx1147), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_11)) ;
    oai32 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix513 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .A0 (
          nx1149), .A1 (RST), .A2 (nx7427), .B0 (nx1097), .B1 (nx1143)) ;
    inv01 ix1148 (.Y (nx1149), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_12)) ;
    oai32 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix523 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .A0 (
          nx1151), .A1 (RST), .A2 (nx7429), .B0 (nx1101), .B1 (nx1143)) ;
    inv01 ix1150 (.Y (nx1151), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_13)) ;
    oai32 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix533 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .A0 (
          nx1153), .A1 (RST), .A2 (nx7429), .B0 (nx1105), .B1 (nx1155)) ;
    inv01 ix1152 (.Y (nx1153), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_14)) ;
    inv01 ix1154 (.Y (nx1155), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566)) ;
    oai32 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix543 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .A0 (
          nx1157), .A1 (RST), .A2 (nx7429), .B0 (nx1109), .B1 (nx1155)) ;
    inv01 ix1156 (.Y (nx1157), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_15)) ;
    oai32 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix553 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .A0 (
          nx1159), .A1 (RST), .A2 (nx7429), .B0 (nx1113), .B1 (nx1155)) ;
    inv01 ix1158 (.Y (nx1159), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_16)) ;
    nand02_2x CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix633 (.Y (
              nx1141), .A0 (nx7339), .A1 (nx7429)) ;
    nand02_2x CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix635 (.Y (
              nx1143), .A0 (nx7339), .A1 (nx7429)) ;
    oai32 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix393 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .A0 (
          nx1161), .A1 (RST), .A2 (nx7431), .B0 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx384), .B1 (nx1163)) ;
    inv01 ix1160 (.Y (nx1161), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_0)) ;
    oai32 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix403 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .A0 (
          nx1165), .A1 (RST), .A2 (nx7431), .B0 (nx981), .B1 (nx1163)) ;
    inv01 ix1164 (.Y (nx1165), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_1)) ;
    oai32 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix413 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .A0 (
          nx1167), .A1 (RST), .A2 (nx7431), .B0 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx387), .B1 (nx1163)) ;
    inv01 ix1166 (.Y (nx1167), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_2)) ;
    oai32 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix423 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .A0 (
          nx1169), .A1 (RST), .A2 (nx7431), .B0 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx399), .B1 (nx1163)) ;
    inv01 ix1168 (.Y (nx1169), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_3)) ;
    oai32 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix433 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .A0 (
          nx1171), .A1 (RST), .A2 (nx7431), .B0 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx409), .B1 (nx1163)) ;
    inv01 ix1170 (.Y (nx1171), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_4)) ;
    oai32 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix443 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .A0 (
          nx1173), .A1 (RST), .A2 (nx7431), .B0 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx419), .B1 (nx1163)) ;
    inv01 ix1172 (.Y (nx1173), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_5)) ;
    oai32 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix453 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .A0 (
          nx1175), .A1 (RST), .A2 (nx7431), .B0 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx429), .B1 (nx1163)) ;
    inv01 ix1174 (.Y (nx1175), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_6)) ;
    oai32 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix463 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .A0 (
          nx1177), .A1 (RST), .A2 (nx7433), .B0 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx439), .B1 (nx1179)) ;
    inv01 ix1176 (.Y (nx1177), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_7)) ;
    oai32 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix473 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .A0 (
          nx1181), .A1 (RST), .A2 (nx7433), .B0 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx449), .B1 (nx1179)) ;
    inv01 ix1180 (.Y (nx1181), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_8)) ;
    oai32 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix483 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .A0 (
          nx1183), .A1 (RST), .A2 (nx7433), .B0 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx469), .B1 (nx1179)) ;
    inv01 ix1182 (.Y (nx1183), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_9)) ;
    oai32 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix493 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .A0 (
          nx1185), .A1 (RST), .A2 (nx7433), .B0 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx477), .B1 (nx1179)) ;
    inv01 ix1184 (.Y (nx1185), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_10)) ;
    oai32 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix503 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .A0 (
          nx1187), .A1 (RST), .A2 (nx7433), .B0 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx485), .B1 (nx1179)) ;
    inv01 ix1186 (.Y (nx1187), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_11)) ;
    oai32 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix513 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .A0 (
          nx1189), .A1 (RST), .A2 (nx7433), .B0 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx493), .B1 (nx1179)) ;
    inv01 ix1188 (.Y (nx1189), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_12)) ;
    oai32 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix523 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .A0 (
          nx1191), .A1 (RST), .A2 (nx7433), .B0 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx501), .B1 (nx1179)) ;
    inv01 ix1190 (.Y (nx1191), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_13)) ;
    oai32 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix533 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .A0 (
          nx1193), .A1 (RST), .A2 (nx7435), .B0 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx509), .B1 (nx1195)) ;
    inv01 ix1192 (.Y (nx1193), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_14)) ;
    inv01 ix1194 (.Y (nx1195), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566)) ;
    oai32 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix543 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .A0 (
          nx1197), .A1 (RST), .A2 (nx7435), .B0 (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_nx517), .B1 (nx1195)) ;
    inv01 ix1196 (.Y (nx1197), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_15)) ;
    oai32 CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix553 (.Y (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .A0 (
          nx1199), .A1 (RST), .A2 (nx7435), .B0 (nx997), .B1 (nx1195)) ;
    inv01 ix1198 (.Y (nx1199), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_16)) ;
    nand02_2x CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix633 (.Y (
              nx1163), .A0 (nx7339), .A1 (nx7435)) ;
    nand02_2x CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix635 (.Y (
              nx1179), .A0 (nx7339), .A1 (nx7435)) ;
    mux21 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix404 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx403), .A0 (nx1201), .A1 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_2), .S0 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx395)) ;
    inv01 ix1200 (.Y (nx1201), .A (CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx391)) ;
    mux21 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix414 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx413), .A0 (nx1203), .A1 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_3), .S0 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx405)) ;
    inv01 ix1202 (.Y (nx1203), .A (CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx403)) ;
    mux21 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix424 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx423), .A0 (nx1205), .A1 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_4), .S0 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx415)) ;
    inv01 ix1204 (.Y (nx1205), .A (CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx413)) ;
    mux21 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix434 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx433), .A0 (nx1207), .A1 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_5), .S0 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx425)) ;
    inv01 ix1206 (.Y (nx1207), .A (CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx423)) ;
    mux21 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix444 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx443), .A0 (nx1209), .A1 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_6), .S0 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx435)) ;
    inv01 ix1208 (.Y (nx1209), .A (CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx433)) ;
    mux21 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix454 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx453), .A0 (nx1211), .A1 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_7), .S0 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx445)) ;
    inv01 ix1210 (.Y (nx1211), .A (CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx443)) ;
    mux21 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix462 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx461), .A0 (nx1213), .A1 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_8), .S0 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx455)) ;
    inv01 ix1212 (.Y (nx1213), .A (CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx453)) ;
    mux21 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix468 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx467), .A0 (nx1215), .A1 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_9), .S0 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx463)) ;
    inv01 ix1214 (.Y (nx1215), .A (CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx461)) ;
    mux21 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix476 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx475), .A0 (nx1217), .A1 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_10), .S0 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx471)) ;
    inv01 ix1216 (.Y (nx1217), .A (CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx467)) ;
    mux21 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix484 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx483), .A0 (nx1219), .A1 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_11), .S0 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx479)) ;
    inv01 ix1218 (.Y (nx1219), .A (CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx475)) ;
    mux21 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix492 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx491), .A0 (nx1221), .A1 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_12), .S0 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx487)) ;
    inv01 ix1220 (.Y (nx1221), .A (CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx483)) ;
    mux21 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix500 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx499), .A0 (nx1223), .A1 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_13), .S0 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx495)) ;
    inv01 ix1222 (.Y (nx1223), .A (CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx491)) ;
    mux21 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix508 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx507), .A0 (nx1225), .A1 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_14), .S0 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx503)) ;
    inv01 ix1224 (.Y (nx1225), .A (CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx499)) ;
    mux21 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix516 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx515), .A0 (nx1227), .A1 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_15), .S0 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx511)) ;
    inv01 ix1226 (.Y (nx1227), .A (CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx507)) ;
    mux21 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix161 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_1), .A0 (nx1229), .A1 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx379), .S0 (nx7439)) ;
    inv01 ix1228 (.Y (nx1229), .A (CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_1)) ;
    mux21 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix181 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_2), .A0 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx387), .A1 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx389), .S0 (nx7439)) ;
    mux21 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix201 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_3), .A0 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx399), .A1 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx401), .S0 (nx7439)) ;
    mux21 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix221 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_4), .A0 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx409), .A1 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx411), .S0 (nx7439)) ;
    mux21 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix241 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_5), .A0 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx419), .A1 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx421), .S0 (nx7439)) ;
    mux21 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix261 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_6), .A0 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx429), .A1 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx431), .S0 (nx7439)) ;
    mux21 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix281 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_7), .A0 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx439), .A1 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx441), .S0 (nx7439)) ;
    mux21 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix301 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_8), .A0 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx449), .A1 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx451), .S0 (nx7441)) ;
    mux21 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix321 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_9), .A0 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx469), .A1 (nx1231), .S0 (nx7441)) ;
    inv01 ix1230 (.Y (nx1231), .A (CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx316)) ;
    mux21 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix341 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_10), .A0 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx477), .A1 (nx1233), .S0 (nx7441)) ;
    inv01 ix1232 (.Y (nx1233), .A (CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx336)) ;
    mux21 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix361 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_11), .A0 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx485), .A1 (nx1235), .S0 (nx7441)) ;
    inv01 ix1234 (.Y (nx1235), .A (CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx356)) ;
    mux21 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix381 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_12), .A0 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx493), .A1 (nx1237), .S0 (nx7441)) ;
    inv01 ix1236 (.Y (nx1237), .A (CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx376)) ;
    mux21 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix401 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_13), .A0 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx501), .A1 (nx1239), .S0 (nx7441)) ;
    inv01 ix1238 (.Y (nx1239), .A (CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx396)) ;
    mux21 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix421 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_14), .A0 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx509), .A1 (nx1241), .S0 (nx7441)) ;
    inv01 ix1240 (.Y (nx1241), .A (CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx416)) ;
    mux21 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix441 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_15), .A0 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx517), .A1 (nx1243), .S0 (nx7443)) ;
    inv01 ix1242 (.Y (nx1243), .A (CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx436)) ;
    mux21 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_ix461 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_16), .A0 (nx1245), 
          .A1 (nx1247), .S0 (nx7443)) ;
    inv01 ix1244 (.Y (nx1245), .A (CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothP_16)
          ) ;
    inv01 ix1246 (.Y (nx1247), .A (CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx456)) ;
    nor02_2x CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix81 (.Y (
             CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx80), .A0 (Instr), .A1 (
             nx7305)) ;
    nor02_2x CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix319 (.Y (
             CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642), .A0 (
             CALCULATOR_Start_dup_1154), .A1 (
             CALCULATOR_CalculatingBooth_dup_1146)) ;
    nor02_2x CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix85 (.Y (
             CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_0), .A0 (
             nx7453), .A1 (nx1249)) ;
    inv01 ix1248 (.Y (nx1249), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_1)) ;
    mux21 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix125 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_1), .A0 (
          nx1251), .A1 (nx1253), .S0 (nx7453)) ;
    inv01 ix1250 (.Y (nx1251), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_2)) ;
    inv01 ix1252 (.Y (nx1253), .A (CacheWindow_0__2__0)) ;
    mux21 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix133 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_2), .A0 (
          nx1255), .A1 (nx1257), .S0 (nx7453)) ;
    inv01 ix1254 (.Y (nx1255), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_3)) ;
    inv01 ix1256 (.Y (nx1257), .A (CacheWindow_0__2__1)) ;
    mux21 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix141 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_3), .A0 (
          nx1259), .A1 (nx1261), .S0 (nx7453)) ;
    inv01 ix1258 (.Y (nx1259), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_4)) ;
    inv01 ix1260 (.Y (nx1261), .A (CacheWindow_0__2__2)) ;
    mux21 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix149 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_4), .A0 (
          nx1263), .A1 (nx1265), .S0 (nx7453)) ;
    inv01 ix1262 (.Y (nx1263), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_5)) ;
    inv01 ix1264 (.Y (nx1265), .A (CacheWindow_0__2__3)) ;
    mux21 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix157 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_5), .A0 (
          nx1267), .A1 (nx1269), .S0 (nx7453)) ;
    inv01 ix1266 (.Y (nx1267), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_6)) ;
    inv01 ix1268 (.Y (nx1269), .A (CacheWindow_0__2__4)) ;
    mux21 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix165 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_6), .A0 (
          nx1271), .A1 (nx1273), .S0 (nx7453)) ;
    inv01 ix1270 (.Y (nx1271), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_7)) ;
    inv01 ix1272 (.Y (nx1273), .A (CacheWindow_0__2__5)) ;
    mux21 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix173 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_7), .A0 (
          nx1275), .A1 (nx1277), .S0 (nx7455)) ;
    inv01 ix1274 (.Y (nx1275), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_8)) ;
    inv01 ix1276 (.Y (nx1277), .A (CacheWindow_0__2__6)) ;
    mux21 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix181 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_8), .A0 (
          nx1279), .A1 (nx1281), .S0 (nx7455)) ;
    inv01 ix1278 (.Y (nx1279), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_9)) ;
    inv01 ix1280 (.Y (nx1281), .A (CacheWindow_0__2__7)) ;
    nor02_2x CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix89 (.Y (
             CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_9), .A0 (
             nx7455), .A1 (nx1283)) ;
    inv01 ix1282 (.Y (nx1283), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_10)) ;
    nor02_2x CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix93 (.Y (
             CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_10), .A0 (
             nx7455), .A1 (nx1285)) ;
    inv01 ix1284 (.Y (nx1285), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_11)) ;
    nor02_2x CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix97 (.Y (
             CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_11), .A0 (
             nx7455), .A1 (nx1287)) ;
    inv01 ix1286 (.Y (nx1287), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_12)) ;
    nor02_2x CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix101 (.Y (
             CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_12), .A0 (
             nx7455), .A1 (nx1289)) ;
    inv01 ix1288 (.Y (nx1289), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_13)) ;
    nor02_2x CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix105 (.Y (
             CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_13), .A0 (
             nx7455), .A1 (nx1291)) ;
    inv01 ix1290 (.Y (nx1291), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_14)) ;
    nor02_2x CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix109 (.Y (
             CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_14), .A0 (
             nx7457), .A1 (nx1293)) ;
    inv01 ix1292 (.Y (nx1293), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_15)) ;
    nor02_2x CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix113 (.Y (
             CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_15), .A0 (
             nx7457), .A1 (nx1295)) ;
    inv01 ix1294 (.Y (nx1295), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_16)) ;
    nor02_2x CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix117 (.Y (
             CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_16), .A0 (
             nx7457), .A1 (nx1295)) ;
    mux21 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix189 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothOperand_0), .A0 (nx1297), .A1 (
          nx1299), .S0 (nx7445)) ;
    inv01 ix1296 (.Y (nx1297), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_0)) ;
    inv01 ix1298 (.Y (nx1299), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_0)) ;
    mux21 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix197 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothOperand_1), .A0 (nx1301), .A1 (
          nx1303), .S0 (nx7445)) ;
    inv01 ix1300 (.Y (nx1301), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_1)) ;
    inv01 ix1302 (.Y (nx1303), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_1)) ;
    mux21 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix205 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothOperand_2), .A0 (nx1305), .A1 (
          nx1307), .S0 (nx7445)) ;
    inv01 ix1304 (.Y (nx1305), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_2)) ;
    inv01 ix1306 (.Y (nx1307), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_2)) ;
    mux21 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix213 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothOperand_3), .A0 (nx1309), .A1 (
          nx1311), .S0 (nx7445)) ;
    inv01 ix1308 (.Y (nx1309), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_3)) ;
    inv01 ix1310 (.Y (nx1311), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_3)) ;
    mux21 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix221 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothOperand_4), .A0 (nx1313), .A1 (
          nx1315), .S0 (nx7445)) ;
    inv01 ix1312 (.Y (nx1313), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_4)) ;
    inv01 ix1314 (.Y (nx1315), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_4)) ;
    mux21 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix229 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothOperand_5), .A0 (nx1317), .A1 (
          nx1319), .S0 (nx7447)) ;
    inv01 ix1316 (.Y (nx1317), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_5)) ;
    inv01 ix1318 (.Y (nx1319), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_5)) ;
    mux21 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix237 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothOperand_6), .A0 (nx1321), .A1 (
          nx1323), .S0 (nx7447)) ;
    inv01 ix1320 (.Y (nx1321), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_6)) ;
    inv01 ix1322 (.Y (nx1323), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_6)) ;
    mux21 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix245 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothOperand_7), .A0 (nx1325), .A1 (
          nx1327), .S0 (nx7447)) ;
    inv01 ix1324 (.Y (nx1325), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_7)) ;
    inv01 ix1326 (.Y (nx1327), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_7)) ;
    mux21 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix253 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothOperand_8), .A0 (nx1329), .A1 (
          nx1331), .S0 (nx7447)) ;
    inv01 ix1328 (.Y (nx1329), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_8)) ;
    inv01 ix1330 (.Y (nx1331), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_8)) ;
    mux21 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix261 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothOperand_9), .A0 (nx1333), .A1 (
          nx1335), .S0 (nx7447)) ;
    inv01 ix1332 (.Y (nx1333), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_9)) ;
    inv01 ix1334 (.Y (nx1335), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_9)) ;
    mux21 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix269 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothOperand_10), .A0 (nx1337), .A1 (
          nx1339), .S0 (nx7447)) ;
    inv01 ix1336 (.Y (nx1337), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_10)) ;
    inv01 ix1338 (.Y (nx1339), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_10)) ;
    mux21 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix277 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothOperand_11), .A0 (nx1341), .A1 (
          nx1343), .S0 (nx7447)) ;
    inv01 ix1340 (.Y (nx1341), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_11)) ;
    inv01 ix1342 (.Y (nx1343), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_11)) ;
    mux21 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix285 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothOperand_12), .A0 (nx1345), .A1 (
          nx1347), .S0 (nx7449)) ;
    inv01 ix1344 (.Y (nx1345), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_12)) ;
    inv01 ix1346 (.Y (nx1347), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_12)) ;
    mux21 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix293 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothOperand_13), .A0 (nx1349), .A1 (
          nx1351), .S0 (nx7449)) ;
    inv01 ix1348 (.Y (nx1349), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_13)) ;
    inv01 ix1350 (.Y (nx1351), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_13)) ;
    mux21 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix301 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothOperand_14), .A0 (nx1353), .A1 (
          nx1355), .S0 (nx7449)) ;
    inv01 ix1352 (.Y (nx1353), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_14)) ;
    inv01 ix1354 (.Y (nx1355), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_14)) ;
    mux21 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix309 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothOperand_15), .A0 (nx1357), .A1 (
          nx1359), .S0 (nx7449)) ;
    inv01 ix1356 (.Y (nx1357), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_15)) ;
    inv01 ix1358 (.Y (nx1359), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_15)) ;
    mux21 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix317 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BoothOperand_16), .A0 (nx1361), .A1 (
          nx1363), .S0 (nx7449)) ;
    inv01 ix1360 (.Y (nx1361), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_16)) ;
    inv01 ix1362 (.Y (nx1363), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_16)) ;
    xnor2 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix321 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_AddPToBoothOperand), .A0 (nx7449), .A1 (
          nx1229)) ;
    oai32 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix393 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .A0 (
          nx8491), .A1 (RST), .A2 (nx7459), .B0 (nx1299), .B1 (nx1367)) ;
    oai32 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix403 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .A0 (
          nx8491), .A1 (RST), .A2 (nx7459), .B0 (nx1303), .B1 (nx1367)) ;
    oai32 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix413 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .A0 (
          nx8491), .A1 (RST), .A2 (nx7459), .B0 (nx1307), .B1 (nx1367)) ;
    oai32 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix423 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .A0 (
          nx8491), .A1 (RST), .A2 (nx7459), .B0 (nx1311), .B1 (nx1367)) ;
    oai32 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix433 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .A0 (
          nx8491), .A1 (RST), .A2 (nx7459), .B0 (nx1315), .B1 (nx1367)) ;
    oai32 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix443 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .A0 (
          nx8491), .A1 (RST), .A2 (nx7459), .B0 (nx1319), .B1 (nx1367)) ;
    oai32 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix453 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .A0 (
          nx8491), .A1 (RST), .A2 (nx7461), .B0 (nx1323), .B1 (nx1367)) ;
    oai32 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix463 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .A0 (
          nx8493), .A1 (RST), .A2 (nx7461), .B0 (nx1327), .B1 (nx1369)) ;
    oai32 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix473 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .A0 (
          nx8493), .A1 (RST), .A2 (nx7461), .B0 (nx1331), .B1 (nx1369)) ;
    oai32 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix483 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .A0 (
          nx1371), .A1 (RST), .A2 (nx7461), .B0 (nx1335), .B1 (nx1369)) ;
    inv01 ix1370 (.Y (nx1371), .A (CacheFilter_0__2__0)) ;
    oai32 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix493 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .A0 (
          nx1373), .A1 (RST), .A2 (nx7461), .B0 (nx1339), .B1 (nx1369)) ;
    inv01 ix1372 (.Y (nx1373), .A (CacheFilter_0__2__1)) ;
    oai32 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix503 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .A0 (
          nx1375), .A1 (RST), .A2 (nx7461), .B0 (nx1343), .B1 (nx1369)) ;
    inv01 ix1374 (.Y (nx1375), .A (CacheFilter_0__2__2)) ;
    oai32 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix513 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .A0 (
          nx1377), .A1 (RST), .A2 (nx7461), .B0 (nx1347), .B1 (nx1369)) ;
    inv01 ix1376 (.Y (nx1377), .A (CacheFilter_0__2__3)) ;
    oai32 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix523 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .A0 (
          nx1379), .A1 (RST), .A2 (nx7463), .B0 (nx1351), .B1 (nx1369)) ;
    inv01 ix1378 (.Y (nx1379), .A (CacheFilter_0__2__4)) ;
    oai32 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix533 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .A0 (
          nx1381), .A1 (RST), .A2 (nx7463), .B0 (nx1355), .B1 (nx1383)) ;
    inv01 ix1380 (.Y (nx1381), .A (CacheFilter_0__2__5)) ;
    inv01 ix1382 (.Y (nx1383), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566)) ;
    oai32 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix543 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .A0 (
          nx1385), .A1 (RST), .A2 (nx7463), .B0 (nx1359), .B1 (nx1383)) ;
    inv01 ix1384 (.Y (nx1385), .A (CacheFilter_0__2__6)) ;
    oai32 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix553 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .A0 (
          nx1387), .A1 (RST), .A2 (nx7463), .B0 (nx1363), .B1 (nx1383)) ;
    inv01 ix1386 (.Y (nx1387), .A (CacheFilter_0__2__7)) ;
    nand02_2x CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix633 (.Y (
              nx1367), .A0 (nx7339), .A1 (nx7463)) ;
    nand02_2x CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix635 (.Y (
              nx1369), .A0 (nx7341), .A1 (nx7463)) ;
    oai32 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix393 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .A0 (
          nx8493), .A1 (RST), .A2 (nx7465), .B0 (nx1297), .B1 (nx1389)) ;
    oai32 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix403 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .A0 (
          nx8493), .A1 (RST), .A2 (nx7465), .B0 (nx1301), .B1 (nx1389)) ;
    oai32 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix413 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .A0 (
          nx8493), .A1 (RST), .A2 (nx7465), .B0 (nx1305), .B1 (nx1389)) ;
    oai32 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix423 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .A0 (
          nx8493), .A1 (RST), .A2 (nx7465), .B0 (nx1309), .B1 (nx1389)) ;
    oai32 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix433 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .A0 (
          nx8493), .A1 (RST), .A2 (nx7465), .B0 (nx1313), .B1 (nx1389)) ;
    oai32 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix443 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .A0 (
          nx8495), .A1 (RST), .A2 (nx7465), .B0 (nx1317), .B1 (nx1389)) ;
    oai32 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix453 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .A0 (
          nx8495), .A1 (RST), .A2 (nx7467), .B0 (nx1321), .B1 (nx1389)) ;
    oai32 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix463 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .A0 (
          nx8495), .A1 (RST), .A2 (nx7467), .B0 (nx1325), .B1 (nx1391)) ;
    oai32 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix473 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .A0 (
          nx8495), .A1 (RST), .A2 (nx7467), .B0 (nx1329), .B1 (nx1391)) ;
    oai32 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix483 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .A0 (
          nx1371), .A1 (RST), .A2 (nx7467), .B0 (nx1333), .B1 (nx1391)) ;
    oai32 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix493 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .A0 (
          nx1393), .A1 (RST), .A2 (nx7467), .B0 (nx1337), .B1 (nx1391)) ;
    inv01 ix1392 (.Y (nx1393), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_10)) ;
    oai32 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix503 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .A0 (
          nx1395), .A1 (RST), .A2 (nx7467), .B0 (nx1341), .B1 (nx1391)) ;
    inv01 ix1394 (.Y (nx1395), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_11)) ;
    oai32 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix513 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .A0 (
          nx1397), .A1 (RST), .A2 (nx7467), .B0 (nx1345), .B1 (nx1391)) ;
    inv01 ix1396 (.Y (nx1397), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_12)) ;
    oai32 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix523 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .A0 (
          nx1399), .A1 (RST), .A2 (nx7469), .B0 (nx1349), .B1 (nx1391)) ;
    inv01 ix1398 (.Y (nx1399), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_13)) ;
    oai32 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix533 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .A0 (
          nx1401), .A1 (RST), .A2 (nx7469), .B0 (nx1353), .B1 (nx1403)) ;
    inv01 ix1400 (.Y (nx1401), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_14)) ;
    inv01 ix1402 (.Y (nx1403), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566)) ;
    oai32 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix543 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .A0 (
          nx1405), .A1 (RST), .A2 (nx7469), .B0 (nx1357), .B1 (nx1403)) ;
    inv01 ix1404 (.Y (nx1405), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_15)) ;
    oai32 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix553 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .A0 (
          nx1407), .A1 (RST), .A2 (nx7469), .B0 (nx1361), .B1 (nx1403)) ;
    inv01 ix1406 (.Y (nx1407), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_16)) ;
    nand02_2x CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix633 (.Y (
              nx1389), .A0 (nx7341), .A1 (nx7469)) ;
    nand02_2x CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix635 (.Y (
              nx1391), .A0 (nx7341), .A1 (nx7469)) ;
    oai32 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix393 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .A0 (
          nx1409), .A1 (RST), .A2 (nx7471), .B0 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx384), .B1 (nx1411)) ;
    inv01 ix1408 (.Y (nx1409), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_0)) ;
    oai32 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix403 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .A0 (
          nx1413), .A1 (RST), .A2 (nx7471), .B0 (nx1229), .B1 (nx1411)) ;
    inv01 ix1412 (.Y (nx1413), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_1)) ;
    oai32 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix413 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .A0 (
          nx1415), .A1 (RST), .A2 (nx7471), .B0 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx387), .B1 (nx1411)) ;
    inv01 ix1414 (.Y (nx1415), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_2)) ;
    oai32 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix423 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .A0 (
          nx1417), .A1 (RST), .A2 (nx7471), .B0 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx399), .B1 (nx1411)) ;
    inv01 ix1416 (.Y (nx1417), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_3)) ;
    oai32 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix433 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .A0 (
          nx1419), .A1 (RST), .A2 (nx7471), .B0 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx409), .B1 (nx1411)) ;
    inv01 ix1418 (.Y (nx1419), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_4)) ;
    oai32 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix443 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .A0 (
          nx1421), .A1 (RST), .A2 (nx7471), .B0 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx419), .B1 (nx1411)) ;
    inv01 ix1420 (.Y (nx1421), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_5)) ;
    oai32 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix453 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .A0 (
          nx1423), .A1 (RST), .A2 (nx7471), .B0 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx429), .B1 (nx1411)) ;
    inv01 ix1422 (.Y (nx1423), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_6)) ;
    oai32 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix463 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .A0 (
          nx1425), .A1 (RST), .A2 (nx7473), .B0 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx439), .B1 (nx1427)) ;
    inv01 ix1424 (.Y (nx1425), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_7)) ;
    oai32 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix473 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .A0 (
          nx1429), .A1 (RST), .A2 (nx7473), .B0 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx449), .B1 (nx1427)) ;
    inv01 ix1428 (.Y (nx1429), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_8)) ;
    oai32 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix483 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .A0 (
          nx1431), .A1 (RST), .A2 (nx7473), .B0 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx469), .B1 (nx1427)) ;
    inv01 ix1430 (.Y (nx1431), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_9)) ;
    oai32 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix493 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .A0 (
          nx1433), .A1 (RST), .A2 (nx7473), .B0 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx477), .B1 (nx1427)) ;
    inv01 ix1432 (.Y (nx1433), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_10)) ;
    oai32 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix503 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .A0 (
          nx1435), .A1 (RST), .A2 (nx7473), .B0 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx485), .B1 (nx1427)) ;
    inv01 ix1434 (.Y (nx1435), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_11)) ;
    oai32 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix513 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .A0 (
          nx1437), .A1 (RST), .A2 (nx7473), .B0 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx493), .B1 (nx1427)) ;
    inv01 ix1436 (.Y (nx1437), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_12)) ;
    oai32 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix523 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .A0 (
          nx1439), .A1 (RST), .A2 (nx7473), .B0 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx501), .B1 (nx1427)) ;
    inv01 ix1438 (.Y (nx1439), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_13)) ;
    oai32 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix533 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .A0 (
          nx1441), .A1 (RST), .A2 (nx7475), .B0 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx509), .B1 (nx1443)) ;
    inv01 ix1440 (.Y (nx1441), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_14)) ;
    inv01 ix1442 (.Y (nx1443), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566)) ;
    oai32 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix543 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .A0 (
          nx1445), .A1 (RST), .A2 (nx7475), .B0 (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_nx517), .B1 (nx1443)) ;
    inv01 ix1444 (.Y (nx1445), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_15)) ;
    oai32 CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix553 (.Y (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .A0 (
          nx1447), .A1 (RST), .A2 (nx7475), .B0 (nx1245), .B1 (nx1443)) ;
    inv01 ix1446 (.Y (nx1447), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_16)) ;
    nand02_2x CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix633 (.Y (
              nx1411), .A0 (nx7341), .A1 (nx7475)) ;
    nand02_2x CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix635 (.Y (
              nx1427), .A0 (nx7341), .A1 (nx7475)) ;
    mux21 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix404 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx403), .A0 (nx1449), .A1 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_2), .S0 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx395)) ;
    inv01 ix1448 (.Y (nx1449), .A (CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx391)) ;
    mux21 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix414 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx413), .A0 (nx1451), .A1 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_3), .S0 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx405)) ;
    inv01 ix1450 (.Y (nx1451), .A (CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx403)) ;
    mux21 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix424 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx423), .A0 (nx1453), .A1 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_4), .S0 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx415)) ;
    inv01 ix1452 (.Y (nx1453), .A (CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx413)) ;
    mux21 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix434 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx433), .A0 (nx1455), .A1 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_5), .S0 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx425)) ;
    inv01 ix1454 (.Y (nx1455), .A (CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx423)) ;
    mux21 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix444 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx443), .A0 (nx1457), .A1 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_6), .S0 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx435)) ;
    inv01 ix1456 (.Y (nx1457), .A (CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx433)) ;
    mux21 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix454 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx453), .A0 (nx1459), .A1 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_7), .S0 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx445)) ;
    inv01 ix1458 (.Y (nx1459), .A (CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx443)) ;
    mux21 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix462 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx461), .A0 (nx1461), .A1 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_8), .S0 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx455)) ;
    inv01 ix1460 (.Y (nx1461), .A (CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx453)) ;
    mux21 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix468 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx467), .A0 (nx1463), .A1 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_9), .S0 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx463)) ;
    inv01 ix1462 (.Y (nx1463), .A (CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx461)) ;
    mux21 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix476 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx475), .A0 (nx1465), .A1 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_10), .S0 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx471)) ;
    inv01 ix1464 (.Y (nx1465), .A (CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx467)) ;
    mux21 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix484 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx483), .A0 (nx1467), .A1 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_11), .S0 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx479)) ;
    inv01 ix1466 (.Y (nx1467), .A (CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx475)) ;
    mux21 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix492 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx491), .A0 (nx1469), .A1 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_12), .S0 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx487)) ;
    inv01 ix1468 (.Y (nx1469), .A (CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx483)) ;
    mux21 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix500 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx499), .A0 (nx1471), .A1 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_13), .S0 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx495)) ;
    inv01 ix1470 (.Y (nx1471), .A (CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx491)) ;
    mux21 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix508 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx507), .A0 (nx1473), .A1 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_14), .S0 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx503)) ;
    inv01 ix1472 (.Y (nx1473), .A (CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx499)) ;
    mux21 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix516 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx515), .A0 (nx1475), .A1 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_15), .S0 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx511)) ;
    inv01 ix1474 (.Y (nx1475), .A (CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx507)) ;
    mux21 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix161 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_1), .A0 (nx1477), .A1 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx379), .S0 (nx7479)) ;
    inv01 ix1476 (.Y (nx1477), .A (CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_1)) ;
    mux21 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix181 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_2), .A0 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx387), .A1 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx389), .S0 (nx7479)) ;
    mux21 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix201 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_3), .A0 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx399), .A1 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx401), .S0 (nx7479)) ;
    mux21 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix221 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_4), .A0 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx409), .A1 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx411), .S0 (nx7479)) ;
    mux21 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix241 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_5), .A0 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx419), .A1 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx421), .S0 (nx7479)) ;
    mux21 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix261 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_6), .A0 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx429), .A1 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx431), .S0 (nx7479)) ;
    mux21 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix281 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_7), .A0 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx439), .A1 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx441), .S0 (nx7479)) ;
    mux21 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix301 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_8), .A0 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx449), .A1 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx451), .S0 (nx7481)) ;
    mux21 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix321 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_9), .A0 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx469), .A1 (nx1479), .S0 (nx7481)) ;
    inv01 ix1478 (.Y (nx1479), .A (CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx316)) ;
    mux21 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix341 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_10), .A0 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx477), .A1 (nx1481), .S0 (nx7481)) ;
    inv01 ix1480 (.Y (nx1481), .A (CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx336)) ;
    mux21 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix361 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_11), .A0 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx485), .A1 (nx1483), .S0 (nx7481)) ;
    inv01 ix1482 (.Y (nx1483), .A (CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx356)) ;
    mux21 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix381 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_12), .A0 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx493), .A1 (nx1485), .S0 (nx7481)) ;
    inv01 ix1484 (.Y (nx1485), .A (CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx376)) ;
    mux21 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix401 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_13), .A0 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx501), .A1 (nx1487), .S0 (nx7481)) ;
    inv01 ix1486 (.Y (nx1487), .A (CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx396)) ;
    mux21 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix421 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_14), .A0 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx509), .A1 (nx1489), .S0 (nx7481)) ;
    inv01 ix1488 (.Y (nx1489), .A (CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx416)) ;
    mux21 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix441 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_15), .A0 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx517), .A1 (nx1491), .S0 (nx7483)) ;
    inv01 ix1490 (.Y (nx1491), .A (CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx436)) ;
    mux21 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_ix461 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_16), .A0 (nx1493), 
          .A1 (nx1495), .S0 (nx7483)) ;
    inv01 ix1492 (.Y (nx1493), .A (CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothP_16)
          ) ;
    inv01 ix1494 (.Y (nx1495), .A (CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx456)) ;
    nor02_2x CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix81 (.Y (
             CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx80), .A0 (Instr), .A1 (
             CALCULATOR_nx1111)) ;
    nor02_2x CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix319 (.Y (
             CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642), .A0 (
             CALCULATOR_Start_dup_1159), .A1 (
             CALCULATOR_CalculatingBooth_dup_1146)) ;
    nor02_2x CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix85 (.Y (
             CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_0), .A0 (
             nx7493), .A1 (nx1497)) ;
    inv01 ix1496 (.Y (nx1497), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_1)) ;
    mux21 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix125 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_1), .A0 (
          nx1499), .A1 (nx1501), .S0 (nx7493)) ;
    inv01 ix1498 (.Y (nx1499), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_2)) ;
    inv01 ix1500 (.Y (nx1501), .A (CacheWindow_0__3__0)) ;
    mux21 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix133 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_2), .A0 (
          nx1503), .A1 (nx1505), .S0 (nx7493)) ;
    inv01 ix1502 (.Y (nx1503), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_3)) ;
    inv01 ix1504 (.Y (nx1505), .A (CacheWindow_0__3__1)) ;
    mux21 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix141 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_3), .A0 (
          nx1507), .A1 (nx1509), .S0 (nx7493)) ;
    inv01 ix1506 (.Y (nx1507), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_4)) ;
    inv01 ix1508 (.Y (nx1509), .A (CacheWindow_0__3__2)) ;
    mux21 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix149 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_4), .A0 (
          nx1511), .A1 (nx1513), .S0 (nx7493)) ;
    inv01 ix1510 (.Y (nx1511), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_5)) ;
    inv01 ix1512 (.Y (nx1513), .A (CacheWindow_0__3__3)) ;
    mux21 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix157 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_5), .A0 (
          nx1515), .A1 (nx1517), .S0 (nx7493)) ;
    inv01 ix1514 (.Y (nx1515), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_6)) ;
    inv01 ix1516 (.Y (nx1517), .A (CacheWindow_0__3__4)) ;
    mux21 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix165 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_6), .A0 (
          nx1519), .A1 (nx1521), .S0 (nx7493)) ;
    inv01 ix1518 (.Y (nx1519), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_7)) ;
    inv01 ix1520 (.Y (nx1521), .A (CacheWindow_0__3__5)) ;
    mux21 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix173 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_7), .A0 (
          nx1523), .A1 (nx1525), .S0 (nx7495)) ;
    inv01 ix1522 (.Y (nx1523), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_8)) ;
    inv01 ix1524 (.Y (nx1525), .A (CacheWindow_0__3__6)) ;
    mux21 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix181 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_8), .A0 (
          nx1527), .A1 (nx1529), .S0 (nx7495)) ;
    inv01 ix1526 (.Y (nx1527), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_9)) ;
    inv01 ix1528 (.Y (nx1529), .A (CacheWindow_0__3__7)) ;
    nor02_2x CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix89 (.Y (
             CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_9), .A0 (
             nx7495), .A1 (nx1531)) ;
    inv01 ix1530 (.Y (nx1531), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_10)) ;
    nor02_2x CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix93 (.Y (
             CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_10), .A0 (
             nx7495), .A1 (nx1533)) ;
    inv01 ix1532 (.Y (nx1533), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_11)) ;
    nor02_2x CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix97 (.Y (
             CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_11), .A0 (
             nx7495), .A1 (nx1535)) ;
    inv01 ix1534 (.Y (nx1535), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_12)) ;
    nor02_2x CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix101 (.Y (
             CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_12), .A0 (
             nx7495), .A1 (nx1537)) ;
    inv01 ix1536 (.Y (nx1537), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_13)) ;
    nor02_2x CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix105 (.Y (
             CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_13), .A0 (
             nx7495), .A1 (nx1539)) ;
    inv01 ix1538 (.Y (nx1539), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_14)) ;
    nor02_2x CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix109 (.Y (
             CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_14), .A0 (
             nx7497), .A1 (nx1541)) ;
    inv01 ix1540 (.Y (nx1541), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_15)) ;
    nor02_2x CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix113 (.Y (
             CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_15), .A0 (
             nx7497), .A1 (nx1543)) ;
    inv01 ix1542 (.Y (nx1543), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_16)) ;
    nor02_2x CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix117 (.Y (
             CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_16), .A0 (
             nx7497), .A1 (nx1543)) ;
    mux21 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix189 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothOperand_0), .A0 (nx1545), .A1 (
          nx1547), .S0 (nx7485)) ;
    inv01 ix1544 (.Y (nx1545), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_0)) ;
    inv01 ix1546 (.Y (nx1547), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_0)) ;
    mux21 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix197 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothOperand_1), .A0 (nx1549), .A1 (
          nx1551), .S0 (nx7485)) ;
    inv01 ix1548 (.Y (nx1549), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_1)) ;
    inv01 ix1550 (.Y (nx1551), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_1)) ;
    mux21 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix205 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothOperand_2), .A0 (nx1553), .A1 (
          nx1555), .S0 (nx7485)) ;
    inv01 ix1552 (.Y (nx1553), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_2)) ;
    inv01 ix1554 (.Y (nx1555), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_2)) ;
    mux21 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix213 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothOperand_3), .A0 (nx1557), .A1 (
          nx1559), .S0 (nx7485)) ;
    inv01 ix1556 (.Y (nx1557), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_3)) ;
    inv01 ix1558 (.Y (nx1559), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_3)) ;
    mux21 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix221 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothOperand_4), .A0 (nx1561), .A1 (
          nx1563), .S0 (nx7485)) ;
    inv01 ix1560 (.Y (nx1561), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_4)) ;
    inv01 ix1562 (.Y (nx1563), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_4)) ;
    mux21 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix229 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothOperand_5), .A0 (nx1565), .A1 (
          nx1567), .S0 (nx7487)) ;
    inv01 ix1564 (.Y (nx1565), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_5)) ;
    inv01 ix1566 (.Y (nx1567), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_5)) ;
    mux21 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix237 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothOperand_6), .A0 (nx1569), .A1 (
          nx1571), .S0 (nx7487)) ;
    inv01 ix1568 (.Y (nx1569), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_6)) ;
    inv01 ix1570 (.Y (nx1571), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_6)) ;
    mux21 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix245 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothOperand_7), .A0 (nx1573), .A1 (
          nx1575), .S0 (nx7487)) ;
    inv01 ix1572 (.Y (nx1573), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_7)) ;
    inv01 ix1574 (.Y (nx1575), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_7)) ;
    mux21 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix253 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothOperand_8), .A0 (nx1577), .A1 (
          nx1579), .S0 (nx7487)) ;
    inv01 ix1576 (.Y (nx1577), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_8)) ;
    inv01 ix1578 (.Y (nx1579), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_8)) ;
    mux21 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix261 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothOperand_9), .A0 (nx1581), .A1 (
          nx1583), .S0 (nx7487)) ;
    inv01 ix1580 (.Y (nx1581), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_9)) ;
    inv01 ix1582 (.Y (nx1583), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_9)) ;
    mux21 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix269 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothOperand_10), .A0 (nx1585), .A1 (
          nx1587), .S0 (nx7487)) ;
    inv01 ix1584 (.Y (nx1585), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_10)) ;
    inv01 ix1586 (.Y (nx1587), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_10)) ;
    mux21 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix277 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothOperand_11), .A0 (nx1589), .A1 (
          nx1591), .S0 (nx7487)) ;
    inv01 ix1588 (.Y (nx1589), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_11)) ;
    inv01 ix1590 (.Y (nx1591), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_11)) ;
    mux21 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix285 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothOperand_12), .A0 (nx1593), .A1 (
          nx1595), .S0 (nx7489)) ;
    inv01 ix1592 (.Y (nx1593), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_12)) ;
    inv01 ix1594 (.Y (nx1595), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_12)) ;
    mux21 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix293 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothOperand_13), .A0 (nx1597), .A1 (
          nx1599), .S0 (nx7489)) ;
    inv01 ix1596 (.Y (nx1597), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_13)) ;
    inv01 ix1598 (.Y (nx1599), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_13)) ;
    mux21 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix301 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothOperand_14), .A0 (nx1601), .A1 (
          nx1603), .S0 (nx7489)) ;
    inv01 ix1600 (.Y (nx1601), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_14)) ;
    inv01 ix1602 (.Y (nx1603), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_14)) ;
    mux21 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix309 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothOperand_15), .A0 (nx1605), .A1 (
          nx1607), .S0 (nx7489)) ;
    inv01 ix1604 (.Y (nx1605), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_15)) ;
    inv01 ix1606 (.Y (nx1607), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_15)) ;
    mux21 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix317 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BoothOperand_16), .A0 (nx1609), .A1 (
          nx1611), .S0 (nx7489)) ;
    inv01 ix1608 (.Y (nx1609), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_16)) ;
    inv01 ix1610 (.Y (nx1611), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_16)) ;
    xnor2 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix321 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_AddPToBoothOperand), .A0 (nx7489), .A1 (
          nx1477)) ;
    oai32 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix393 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .A0 (
          nx8497), .A1 (RST), .A2 (nx7499), .B0 (nx1547), .B1 (nx1615)) ;
    oai32 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix403 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .A0 (
          nx8497), .A1 (RST), .A2 (nx7499), .B0 (nx1551), .B1 (nx1615)) ;
    oai32 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix413 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .A0 (
          nx8497), .A1 (RST), .A2 (nx7499), .B0 (nx1555), .B1 (nx1615)) ;
    oai32 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix423 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .A0 (
          nx8497), .A1 (RST), .A2 (nx7499), .B0 (nx1559), .B1 (nx1615)) ;
    oai32 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix433 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .A0 (
          nx8497), .A1 (RST), .A2 (nx7499), .B0 (nx1563), .B1 (nx1615)) ;
    oai32 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix443 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .A0 (
          nx8497), .A1 (RST), .A2 (nx7499), .B0 (nx1567), .B1 (nx1615)) ;
    oai32 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix453 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .A0 (
          nx8497), .A1 (RST), .A2 (nx7501), .B0 (nx1571), .B1 (nx1615)) ;
    oai32 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix463 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .A0 (
          nx8499), .A1 (RST), .A2 (nx7501), .B0 (nx1575), .B1 (nx1617)) ;
    oai32 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix473 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .A0 (
          nx8499), .A1 (RST), .A2 (nx7501), .B0 (nx1579), .B1 (nx1617)) ;
    oai32 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix483 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .A0 (
          nx1619), .A1 (RST), .A2 (nx7501), .B0 (nx1583), .B1 (nx1617)) ;
    inv01 ix1618 (.Y (nx1619), .A (CacheFilter_0__3__0)) ;
    oai32 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix493 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .A0 (
          nx1621), .A1 (RST), .A2 (nx7501), .B0 (nx1587), .B1 (nx1617)) ;
    inv01 ix1620 (.Y (nx1621), .A (CacheFilter_0__3__1)) ;
    oai32 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix503 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .A0 (
          nx1623), .A1 (RST), .A2 (nx7501), .B0 (nx1591), .B1 (nx1617)) ;
    inv01 ix1622 (.Y (nx1623), .A (CacheFilter_0__3__2)) ;
    oai32 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix513 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .A0 (
          nx1625), .A1 (RST), .A2 (nx7501), .B0 (nx1595), .B1 (nx1617)) ;
    inv01 ix1624 (.Y (nx1625), .A (CacheFilter_0__3__3)) ;
    oai32 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix523 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .A0 (
          nx1627), .A1 (RST), .A2 (nx7503), .B0 (nx1599), .B1 (nx1617)) ;
    inv01 ix1626 (.Y (nx1627), .A (CacheFilter_0__3__4)) ;
    oai32 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix533 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .A0 (
          nx1629), .A1 (RST), .A2 (nx7503), .B0 (nx1603), .B1 (nx1631)) ;
    inv01 ix1628 (.Y (nx1629), .A (CacheFilter_0__3__5)) ;
    inv01 ix1630 (.Y (nx1631), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566)) ;
    oai32 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix543 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .A0 (
          nx1633), .A1 (RST), .A2 (nx7503), .B0 (nx1607), .B1 (nx1631)) ;
    inv01 ix1632 (.Y (nx1633), .A (CacheFilter_0__3__6)) ;
    oai32 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix553 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .A0 (
          nx1635), .A1 (RST), .A2 (nx7503), .B0 (nx1611), .B1 (nx1631)) ;
    inv01 ix1634 (.Y (nx1635), .A (CacheFilter_0__3__7)) ;
    nand02_2x CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix633 (.Y (
              nx1615), .A0 (nx7341), .A1 (nx7503)) ;
    nand02_2x CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix635 (.Y (
              nx1617), .A0 (nx7341), .A1 (nx7503)) ;
    oai32 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix393 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .A0 (
          nx8499), .A1 (RST), .A2 (nx7505), .B0 (nx1545), .B1 (nx1637)) ;
    oai32 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix403 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .A0 (
          nx8499), .A1 (RST), .A2 (nx7505), .B0 (nx1549), .B1 (nx1637)) ;
    oai32 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix413 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .A0 (
          nx8499), .A1 (RST), .A2 (nx7505), .B0 (nx1553), .B1 (nx1637)) ;
    oai32 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix423 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .A0 (
          nx8499), .A1 (RST), .A2 (nx7505), .B0 (nx1557), .B1 (nx1637)) ;
    oai32 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix433 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .A0 (
          nx8499), .A1 (RST), .A2 (nx7505), .B0 (nx1561), .B1 (nx1637)) ;
    oai32 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix443 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .A0 (
          nx8501), .A1 (RST), .A2 (nx7505), .B0 (nx1565), .B1 (nx1637)) ;
    oai32 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix453 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .A0 (
          nx8501), .A1 (RST), .A2 (nx7507), .B0 (nx1569), .B1 (nx1637)) ;
    oai32 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix463 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .A0 (
          nx8501), .A1 (RST), .A2 (nx7507), .B0 (nx1573), .B1 (nx1639)) ;
    oai32 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix473 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .A0 (
          nx8501), .A1 (RST), .A2 (nx7507), .B0 (nx1577), .B1 (nx1639)) ;
    oai32 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix483 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .A0 (
          nx1619), .A1 (RST), .A2 (nx7507), .B0 (nx1581), .B1 (nx1639)) ;
    oai32 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix493 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .A0 (
          nx1641), .A1 (RST), .A2 (nx7507), .B0 (nx1585), .B1 (nx1639)) ;
    inv01 ix1640 (.Y (nx1641), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_10)) ;
    oai32 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix503 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .A0 (
          nx1643), .A1 (RST), .A2 (nx7507), .B0 (nx1589), .B1 (nx1639)) ;
    inv01 ix1642 (.Y (nx1643), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_11)) ;
    oai32 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix513 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .A0 (
          nx1645), .A1 (RST), .A2 (nx7507), .B0 (nx1593), .B1 (nx1639)) ;
    inv01 ix1644 (.Y (nx1645), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_12)) ;
    oai32 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix523 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .A0 (
          nx1647), .A1 (RST), .A2 (nx7509), .B0 (nx1597), .B1 (nx1639)) ;
    inv01 ix1646 (.Y (nx1647), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_13)) ;
    oai32 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix533 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .A0 (
          nx1649), .A1 (RST), .A2 (nx7509), .B0 (nx1601), .B1 (nx1651)) ;
    inv01 ix1648 (.Y (nx1649), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_14)) ;
    inv01 ix1650 (.Y (nx1651), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566)) ;
    oai32 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix543 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .A0 (
          nx1653), .A1 (RST), .A2 (nx7509), .B0 (nx1605), .B1 (nx1651)) ;
    inv01 ix1652 (.Y (nx1653), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_15)) ;
    oai32 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix553 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .A0 (
          nx1655), .A1 (RST), .A2 (nx7509), .B0 (nx1609), .B1 (nx1651)) ;
    inv01 ix1654 (.Y (nx1655), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_16)) ;
    nand02_2x CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix633 (.Y (
              nx1637), .A0 (nx7343), .A1 (nx7509)) ;
    nand02_2x CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix635 (.Y (
              nx1639), .A0 (nx7343), .A1 (nx7509)) ;
    oai32 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix393 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .A0 (
          nx1657), .A1 (RST), .A2 (nx7511), .B0 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx384), .B1 (nx1659)) ;
    inv01 ix1656 (.Y (nx1657), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_0)) ;
    oai32 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix403 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .A0 (
          nx1661), .A1 (RST), .A2 (nx7511), .B0 (nx1477), .B1 (nx1659)) ;
    inv01 ix1660 (.Y (nx1661), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_1)) ;
    oai32 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix413 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .A0 (
          nx1663), .A1 (RST), .A2 (nx7511), .B0 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx387), .B1 (nx1659)) ;
    inv01 ix1662 (.Y (nx1663), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_2)) ;
    oai32 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix423 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .A0 (
          nx1665), .A1 (RST), .A2 (nx7511), .B0 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx399), .B1 (nx1659)) ;
    inv01 ix1664 (.Y (nx1665), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_3)) ;
    oai32 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix433 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .A0 (
          nx1667), .A1 (RST), .A2 (nx7511), .B0 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx409), .B1 (nx1659)) ;
    inv01 ix1666 (.Y (nx1667), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_4)) ;
    oai32 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix443 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .A0 (
          nx1669), .A1 (RST), .A2 (nx7511), .B0 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx419), .B1 (nx1659)) ;
    inv01 ix1668 (.Y (nx1669), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_5)) ;
    oai32 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix453 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .A0 (
          nx1671), .A1 (RST), .A2 (nx7511), .B0 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx429), .B1 (nx1659)) ;
    inv01 ix1670 (.Y (nx1671), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_6)) ;
    oai32 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix463 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .A0 (
          nx1673), .A1 (RST), .A2 (nx7513), .B0 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx439), .B1 (nx1675)) ;
    inv01 ix1672 (.Y (nx1673), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_7)) ;
    oai32 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix473 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .A0 (
          nx1677), .A1 (RST), .A2 (nx7513), .B0 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx449), .B1 (nx1675)) ;
    inv01 ix1676 (.Y (nx1677), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_8)) ;
    oai32 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix483 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .A0 (
          nx1679), .A1 (RST), .A2 (nx7513), .B0 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx469), .B1 (nx1675)) ;
    inv01 ix1678 (.Y (nx1679), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_9)) ;
    oai32 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix493 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .A0 (
          nx1681), .A1 (RST), .A2 (nx7513), .B0 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx477), .B1 (nx1675)) ;
    inv01 ix1680 (.Y (nx1681), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_10)) ;
    oai32 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix503 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .A0 (
          nx1683), .A1 (RST), .A2 (nx7513), .B0 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx485), .B1 (nx1675)) ;
    inv01 ix1682 (.Y (nx1683), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_11)) ;
    oai32 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix513 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .A0 (
          nx1685), .A1 (RST), .A2 (nx7513), .B0 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx493), .B1 (nx1675)) ;
    inv01 ix1684 (.Y (nx1685), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_12)) ;
    oai32 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix523 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .A0 (
          nx1687), .A1 (RST), .A2 (nx7513), .B0 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx501), .B1 (nx1675)) ;
    inv01 ix1686 (.Y (nx1687), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_13)) ;
    oai32 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix533 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .A0 (
          nx1689), .A1 (RST), .A2 (nx7515), .B0 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx509), .B1 (nx1691)) ;
    inv01 ix1688 (.Y (nx1689), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_14)) ;
    inv01 ix1690 (.Y (nx1691), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566)) ;
    oai32 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix543 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .A0 (
          nx1693), .A1 (RST), .A2 (nx7515), .B0 (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_nx517), .B1 (nx1691)) ;
    inv01 ix1692 (.Y (nx1693), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_15)) ;
    oai32 CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix553 (.Y (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .A0 (
          nx1695), .A1 (RST), .A2 (nx7515), .B0 (nx1493), .B1 (nx1691)) ;
    inv01 ix1694 (.Y (nx1695), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_16)) ;
    nand02_2x CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix633 (.Y (
              nx1659), .A0 (nx7343), .A1 (nx7515)) ;
    nand02_2x CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix635 (.Y (
              nx1675), .A0 (nx7343), .A1 (nx7515)) ;
    mux21 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix404 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx403), .A0 (nx1697), .A1 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_2), .S0 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx395)) ;
    inv01 ix1696 (.Y (nx1697), .A (CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx391)) ;
    mux21 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix414 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx413), .A0 (nx1699), .A1 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_3), .S0 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx405)) ;
    inv01 ix1698 (.Y (nx1699), .A (CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx403)) ;
    mux21 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix424 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx423), .A0 (nx1701), .A1 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_4), .S0 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx415)) ;
    inv01 ix1700 (.Y (nx1701), .A (CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx413)) ;
    mux21 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix434 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx433), .A0 (nx1703), .A1 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_5), .S0 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx425)) ;
    inv01 ix1702 (.Y (nx1703), .A (CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx423)) ;
    mux21 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix444 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx443), .A0 (nx1705), .A1 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_6), .S0 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx435)) ;
    inv01 ix1704 (.Y (nx1705), .A (CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx433)) ;
    mux21 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix454 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx453), .A0 (nx1707), .A1 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_7), .S0 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx445)) ;
    inv01 ix1706 (.Y (nx1707), .A (CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx443)) ;
    mux21 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix462 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx461), .A0 (nx1709), .A1 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_8), .S0 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx455)) ;
    inv01 ix1708 (.Y (nx1709), .A (CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx453)) ;
    mux21 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix468 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx467), .A0 (nx1711), .A1 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_9), .S0 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx463)) ;
    inv01 ix1710 (.Y (nx1711), .A (CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx461)) ;
    mux21 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix476 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx475), .A0 (nx1713), .A1 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_10), .S0 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx471)) ;
    inv01 ix1712 (.Y (nx1713), .A (CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx467)) ;
    mux21 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix484 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx483), .A0 (nx1715), .A1 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_11), .S0 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx479)) ;
    inv01 ix1714 (.Y (nx1715), .A (CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx475)) ;
    mux21 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix492 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx491), .A0 (nx1717), .A1 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_12), .S0 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx487)) ;
    inv01 ix1716 (.Y (nx1717), .A (CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx483)) ;
    mux21 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix500 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx499), .A0 (nx1719), .A1 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_13), .S0 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx495)) ;
    inv01 ix1718 (.Y (nx1719), .A (CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx491)) ;
    mux21 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix508 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx507), .A0 (nx1721), .A1 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_14), .S0 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx503)) ;
    inv01 ix1720 (.Y (nx1721), .A (CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx499)) ;
    mux21 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix516 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx515), .A0 (nx1723), .A1 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_15), .S0 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx511)) ;
    inv01 ix1722 (.Y (nx1723), .A (CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx507)) ;
    mux21 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix161 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_1), .A0 (nx1725), .A1 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx379), .S0 (nx7519)) ;
    inv01 ix1724 (.Y (nx1725), .A (CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_1)) ;
    mux21 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix181 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_2), .A0 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx387), .A1 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx389), .S0 (nx7519)) ;
    mux21 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix201 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_3), .A0 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx399), .A1 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx401), .S0 (nx7519)) ;
    mux21 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix221 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_4), .A0 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx409), .A1 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx411), .S0 (nx7519)) ;
    mux21 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix241 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_5), .A0 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx419), .A1 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx421), .S0 (nx7519)) ;
    mux21 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix261 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_6), .A0 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx429), .A1 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx431), .S0 (nx7519)) ;
    mux21 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix281 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_7), .A0 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx439), .A1 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx441), .S0 (nx7519)) ;
    mux21 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix301 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_8), .A0 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx449), .A1 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx451), .S0 (nx7521)) ;
    mux21 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix321 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_9), .A0 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx469), .A1 (nx1727), .S0 (nx7521)) ;
    inv01 ix1726 (.Y (nx1727), .A (CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx316)) ;
    mux21 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix341 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_10), .A0 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx477), .A1 (nx1729), .S0 (nx7521)) ;
    inv01 ix1728 (.Y (nx1729), .A (CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx336)) ;
    mux21 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix361 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_11), .A0 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx485), .A1 (nx1731), .S0 (nx7521)) ;
    inv01 ix1730 (.Y (nx1731), .A (CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx356)) ;
    mux21 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix381 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_12), .A0 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx493), .A1 (nx1733), .S0 (nx7521)) ;
    inv01 ix1732 (.Y (nx1733), .A (CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx376)) ;
    mux21 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix401 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_13), .A0 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx501), .A1 (nx1735), .S0 (nx7521)) ;
    inv01 ix1734 (.Y (nx1735), .A (CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx396)) ;
    mux21 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix421 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_14), .A0 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx509), .A1 (nx1737), .S0 (nx7521)) ;
    inv01 ix1736 (.Y (nx1737), .A (CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx416)) ;
    mux21 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix441 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_15), .A0 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx517), .A1 (nx1739), .S0 (nx7523)) ;
    inv01 ix1738 (.Y (nx1739), .A (CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx436)) ;
    mux21 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_ix461 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_16), .A0 (nx1741), 
          .A1 (nx1743), .S0 (nx7523)) ;
    inv01 ix1740 (.Y (nx1741), .A (CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothP_16)
          ) ;
    inv01 ix1742 (.Y (nx1743), .A (CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx456)) ;
    nor02_2x CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix81 (.Y (
             CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx80), .A0 (Instr), .A1 (
             CALCULATOR_nx1111)) ;
    nor02_2x CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix319 (.Y (
             CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642), .A0 (
             CALCULATOR_Start_dup_1164), .A1 (
             CALCULATOR_CalculatingBooth_dup_1146)) ;
    nor02_2x CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix85 (.Y (
             CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_0), .A0 (
             nx7533), .A1 (nx1745)) ;
    inv01 ix1744 (.Y (nx1745), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_1)) ;
    mux21 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix125 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_1), .A0 (
          nx1747), .A1 (nx1749), .S0 (nx7533)) ;
    inv01 ix1746 (.Y (nx1747), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_2)) ;
    inv01 ix1748 (.Y (nx1749), .A (CacheWindow_0__4__0)) ;
    mux21 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix133 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_2), .A0 (
          nx1751), .A1 (nx1753), .S0 (nx7533)) ;
    inv01 ix1750 (.Y (nx1751), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_3)) ;
    inv01 ix1752 (.Y (nx1753), .A (CacheWindow_0__4__1)) ;
    mux21 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix141 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_3), .A0 (
          nx1755), .A1 (nx1757), .S0 (nx7533)) ;
    inv01 ix1754 (.Y (nx1755), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_4)) ;
    inv01 ix1756 (.Y (nx1757), .A (CacheWindow_0__4__2)) ;
    mux21 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix149 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_4), .A0 (
          nx1759), .A1 (nx1761), .S0 (nx7533)) ;
    inv01 ix1758 (.Y (nx1759), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_5)) ;
    inv01 ix1760 (.Y (nx1761), .A (CacheWindow_0__4__3)) ;
    mux21 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix157 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_5), .A0 (
          nx1763), .A1 (nx1765), .S0 (nx7533)) ;
    inv01 ix1762 (.Y (nx1763), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_6)) ;
    inv01 ix1764 (.Y (nx1765), .A (CacheWindow_0__4__4)) ;
    mux21 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix165 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_6), .A0 (
          nx1767), .A1 (nx1769), .S0 (nx7533)) ;
    inv01 ix1766 (.Y (nx1767), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_7)) ;
    inv01 ix1768 (.Y (nx1769), .A (CacheWindow_0__4__5)) ;
    mux21 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix173 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_7), .A0 (
          nx1771), .A1 (nx1773), .S0 (nx7535)) ;
    inv01 ix1770 (.Y (nx1771), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_8)) ;
    inv01 ix1772 (.Y (nx1773), .A (CacheWindow_0__4__6)) ;
    mux21 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix181 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_8), .A0 (
          nx1775), .A1 (nx1777), .S0 (nx7535)) ;
    inv01 ix1774 (.Y (nx1775), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_9)) ;
    inv01 ix1776 (.Y (nx1777), .A (CacheWindow_0__4__7)) ;
    nor02_2x CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix89 (.Y (
             CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_9), .A0 (
             nx7535), .A1 (nx1779)) ;
    inv01 ix1778 (.Y (nx1779), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_10)) ;
    nor02_2x CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix93 (.Y (
             CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_10), .A0 (
             nx7535), .A1 (nx1781)) ;
    inv01 ix1780 (.Y (nx1781), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_11)) ;
    nor02_2x CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix97 (.Y (
             CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_11), .A0 (
             nx7535), .A1 (nx1783)) ;
    inv01 ix1782 (.Y (nx1783), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_12)) ;
    nor02_2x CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix101 (.Y (
             CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_12), .A0 (
             nx7535), .A1 (nx1785)) ;
    inv01 ix1784 (.Y (nx1785), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_13)) ;
    nor02_2x CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix105 (.Y (
             CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_13), .A0 (
             nx7535), .A1 (nx1787)) ;
    inv01 ix1786 (.Y (nx1787), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_14)) ;
    nor02_2x CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix109 (.Y (
             CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_14), .A0 (
             nx7537), .A1 (nx1789)) ;
    inv01 ix1788 (.Y (nx1789), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_15)) ;
    nor02_2x CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix113 (.Y (
             CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_15), .A0 (
             nx7537), .A1 (nx1791)) ;
    inv01 ix1790 (.Y (nx1791), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_16)) ;
    nor02_2x CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix117 (.Y (
             CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_16), .A0 (
             nx7537), .A1 (nx1791)) ;
    mux21 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix189 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothOperand_0), .A0 (nx1793), .A1 (
          nx1795), .S0 (nx7525)) ;
    inv01 ix1792 (.Y (nx1793), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_0)) ;
    inv01 ix1794 (.Y (nx1795), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_0)) ;
    mux21 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix197 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothOperand_1), .A0 (nx1797), .A1 (
          nx1799), .S0 (nx7525)) ;
    inv01 ix1796 (.Y (nx1797), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_1)) ;
    inv01 ix1798 (.Y (nx1799), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_1)) ;
    mux21 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix205 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothOperand_2), .A0 (nx1801), .A1 (
          nx1803), .S0 (nx7525)) ;
    inv01 ix1800 (.Y (nx1801), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_2)) ;
    inv01 ix1802 (.Y (nx1803), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_2)) ;
    mux21 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix213 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothOperand_3), .A0 (nx1805), .A1 (
          nx1807), .S0 (nx7525)) ;
    inv01 ix1804 (.Y (nx1805), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_3)) ;
    inv01 ix1806 (.Y (nx1807), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_3)) ;
    mux21 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix221 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothOperand_4), .A0 (nx1809), .A1 (
          nx1811), .S0 (nx7525)) ;
    inv01 ix1808 (.Y (nx1809), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_4)) ;
    inv01 ix1810 (.Y (nx1811), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_4)) ;
    mux21 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix229 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothOperand_5), .A0 (nx1813), .A1 (
          nx1815), .S0 (nx7527)) ;
    inv01 ix1812 (.Y (nx1813), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_5)) ;
    inv01 ix1814 (.Y (nx1815), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_5)) ;
    mux21 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix237 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothOperand_6), .A0 (nx1817), .A1 (
          nx1819), .S0 (nx7527)) ;
    inv01 ix1816 (.Y (nx1817), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_6)) ;
    inv01 ix1818 (.Y (nx1819), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_6)) ;
    mux21 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix245 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothOperand_7), .A0 (nx1821), .A1 (
          nx1823), .S0 (nx7527)) ;
    inv01 ix1820 (.Y (nx1821), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_7)) ;
    inv01 ix1822 (.Y (nx1823), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_7)) ;
    mux21 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix253 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothOperand_8), .A0 (nx1825), .A1 (
          nx1827), .S0 (nx7527)) ;
    inv01 ix1824 (.Y (nx1825), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_8)) ;
    inv01 ix1826 (.Y (nx1827), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_8)) ;
    mux21 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix261 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothOperand_9), .A0 (nx1829), .A1 (
          nx1831), .S0 (nx7527)) ;
    inv01 ix1828 (.Y (nx1829), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_9)) ;
    inv01 ix1830 (.Y (nx1831), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_9)) ;
    mux21 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix269 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothOperand_10), .A0 (nx1833), .A1 (
          nx1835), .S0 (nx7527)) ;
    inv01 ix1832 (.Y (nx1833), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_10)) ;
    inv01 ix1834 (.Y (nx1835), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_10)) ;
    mux21 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix277 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothOperand_11), .A0 (nx1837), .A1 (
          nx1839), .S0 (nx7527)) ;
    inv01 ix1836 (.Y (nx1837), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_11)) ;
    inv01 ix1838 (.Y (nx1839), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_11)) ;
    mux21 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix285 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothOperand_12), .A0 (nx1841), .A1 (
          nx1843), .S0 (nx7529)) ;
    inv01 ix1840 (.Y (nx1841), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_12)) ;
    inv01 ix1842 (.Y (nx1843), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_12)) ;
    mux21 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix293 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothOperand_13), .A0 (nx1845), .A1 (
          nx1847), .S0 (nx7529)) ;
    inv01 ix1844 (.Y (nx1845), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_13)) ;
    inv01 ix1846 (.Y (nx1847), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_13)) ;
    mux21 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix301 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothOperand_14), .A0 (nx1849), .A1 (
          nx1851), .S0 (nx7529)) ;
    inv01 ix1848 (.Y (nx1849), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_14)) ;
    inv01 ix1850 (.Y (nx1851), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_14)) ;
    mux21 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix309 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothOperand_15), .A0 (nx1853), .A1 (
          nx1855), .S0 (nx7529)) ;
    inv01 ix1852 (.Y (nx1853), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_15)) ;
    inv01 ix1854 (.Y (nx1855), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_15)) ;
    mux21 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix317 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BoothOperand_16), .A0 (nx1857), .A1 (
          nx1859), .S0 (nx7529)) ;
    inv01 ix1856 (.Y (nx1857), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_16)) ;
    inv01 ix1858 (.Y (nx1859), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_16)) ;
    xnor2 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix321 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_AddPToBoothOperand), .A0 (nx7529), .A1 (
          nx1725)) ;
    oai32 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix393 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .A0 (
          nx8503), .A1 (RST), .A2 (nx7539), .B0 (nx1795), .B1 (nx1863)) ;
    oai32 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix403 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .A0 (
          nx8503), .A1 (RST), .A2 (nx7539), .B0 (nx1799), .B1 (nx1863)) ;
    oai32 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix413 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .A0 (
          nx8503), .A1 (RST), .A2 (nx7539), .B0 (nx1803), .B1 (nx1863)) ;
    oai32 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix423 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .A0 (
          nx8503), .A1 (RST), .A2 (nx7539), .B0 (nx1807), .B1 (nx1863)) ;
    oai32 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix433 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .A0 (
          nx8503), .A1 (RST), .A2 (nx7539), .B0 (nx1811), .B1 (nx1863)) ;
    oai32 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix443 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .A0 (
          nx8503), .A1 (RST), .A2 (nx7539), .B0 (nx1815), .B1 (nx1863)) ;
    oai32 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix453 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .A0 (
          nx8503), .A1 (RST), .A2 (nx7541), .B0 (nx1819), .B1 (nx1863)) ;
    oai32 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix463 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .A0 (
          nx8505), .A1 (RST), .A2 (nx7541), .B0 (nx1823), .B1 (nx1865)) ;
    oai32 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix473 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .A0 (
          nx8505), .A1 (RST), .A2 (nx7541), .B0 (nx1827), .B1 (nx1865)) ;
    oai32 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix483 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .A0 (
          nx1867), .A1 (RST), .A2 (nx7541), .B0 (nx1831), .B1 (nx1865)) ;
    inv01 ix1866 (.Y (nx1867), .A (CacheFilter_0__4__0)) ;
    oai32 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix493 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .A0 (
          nx1869), .A1 (RST), .A2 (nx7541), .B0 (nx1835), .B1 (nx1865)) ;
    inv01 ix1868 (.Y (nx1869), .A (CacheFilter_0__4__1)) ;
    oai32 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix503 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .A0 (
          nx1871), .A1 (RST), .A2 (nx7541), .B0 (nx1839), .B1 (nx1865)) ;
    inv01 ix1870 (.Y (nx1871), .A (CacheFilter_0__4__2)) ;
    oai32 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix513 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .A0 (
          nx1873), .A1 (RST), .A2 (nx7541), .B0 (nx1843), .B1 (nx1865)) ;
    inv01 ix1872 (.Y (nx1873), .A (CacheFilter_0__4__3)) ;
    oai32 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix523 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .A0 (
          nx1875), .A1 (RST), .A2 (nx7543), .B0 (nx1847), .B1 (nx1865)) ;
    inv01 ix1874 (.Y (nx1875), .A (CacheFilter_0__4__4)) ;
    oai32 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix533 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .A0 (
          nx1877), .A1 (RST), .A2 (nx7543), .B0 (nx1851), .B1 (nx1879)) ;
    inv01 ix1876 (.Y (nx1877), .A (CacheFilter_0__4__5)) ;
    inv01 ix1878 (.Y (nx1879), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566)) ;
    oai32 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix543 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .A0 (
          nx1881), .A1 (RST), .A2 (nx7543), .B0 (nx1855), .B1 (nx1879)) ;
    inv01 ix1880 (.Y (nx1881), .A (CacheFilter_0__4__6)) ;
    oai32 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix553 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .A0 (
          nx1883), .A1 (RST), .A2 (nx7543), .B0 (nx1859), .B1 (nx1879)) ;
    inv01 ix1882 (.Y (nx1883), .A (CacheFilter_0__4__7)) ;
    nand02_2x CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix633 (.Y (
              nx1863), .A0 (nx7343), .A1 (nx7543)) ;
    nand02_2x CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix635 (.Y (
              nx1865), .A0 (nx7343), .A1 (nx7543)) ;
    oai32 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix393 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .A0 (
          nx8505), .A1 (RST), .A2 (nx7545), .B0 (nx1793), .B1 (nx1885)) ;
    oai32 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix403 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .A0 (
          nx8505), .A1 (RST), .A2 (nx7545), .B0 (nx1797), .B1 (nx1885)) ;
    oai32 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix413 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .A0 (
          nx8505), .A1 (RST), .A2 (nx7545), .B0 (nx1801), .B1 (nx1885)) ;
    oai32 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix423 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .A0 (
          nx8505), .A1 (RST), .A2 (nx7545), .B0 (nx1805), .B1 (nx1885)) ;
    oai32 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix433 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .A0 (
          nx8505), .A1 (RST), .A2 (nx7545), .B0 (nx1809), .B1 (nx1885)) ;
    oai32 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix443 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .A0 (
          nx8507), .A1 (RST), .A2 (nx7545), .B0 (nx1813), .B1 (nx1885)) ;
    oai32 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix453 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .A0 (
          nx8507), .A1 (RST), .A2 (nx7547), .B0 (nx1817), .B1 (nx1885)) ;
    oai32 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix463 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .A0 (
          nx8507), .A1 (RST), .A2 (nx7547), .B0 (nx1821), .B1 (nx1887)) ;
    oai32 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix473 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .A0 (
          nx8507), .A1 (RST), .A2 (nx7547), .B0 (nx1825), .B1 (nx1887)) ;
    oai32 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix483 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .A0 (
          nx1867), .A1 (RST), .A2 (nx7547), .B0 (nx1829), .B1 (nx1887)) ;
    oai32 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix493 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .A0 (
          nx1889), .A1 (RST), .A2 (nx7547), .B0 (nx1833), .B1 (nx1887)) ;
    inv01 ix1888 (.Y (nx1889), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_10)) ;
    oai32 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix503 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .A0 (
          nx1891), .A1 (RST), .A2 (nx7547), .B0 (nx1837), .B1 (nx1887)) ;
    inv01 ix1890 (.Y (nx1891), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_11)) ;
    oai32 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix513 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .A0 (
          nx1893), .A1 (RST), .A2 (nx7547), .B0 (nx1841), .B1 (nx1887)) ;
    inv01 ix1892 (.Y (nx1893), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_12)) ;
    oai32 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix523 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .A0 (
          nx1895), .A1 (RST), .A2 (nx7549), .B0 (nx1845), .B1 (nx1887)) ;
    inv01 ix1894 (.Y (nx1895), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_13)) ;
    oai32 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix533 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .A0 (
          nx1897), .A1 (RST), .A2 (nx7549), .B0 (nx1849), .B1 (nx1899)) ;
    inv01 ix1896 (.Y (nx1897), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_14)) ;
    inv01 ix1898 (.Y (nx1899), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566)) ;
    oai32 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix543 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .A0 (
          nx1901), .A1 (RST), .A2 (nx7549), .B0 (nx1853), .B1 (nx1899)) ;
    inv01 ix1900 (.Y (nx1901), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_15)) ;
    oai32 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix553 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .A0 (
          nx1903), .A1 (RST), .A2 (nx7549), .B0 (nx1857), .B1 (nx1899)) ;
    inv01 ix1902 (.Y (nx1903), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_16)) ;
    nand02_2x CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix633 (.Y (
              nx1885), .A0 (nx7343), .A1 (nx7549)) ;
    nand02_2x CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix635 (.Y (
              nx1887), .A0 (nx7345), .A1 (nx7549)) ;
    oai32 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix393 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .A0 (
          nx1905), .A1 (RST), .A2 (nx7551), .B0 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx384), .B1 (nx1907)) ;
    inv01 ix1904 (.Y (nx1905), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_0)) ;
    oai32 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix403 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .A0 (
          nx1909), .A1 (RST), .A2 (nx7551), .B0 (nx1725), .B1 (nx1907)) ;
    inv01 ix1908 (.Y (nx1909), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_1)) ;
    oai32 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix413 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .A0 (
          nx1911), .A1 (RST), .A2 (nx7551), .B0 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx387), .B1 (nx1907)) ;
    inv01 ix1910 (.Y (nx1911), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_2)) ;
    oai32 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix423 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .A0 (
          nx1913), .A1 (RST), .A2 (nx7551), .B0 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx399), .B1 (nx1907)) ;
    inv01 ix1912 (.Y (nx1913), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_3)) ;
    oai32 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix433 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .A0 (
          nx1915), .A1 (RST), .A2 (nx7551), .B0 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx409), .B1 (nx1907)) ;
    inv01 ix1914 (.Y (nx1915), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_4)) ;
    oai32 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix443 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .A0 (
          nx1917), .A1 (RST), .A2 (nx7551), .B0 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx419), .B1 (nx1907)) ;
    inv01 ix1916 (.Y (nx1917), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_5)) ;
    oai32 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix453 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .A0 (
          nx1919), .A1 (RST), .A2 (nx7551), .B0 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx429), .B1 (nx1907)) ;
    inv01 ix1918 (.Y (nx1919), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_6)) ;
    oai32 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix463 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .A0 (
          nx1921), .A1 (RST), .A2 (nx7553), .B0 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx439), .B1 (nx1923)) ;
    inv01 ix1920 (.Y (nx1921), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_7)) ;
    oai32 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix473 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .A0 (
          nx1925), .A1 (RST), .A2 (nx7553), .B0 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx449), .B1 (nx1923)) ;
    inv01 ix1924 (.Y (nx1925), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_8)) ;
    oai32 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix483 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .A0 (
          nx1927), .A1 (RST), .A2 (nx7553), .B0 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx469), .B1 (nx1923)) ;
    inv01 ix1926 (.Y (nx1927), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_9)) ;
    oai32 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix493 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .A0 (
          nx1929), .A1 (RST), .A2 (nx7553), .B0 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx477), .B1 (nx1923)) ;
    inv01 ix1928 (.Y (nx1929), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_10)) ;
    oai32 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix503 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .A0 (
          nx1931), .A1 (RST), .A2 (nx7553), .B0 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx485), .B1 (nx1923)) ;
    inv01 ix1930 (.Y (nx1931), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_11)) ;
    oai32 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix513 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .A0 (
          nx1933), .A1 (RST), .A2 (nx7553), .B0 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx493), .B1 (nx1923)) ;
    inv01 ix1932 (.Y (nx1933), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_12)) ;
    oai32 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix523 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .A0 (
          nx1935), .A1 (RST), .A2 (nx7553), .B0 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx501), .B1 (nx1923)) ;
    inv01 ix1934 (.Y (nx1935), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_13)) ;
    oai32 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix533 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .A0 (
          nx1937), .A1 (RST), .A2 (nx7555), .B0 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx509), .B1 (nx1939)) ;
    inv01 ix1936 (.Y (nx1937), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_14)) ;
    inv01 ix1938 (.Y (nx1939), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566)) ;
    oai32 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix543 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .A0 (
          nx1941), .A1 (RST), .A2 (nx7555), .B0 (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_nx517), .B1 (nx1939)) ;
    inv01 ix1940 (.Y (nx1941), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_15)) ;
    oai32 CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix553 (.Y (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .A0 (
          nx1943), .A1 (RST), .A2 (nx7555), .B0 (nx1741), .B1 (nx1939)) ;
    inv01 ix1942 (.Y (nx1943), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_16)) ;
    nand02_2x CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix633 (.Y (
              nx1907), .A0 (nx7345), .A1 (nx7555)) ;
    nand02_2x CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix635 (.Y (
              nx1923), .A0 (nx7345), .A1 (nx7555)) ;
    mux21 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix404 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx403), .A0 (nx1945), .A1 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_2), .S0 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx395)) ;
    inv01 ix1944 (.Y (nx1945), .A (CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx391)) ;
    mux21 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix414 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx413), .A0 (nx1947), .A1 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_3), .S0 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx405)) ;
    inv01 ix1946 (.Y (nx1947), .A (CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx403)) ;
    mux21 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix424 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx423), .A0 (nx1949), .A1 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_4), .S0 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx415)) ;
    inv01 ix1948 (.Y (nx1949), .A (CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx413)) ;
    mux21 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix434 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx433), .A0 (nx1951), .A1 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_5), .S0 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx425)) ;
    inv01 ix1950 (.Y (nx1951), .A (CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx423)) ;
    mux21 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix444 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx443), .A0 (nx1953), .A1 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_6), .S0 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx435)) ;
    inv01 ix1952 (.Y (nx1953), .A (CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx433)) ;
    mux21 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix454 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx453), .A0 (nx1955), .A1 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_7), .S0 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx445)) ;
    inv01 ix1954 (.Y (nx1955), .A (CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx443)) ;
    mux21 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix462 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx461), .A0 (nx1957), .A1 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_8), .S0 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx455)) ;
    inv01 ix1956 (.Y (nx1957), .A (CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx453)) ;
    mux21 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix468 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx467), .A0 (nx1959), .A1 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_9), .S0 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx463)) ;
    inv01 ix1958 (.Y (nx1959), .A (CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx461)) ;
    mux21 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix476 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx475), .A0 (nx1961), .A1 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_10), .S0 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx471)) ;
    inv01 ix1960 (.Y (nx1961), .A (CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx467)) ;
    mux21 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix484 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx483), .A0 (nx1963), .A1 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_11), .S0 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx479)) ;
    inv01 ix1962 (.Y (nx1963), .A (CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx475)) ;
    mux21 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix492 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx491), .A0 (nx1965), .A1 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_12), .S0 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx487)) ;
    inv01 ix1964 (.Y (nx1965), .A (CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx483)) ;
    mux21 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix500 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx499), .A0 (nx1967), .A1 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_13), .S0 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx495)) ;
    inv01 ix1966 (.Y (nx1967), .A (CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx491)) ;
    mux21 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix508 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx507), .A0 (nx1969), .A1 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_14), .S0 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx503)) ;
    inv01 ix1968 (.Y (nx1969), .A (CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx499)) ;
    mux21 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix516 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx515), .A0 (nx1971), .A1 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_15), .S0 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx511)) ;
    inv01 ix1970 (.Y (nx1971), .A (CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx507)) ;
    mux21 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix161 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_1), .A0 (nx1973), .A1 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx379), .S0 (nx7559)) ;
    inv01 ix1972 (.Y (nx1973), .A (CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_1)) ;
    mux21 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix181 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_2), .A0 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx387), .A1 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx389), .S0 (nx7559)) ;
    mux21 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix201 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_3), .A0 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx399), .A1 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx401), .S0 (nx7559)) ;
    mux21 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix221 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_4), .A0 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx409), .A1 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx411), .S0 (nx7559)) ;
    mux21 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix241 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_5), .A0 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx419), .A1 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx421), .S0 (nx7559)) ;
    mux21 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix261 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_6), .A0 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx429), .A1 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx431), .S0 (nx7559)) ;
    mux21 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix281 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_7), .A0 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx439), .A1 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx441), .S0 (nx7559)) ;
    mux21 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix301 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_8), .A0 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx449), .A1 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx451), .S0 (nx7561)) ;
    mux21 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix321 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_9), .A0 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx469), .A1 (nx1975), .S0 (nx7561)) ;
    inv01 ix1974 (.Y (nx1975), .A (CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx316)) ;
    mux21 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix341 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_10), .A0 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx477), .A1 (nx1977), .S0 (nx7561)) ;
    inv01 ix1976 (.Y (nx1977), .A (CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx336)) ;
    mux21 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix361 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_11), .A0 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx485), .A1 (nx1979), .S0 (nx7561)) ;
    inv01 ix1978 (.Y (nx1979), .A (CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx356)) ;
    mux21 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix381 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_12), .A0 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx493), .A1 (nx1981), .S0 (nx7561)) ;
    inv01 ix1980 (.Y (nx1981), .A (CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx376)) ;
    mux21 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix401 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_13), .A0 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx501), .A1 (nx1983), .S0 (nx7561)) ;
    inv01 ix1982 (.Y (nx1983), .A (CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx396)) ;
    mux21 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix421 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_14), .A0 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx509), .A1 (nx1985), .S0 (nx7561)) ;
    inv01 ix1984 (.Y (nx1985), .A (CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx416)) ;
    mux21 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix441 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_15), .A0 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx517), .A1 (nx1987), .S0 (nx7563)) ;
    inv01 ix1986 (.Y (nx1987), .A (CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx436)) ;
    mux21 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_ix461 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_16), .A0 (nx1989), 
          .A1 (nx1991), .S0 (nx7563)) ;
    inv01 ix1988 (.Y (nx1989), .A (CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothP_16)
          ) ;
    inv01 ix1990 (.Y (nx1991), .A (CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx456)) ;
    nor02_2x CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix81 (.Y (
             CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx80), .A0 (Instr), .A1 (
             CALCULATOR_nx1111)) ;
    nor02_2x CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix319 (.Y (
             CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642), .A0 (
             CALCULATOR_Start_dup_1169), .A1 (
             CALCULATOR_CalculatingBooth_dup_1146)) ;
    nor02_2x CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix85 (.Y (
             CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_0), .A0 (
             nx7573), .A1 (nx1993)) ;
    inv01 ix1992 (.Y (nx1993), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_1)) ;
    mux21 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix125 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_1), .A0 (
          nx1995), .A1 (nx1997), .S0 (nx7573)) ;
    inv01 ix1994 (.Y (nx1995), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_2)) ;
    inv01 ix1996 (.Y (nx1997), .A (CacheWindow_1__0__0)) ;
    mux21 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix133 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_2), .A0 (
          nx1999), .A1 (nx2001), .S0 (nx7573)) ;
    inv01 ix1998 (.Y (nx1999), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_3)) ;
    inv01 ix2000 (.Y (nx2001), .A (CacheWindow_1__0__1)) ;
    mux21 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix141 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_3), .A0 (
          nx2003), .A1 (nx2005), .S0 (nx7573)) ;
    inv01 ix2002 (.Y (nx2003), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_4)) ;
    inv01 ix2004 (.Y (nx2005), .A (CacheWindow_1__0__2)) ;
    mux21 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix149 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_4), .A0 (
          nx2007), .A1 (nx2009), .S0 (nx7573)) ;
    inv01 ix2006 (.Y (nx2007), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_5)) ;
    inv01 ix2008 (.Y (nx2009), .A (CacheWindow_1__0__3)) ;
    mux21 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix157 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_5), .A0 (
          nx2011), .A1 (nx2013), .S0 (nx7573)) ;
    inv01 ix2010 (.Y (nx2011), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_6)) ;
    inv01 ix2012 (.Y (nx2013), .A (CacheWindow_1__0__4)) ;
    mux21 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix165 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_6), .A0 (
          nx2015), .A1 (nx2017), .S0 (nx7573)) ;
    inv01 ix2014 (.Y (nx2015), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_7)) ;
    inv01 ix2016 (.Y (nx2017), .A (CacheWindow_1__0__5)) ;
    mux21 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix173 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_7), .A0 (
          nx2019), .A1 (nx2021), .S0 (nx7575)) ;
    inv01 ix2018 (.Y (nx2019), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_8)) ;
    inv01 ix2020 (.Y (nx2021), .A (CacheWindow_1__0__6)) ;
    mux21 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix181 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_8), .A0 (
          nx2023), .A1 (nx2025), .S0 (nx7575)) ;
    inv01 ix2022 (.Y (nx2023), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_9)) ;
    inv01 ix2024 (.Y (nx2025), .A (CacheWindow_1__0__7)) ;
    nor02_2x CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix89 (.Y (
             CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_9), .A0 (
             nx7575), .A1 (nx2027)) ;
    inv01 ix2026 (.Y (nx2027), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_10)) ;
    nor02_2x CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix93 (.Y (
             CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_10), .A0 (
             nx7575), .A1 (nx2029)) ;
    inv01 ix2028 (.Y (nx2029), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_11)) ;
    nor02_2x CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix97 (.Y (
             CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_11), .A0 (
             nx7575), .A1 (nx2031)) ;
    inv01 ix2030 (.Y (nx2031), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_12)) ;
    nor02_2x CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix101 (.Y (
             CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_12), .A0 (
             nx7575), .A1 (nx2033)) ;
    inv01 ix2032 (.Y (nx2033), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_13)) ;
    nor02_2x CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix105 (.Y (
             CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_13), .A0 (
             nx7575), .A1 (nx2035)) ;
    inv01 ix2034 (.Y (nx2035), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_14)) ;
    nor02_2x CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix109 (.Y (
             CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_14), .A0 (
             nx7577), .A1 (nx2037)) ;
    inv01 ix2036 (.Y (nx2037), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_15)) ;
    nor02_2x CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix113 (.Y (
             CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_15), .A0 (
             nx7577), .A1 (nx2039)) ;
    inv01 ix2038 (.Y (nx2039), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_16)) ;
    nor02_2x CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix117 (.Y (
             CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_16), .A0 (
             nx7577), .A1 (nx2039)) ;
    mux21 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix189 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothOperand_0), .A0 (nx2041), .A1 (
          nx2043), .S0 (nx7565)) ;
    inv01 ix2040 (.Y (nx2041), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_0)) ;
    inv01 ix2042 (.Y (nx2043), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_0)) ;
    mux21 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix197 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothOperand_1), .A0 (nx2045), .A1 (
          nx2047), .S0 (nx7565)) ;
    inv01 ix2044 (.Y (nx2045), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_1)) ;
    inv01 ix2046 (.Y (nx2047), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_1)) ;
    mux21 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix205 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothOperand_2), .A0 (nx2049), .A1 (
          nx2051), .S0 (nx7565)) ;
    inv01 ix2048 (.Y (nx2049), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_2)) ;
    inv01 ix2050 (.Y (nx2051), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_2)) ;
    mux21 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix213 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothOperand_3), .A0 (nx2053), .A1 (
          nx2055), .S0 (nx7565)) ;
    inv01 ix2052 (.Y (nx2053), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_3)) ;
    inv01 ix2054 (.Y (nx2055), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_3)) ;
    mux21 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix221 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothOperand_4), .A0 (nx2057), .A1 (
          nx2059), .S0 (nx7565)) ;
    inv01 ix2056 (.Y (nx2057), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_4)) ;
    inv01 ix2058 (.Y (nx2059), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_4)) ;
    mux21 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix229 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothOperand_5), .A0 (nx2061), .A1 (
          nx2063), .S0 (nx7567)) ;
    inv01 ix2060 (.Y (nx2061), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_5)) ;
    inv01 ix2062 (.Y (nx2063), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_5)) ;
    mux21 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix237 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothOperand_6), .A0 (nx2065), .A1 (
          nx2067), .S0 (nx7567)) ;
    inv01 ix2064 (.Y (nx2065), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_6)) ;
    inv01 ix2066 (.Y (nx2067), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_6)) ;
    mux21 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix245 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothOperand_7), .A0 (nx2069), .A1 (
          nx2071), .S0 (nx7567)) ;
    inv01 ix2068 (.Y (nx2069), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_7)) ;
    inv01 ix2070 (.Y (nx2071), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_7)) ;
    mux21 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix253 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothOperand_8), .A0 (nx2073), .A1 (
          nx2075), .S0 (nx7567)) ;
    inv01 ix2072 (.Y (nx2073), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_8)) ;
    inv01 ix2074 (.Y (nx2075), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_8)) ;
    mux21 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix261 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothOperand_9), .A0 (nx2077), .A1 (
          nx2079), .S0 (nx7567)) ;
    inv01 ix2076 (.Y (nx2077), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_9)) ;
    inv01 ix2078 (.Y (nx2079), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_9)) ;
    mux21 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix269 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothOperand_10), .A0 (nx2081), .A1 (
          nx2083), .S0 (nx7567)) ;
    inv01 ix2080 (.Y (nx2081), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_10)) ;
    inv01 ix2082 (.Y (nx2083), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_10)) ;
    mux21 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix277 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothOperand_11), .A0 (nx2085), .A1 (
          nx2087), .S0 (nx7567)) ;
    inv01 ix2084 (.Y (nx2085), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_11)) ;
    inv01 ix2086 (.Y (nx2087), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_11)) ;
    mux21 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix285 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothOperand_12), .A0 (nx2089), .A1 (
          nx2091), .S0 (nx7569)) ;
    inv01 ix2088 (.Y (nx2089), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_12)) ;
    inv01 ix2090 (.Y (nx2091), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_12)) ;
    mux21 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix293 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothOperand_13), .A0 (nx2093), .A1 (
          nx2095), .S0 (nx7569)) ;
    inv01 ix2092 (.Y (nx2093), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_13)) ;
    inv01 ix2094 (.Y (nx2095), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_13)) ;
    mux21 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix301 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothOperand_14), .A0 (nx2097), .A1 (
          nx2099), .S0 (nx7569)) ;
    inv01 ix2096 (.Y (nx2097), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_14)) ;
    inv01 ix2098 (.Y (nx2099), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_14)) ;
    mux21 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix309 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothOperand_15), .A0 (nx2101), .A1 (
          nx2103), .S0 (nx7569)) ;
    inv01 ix2100 (.Y (nx2101), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_15)) ;
    inv01 ix2102 (.Y (nx2103), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_15)) ;
    mux21 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix317 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BoothOperand_16), .A0 (nx2105), .A1 (
          nx2107), .S0 (nx7569)) ;
    inv01 ix2104 (.Y (nx2105), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_16)) ;
    inv01 ix2106 (.Y (nx2107), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_16)) ;
    xnor2 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix321 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_AddPToBoothOperand), .A0 (nx7569), .A1 (
          nx1973)) ;
    oai32 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix393 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .A0 (
          nx8509), .A1 (RST), .A2 (nx7579), .B0 (nx2043), .B1 (nx2111)) ;
    oai32 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix403 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .A0 (
          nx8509), .A1 (RST), .A2 (nx7579), .B0 (nx2047), .B1 (nx2111)) ;
    oai32 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix413 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .A0 (
          nx8509), .A1 (RST), .A2 (nx7579), .B0 (nx2051), .B1 (nx2111)) ;
    oai32 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix423 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .A0 (
          nx8509), .A1 (RST), .A2 (nx7579), .B0 (nx2055), .B1 (nx2111)) ;
    oai32 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix433 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .A0 (
          nx8509), .A1 (RST), .A2 (nx7579), .B0 (nx2059), .B1 (nx2111)) ;
    oai32 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix443 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .A0 (
          nx8509), .A1 (RST), .A2 (nx7579), .B0 (nx2063), .B1 (nx2111)) ;
    oai32 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix453 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .A0 (
          nx8509), .A1 (RST), .A2 (nx7581), .B0 (nx2067), .B1 (nx2111)) ;
    oai32 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix463 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .A0 (
          nx8511), .A1 (RST), .A2 (nx7581), .B0 (nx2071), .B1 (nx2113)) ;
    oai32 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix473 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .A0 (
          nx8511), .A1 (RST), .A2 (nx7581), .B0 (nx2075), .B1 (nx2113)) ;
    oai32 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix483 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .A0 (
          nx2115), .A1 (RST), .A2 (nx7581), .B0 (nx2079), .B1 (nx2113)) ;
    inv01 ix2114 (.Y (nx2115), .A (CacheFilter_1__0__0)) ;
    oai32 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix493 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .A0 (
          nx2117), .A1 (RST), .A2 (nx7581), .B0 (nx2083), .B1 (nx2113)) ;
    inv01 ix2116 (.Y (nx2117), .A (CacheFilter_1__0__1)) ;
    oai32 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix503 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .A0 (
          nx2119), .A1 (RST), .A2 (nx7581), .B0 (nx2087), .B1 (nx2113)) ;
    inv01 ix2118 (.Y (nx2119), .A (CacheFilter_1__0__2)) ;
    oai32 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix513 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .A0 (
          nx2121), .A1 (RST), .A2 (nx7581), .B0 (nx2091), .B1 (nx2113)) ;
    inv01 ix2120 (.Y (nx2121), .A (CacheFilter_1__0__3)) ;
    oai32 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix523 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .A0 (
          nx2123), .A1 (RST), .A2 (nx7583), .B0 (nx2095), .B1 (nx2113)) ;
    inv01 ix2122 (.Y (nx2123), .A (CacheFilter_1__0__4)) ;
    oai32 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix533 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .A0 (
          nx2125), .A1 (RST), .A2 (nx7583), .B0 (nx2099), .B1 (nx2127)) ;
    inv01 ix2124 (.Y (nx2125), .A (CacheFilter_1__0__5)) ;
    inv01 ix2126 (.Y (nx2127), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566)) ;
    oai32 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix543 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .A0 (
          nx2129), .A1 (RST), .A2 (nx7583), .B0 (nx2103), .B1 (nx2127)) ;
    inv01 ix2128 (.Y (nx2129), .A (CacheFilter_1__0__6)) ;
    oai32 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix553 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .A0 (
          nx2131), .A1 (RST), .A2 (nx7583), .B0 (nx2107), .B1 (nx2127)) ;
    inv01 ix2130 (.Y (nx2131), .A (CacheFilter_1__0__7)) ;
    nand02_2x CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix633 (.Y (
              nx2111), .A0 (nx7345), .A1 (nx7583)) ;
    nand02_2x CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix635 (.Y (
              nx2113), .A0 (nx7345), .A1 (nx7583)) ;
    oai32 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix393 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .A0 (
          nx8511), .A1 (RST), .A2 (nx7585), .B0 (nx2041), .B1 (nx2133)) ;
    oai32 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix403 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .A0 (
          nx8511), .A1 (RST), .A2 (nx7585), .B0 (nx2045), .B1 (nx2133)) ;
    oai32 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix413 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .A0 (
          nx8511), .A1 (RST), .A2 (nx7585), .B0 (nx2049), .B1 (nx2133)) ;
    oai32 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix423 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .A0 (
          nx8511), .A1 (RST), .A2 (nx7585), .B0 (nx2053), .B1 (nx2133)) ;
    oai32 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix433 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .A0 (
          nx8511), .A1 (RST), .A2 (nx7585), .B0 (nx2057), .B1 (nx2133)) ;
    oai32 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix443 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .A0 (
          nx8513), .A1 (RST), .A2 (nx7585), .B0 (nx2061), .B1 (nx2133)) ;
    oai32 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix453 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .A0 (
          nx8513), .A1 (RST), .A2 (nx7587), .B0 (nx2065), .B1 (nx2133)) ;
    oai32 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix463 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .A0 (
          nx8513), .A1 (RST), .A2 (nx7587), .B0 (nx2069), .B1 (nx2135)) ;
    oai32 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix473 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .A0 (
          nx8513), .A1 (RST), .A2 (nx7587), .B0 (nx2073), .B1 (nx2135)) ;
    oai32 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix483 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .A0 (
          nx2115), .A1 (RST), .A2 (nx7587), .B0 (nx2077), .B1 (nx2135)) ;
    oai32 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix493 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .A0 (
          nx2137), .A1 (RST), .A2 (nx7587), .B0 (nx2081), .B1 (nx2135)) ;
    inv01 ix2136 (.Y (nx2137), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_10)) ;
    oai32 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix503 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .A0 (
          nx2139), .A1 (RST), .A2 (nx7587), .B0 (nx2085), .B1 (nx2135)) ;
    inv01 ix2138 (.Y (nx2139), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_11)) ;
    oai32 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix513 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .A0 (
          nx2141), .A1 (RST), .A2 (nx7587), .B0 (nx2089), .B1 (nx2135)) ;
    inv01 ix2140 (.Y (nx2141), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_12)) ;
    oai32 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix523 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .A0 (
          nx2143), .A1 (RST), .A2 (nx7589), .B0 (nx2093), .B1 (nx2135)) ;
    inv01 ix2142 (.Y (nx2143), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_13)) ;
    oai32 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix533 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .A0 (
          nx2145), .A1 (RST), .A2 (nx7589), .B0 (nx2097), .B1 (nx2147)) ;
    inv01 ix2144 (.Y (nx2145), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_14)) ;
    inv01 ix2146 (.Y (nx2147), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566)) ;
    oai32 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix543 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .A0 (
          nx2149), .A1 (RST), .A2 (nx7589), .B0 (nx2101), .B1 (nx2147)) ;
    inv01 ix2148 (.Y (nx2149), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_15)) ;
    oai32 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix553 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .A0 (
          nx2151), .A1 (RST), .A2 (nx7589), .B0 (nx2105), .B1 (nx2147)) ;
    inv01 ix2150 (.Y (nx2151), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_16)) ;
    nand02_2x CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix633 (.Y (
              nx2133), .A0 (nx7345), .A1 (nx7589)) ;
    nand02_2x CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix635 (.Y (
              nx2135), .A0 (nx7345), .A1 (nx7589)) ;
    oai32 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix393 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .A0 (
          nx2153), .A1 (RST), .A2 (nx7591), .B0 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx384), .B1 (nx2155)) ;
    inv01 ix2152 (.Y (nx2153), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_0)) ;
    oai32 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix403 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .A0 (
          nx2157), .A1 (RST), .A2 (nx7591), .B0 (nx1973), .B1 (nx2155)) ;
    inv01 ix2156 (.Y (nx2157), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_1)) ;
    oai32 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix413 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .A0 (
          nx2159), .A1 (RST), .A2 (nx7591), .B0 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx387), .B1 (nx2155)) ;
    inv01 ix2158 (.Y (nx2159), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_2)) ;
    oai32 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix423 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .A0 (
          nx2161), .A1 (RST), .A2 (nx7591), .B0 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx399), .B1 (nx2155)) ;
    inv01 ix2160 (.Y (nx2161), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_3)) ;
    oai32 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix433 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .A0 (
          nx2163), .A1 (RST), .A2 (nx7591), .B0 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx409), .B1 (nx2155)) ;
    inv01 ix2162 (.Y (nx2163), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_4)) ;
    oai32 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix443 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .A0 (
          nx2165), .A1 (RST), .A2 (nx7591), .B0 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx419), .B1 (nx2155)) ;
    inv01 ix2164 (.Y (nx2165), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_5)) ;
    oai32 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix453 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .A0 (
          nx2167), .A1 (RST), .A2 (nx7591), .B0 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx429), .B1 (nx2155)) ;
    inv01 ix2166 (.Y (nx2167), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_6)) ;
    oai32 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix463 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .A0 (
          nx2169), .A1 (RST), .A2 (nx7593), .B0 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx439), .B1 (nx2171)) ;
    inv01 ix2168 (.Y (nx2169), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_7)) ;
    oai32 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix473 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .A0 (
          nx2173), .A1 (RST), .A2 (nx7593), .B0 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx449), .B1 (nx2171)) ;
    inv01 ix2172 (.Y (nx2173), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_8)) ;
    oai32 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix483 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .A0 (
          nx2175), .A1 (RST), .A2 (nx7593), .B0 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx469), .B1 (nx2171)) ;
    inv01 ix2174 (.Y (nx2175), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_9)) ;
    oai32 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix493 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .A0 (
          nx2177), .A1 (RST), .A2 (nx7593), .B0 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx477), .B1 (nx2171)) ;
    inv01 ix2176 (.Y (nx2177), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_10)) ;
    oai32 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix503 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .A0 (
          nx2179), .A1 (RST), .A2 (nx7593), .B0 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx485), .B1 (nx2171)) ;
    inv01 ix2178 (.Y (nx2179), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_11)) ;
    oai32 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix513 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .A0 (
          nx2181), .A1 (RST), .A2 (nx7593), .B0 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx493), .B1 (nx2171)) ;
    inv01 ix2180 (.Y (nx2181), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_12)) ;
    oai32 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix523 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .A0 (
          nx2183), .A1 (RST), .A2 (nx7593), .B0 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx501), .B1 (nx2171)) ;
    inv01 ix2182 (.Y (nx2183), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_13)) ;
    oai32 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix533 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .A0 (
          nx2185), .A1 (RST), .A2 (nx7595), .B0 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx509), .B1 (nx2187)) ;
    inv01 ix2184 (.Y (nx2185), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_14)) ;
    inv01 ix2186 (.Y (nx2187), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566)) ;
    oai32 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix543 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .A0 (
          nx2189), .A1 (RST), .A2 (nx7595), .B0 (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_nx517), .B1 (nx2187)) ;
    inv01 ix2188 (.Y (nx2189), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_15)) ;
    oai32 CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix553 (.Y (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .A0 (
          nx2191), .A1 (RST), .A2 (nx7595), .B0 (nx1989), .B1 (nx2187)) ;
    inv01 ix2190 (.Y (nx2191), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_16)) ;
    nand02_2x CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix633 (.Y (
              nx2155), .A0 (nx7347), .A1 (nx7595)) ;
    nand02_2x CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix635 (.Y (
              nx2171), .A0 (nx7347), .A1 (nx7595)) ;
    mux21 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix404 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx403), .A0 (nx2193), .A1 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_2), .S0 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx395)) ;
    inv01 ix2192 (.Y (nx2193), .A (CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx391)) ;
    mux21 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix414 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx413), .A0 (nx2195), .A1 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_3), .S0 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx405)) ;
    inv01 ix2194 (.Y (nx2195), .A (CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx403)) ;
    mux21 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix424 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx423), .A0 (nx2197), .A1 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_4), .S0 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx415)) ;
    inv01 ix2196 (.Y (nx2197), .A (CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx413)) ;
    mux21 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix434 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx433), .A0 (nx2199), .A1 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_5), .S0 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx425)) ;
    inv01 ix2198 (.Y (nx2199), .A (CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx423)) ;
    mux21 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix444 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx443), .A0 (nx2201), .A1 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_6), .S0 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx435)) ;
    inv01 ix2200 (.Y (nx2201), .A (CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx433)) ;
    mux21 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix454 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx453), .A0 (nx2203), .A1 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_7), .S0 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx445)) ;
    inv01 ix2202 (.Y (nx2203), .A (CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx443)) ;
    mux21 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix462 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx461), .A0 (nx2205), .A1 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_8), .S0 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx455)) ;
    inv01 ix2204 (.Y (nx2205), .A (CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx453)) ;
    mux21 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix468 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx467), .A0 (nx2207), .A1 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_9), .S0 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx463)) ;
    inv01 ix2206 (.Y (nx2207), .A (CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx461)) ;
    mux21 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix476 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx475), .A0 (nx2209), .A1 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_10), .S0 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx471)) ;
    inv01 ix2208 (.Y (nx2209), .A (CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx467)) ;
    mux21 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix484 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx483), .A0 (nx2211), .A1 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_11), .S0 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx479)) ;
    inv01 ix2210 (.Y (nx2211), .A (CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx475)) ;
    mux21 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix492 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx491), .A0 (nx2213), .A1 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_12), .S0 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx487)) ;
    inv01 ix2212 (.Y (nx2213), .A (CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx483)) ;
    mux21 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix500 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx499), .A0 (nx2215), .A1 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_13), .S0 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx495)) ;
    inv01 ix2214 (.Y (nx2215), .A (CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx491)) ;
    mux21 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix508 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx507), .A0 (nx2217), .A1 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_14), .S0 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx503)) ;
    inv01 ix2216 (.Y (nx2217), .A (CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx499)) ;
    mux21 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix516 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx515), .A0 (nx2219), .A1 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_15), .S0 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx511)) ;
    inv01 ix2218 (.Y (nx2219), .A (CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx507)) ;
    mux21 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix161 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_1), .A0 (nx2221), .A1 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx379), .S0 (nx7599)) ;
    inv01 ix2220 (.Y (nx2221), .A (CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_1)) ;
    mux21 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix181 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_2), .A0 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx387), .A1 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx389), .S0 (nx7599)) ;
    mux21 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix201 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_3), .A0 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx399), .A1 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx401), .S0 (nx7599)) ;
    mux21 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix221 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_4), .A0 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx409), .A1 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx411), .S0 (nx7599)) ;
    mux21 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix241 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_5), .A0 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx419), .A1 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx421), .S0 (nx7599)) ;
    mux21 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix261 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_6), .A0 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx429), .A1 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx431), .S0 (nx7599)) ;
    mux21 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix281 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_7), .A0 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx439), .A1 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx441), .S0 (nx7599)) ;
    mux21 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix301 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_8), .A0 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx449), .A1 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx451), .S0 (nx7601)) ;
    mux21 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix321 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_9), .A0 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx469), .A1 (nx2223), .S0 (nx7601)) ;
    inv01 ix2222 (.Y (nx2223), .A (CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx316)) ;
    mux21 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix341 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_10), .A0 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx477), .A1 (nx2225), .S0 (nx7601)) ;
    inv01 ix2224 (.Y (nx2225), .A (CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx336)) ;
    mux21 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix361 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_11), .A0 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx485), .A1 (nx2227), .S0 (nx7601)) ;
    inv01 ix2226 (.Y (nx2227), .A (CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx356)) ;
    mux21 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix381 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_12), .A0 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx493), .A1 (nx2229), .S0 (nx7601)) ;
    inv01 ix2228 (.Y (nx2229), .A (CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx376)) ;
    mux21 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix401 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_13), .A0 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx501), .A1 (nx2231), .S0 (nx7601)) ;
    inv01 ix2230 (.Y (nx2231), .A (CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx396)) ;
    mux21 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix421 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_14), .A0 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx509), .A1 (nx2233), .S0 (nx7601)) ;
    inv01 ix2232 (.Y (nx2233), .A (CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx416)) ;
    mux21 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix441 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_15), .A0 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx517), .A1 (nx2235), .S0 (nx7603)) ;
    inv01 ix2234 (.Y (nx2235), .A (CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx436)) ;
    mux21 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_ix461 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_16), .A0 (nx2237), 
          .A1 (nx2239), .S0 (nx7603)) ;
    inv01 ix2236 (.Y (nx2237), .A (CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothP_16)
          ) ;
    inv01 ix2238 (.Y (nx2239), .A (CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx456)) ;
    nor02_2x CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix81 (.Y (
             CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx80), .A0 (Instr), .A1 (
             CALCULATOR_nx1111)) ;
    nor02_2x CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix319 (.Y (
             CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642), .A0 (
             CALCULATOR_Start_dup_1174), .A1 (
             CALCULATOR_CalculatingBooth_dup_1146)) ;
    nor02_2x CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix85 (.Y (
             CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_0), .A0 (
             nx7613), .A1 (nx2241)) ;
    inv01 ix2240 (.Y (nx2241), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_1)) ;
    mux21 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix125 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_1), .A0 (
          nx2243), .A1 (nx2245), .S0 (nx7613)) ;
    inv01 ix2242 (.Y (nx2243), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_2)) ;
    inv01 ix2244 (.Y (nx2245), .A (CacheWindow_1__1__0)) ;
    mux21 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix133 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_2), .A0 (
          nx2247), .A1 (nx2249), .S0 (nx7613)) ;
    inv01 ix2246 (.Y (nx2247), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_3)) ;
    inv01 ix2248 (.Y (nx2249), .A (CacheWindow_1__1__1)) ;
    mux21 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix141 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_3), .A0 (
          nx2251), .A1 (nx2253), .S0 (nx7613)) ;
    inv01 ix2250 (.Y (nx2251), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_4)) ;
    inv01 ix2252 (.Y (nx2253), .A (CacheWindow_1__1__2)) ;
    mux21 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix149 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_4), .A0 (
          nx2255), .A1 (nx2257), .S0 (nx7613)) ;
    inv01 ix2254 (.Y (nx2255), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_5)) ;
    inv01 ix2256 (.Y (nx2257), .A (CacheWindow_1__1__3)) ;
    mux21 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix157 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_5), .A0 (
          nx2259), .A1 (nx2261), .S0 (nx7613)) ;
    inv01 ix2258 (.Y (nx2259), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_6)) ;
    inv01 ix2260 (.Y (nx2261), .A (CacheWindow_1__1__4)) ;
    mux21 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix165 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_6), .A0 (
          nx2263), .A1 (nx2265), .S0 (nx7613)) ;
    inv01 ix2262 (.Y (nx2263), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_7)) ;
    inv01 ix2264 (.Y (nx2265), .A (CacheWindow_1__1__5)) ;
    mux21 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix173 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_7), .A0 (
          nx2267), .A1 (nx2269), .S0 (nx7615)) ;
    inv01 ix2266 (.Y (nx2267), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_8)) ;
    inv01 ix2268 (.Y (nx2269), .A (CacheWindow_1__1__6)) ;
    mux21 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix181 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_8), .A0 (
          nx2271), .A1 (nx2273), .S0 (nx7615)) ;
    inv01 ix2270 (.Y (nx2271), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_9)) ;
    inv01 ix2272 (.Y (nx2273), .A (CacheWindow_1__1__7)) ;
    nor02_2x CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix89 (.Y (
             CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_9), .A0 (
             nx7615), .A1 (nx2275)) ;
    inv01 ix2274 (.Y (nx2275), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_10)) ;
    nor02_2x CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix93 (.Y (
             CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_10), .A0 (
             nx7615), .A1 (nx2277)) ;
    inv01 ix2276 (.Y (nx2277), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_11)) ;
    nor02_2x CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix97 (.Y (
             CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_11), .A0 (
             nx7615), .A1 (nx2279)) ;
    inv01 ix2278 (.Y (nx2279), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_12)) ;
    nor02_2x CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix101 (.Y (
             CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_12), .A0 (
             nx7615), .A1 (nx2281)) ;
    inv01 ix2280 (.Y (nx2281), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_13)) ;
    nor02_2x CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix105 (.Y (
             CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_13), .A0 (
             nx7615), .A1 (nx2283)) ;
    inv01 ix2282 (.Y (nx2283), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_14)) ;
    nor02_2x CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix109 (.Y (
             CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_14), .A0 (
             nx7617), .A1 (nx2285)) ;
    inv01 ix2284 (.Y (nx2285), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_15)) ;
    nor02_2x CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix113 (.Y (
             CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_15), .A0 (
             nx7617), .A1 (nx2287)) ;
    inv01 ix2286 (.Y (nx2287), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_16)) ;
    nor02_2x CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix117 (.Y (
             CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_16), .A0 (
             nx7617), .A1 (nx2287)) ;
    mux21 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix189 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothOperand_0), .A0 (nx2289), .A1 (
          nx2291), .S0 (nx7605)) ;
    inv01 ix2288 (.Y (nx2289), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_0)) ;
    inv01 ix2290 (.Y (nx2291), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_0)) ;
    mux21 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix197 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothOperand_1), .A0 (nx2293), .A1 (
          nx2295), .S0 (nx7605)) ;
    inv01 ix2292 (.Y (nx2293), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_1)) ;
    inv01 ix2294 (.Y (nx2295), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_1)) ;
    mux21 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix205 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothOperand_2), .A0 (nx2297), .A1 (
          nx2299), .S0 (nx7605)) ;
    inv01 ix2296 (.Y (nx2297), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_2)) ;
    inv01 ix2298 (.Y (nx2299), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_2)) ;
    mux21 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix213 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothOperand_3), .A0 (nx2301), .A1 (
          nx2303), .S0 (nx7605)) ;
    inv01 ix2300 (.Y (nx2301), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_3)) ;
    inv01 ix2302 (.Y (nx2303), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_3)) ;
    mux21 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix221 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothOperand_4), .A0 (nx2305), .A1 (
          nx2307), .S0 (nx7605)) ;
    inv01 ix2304 (.Y (nx2305), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_4)) ;
    inv01 ix2306 (.Y (nx2307), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_4)) ;
    mux21 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix229 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothOperand_5), .A0 (nx2309), .A1 (
          nx2311), .S0 (nx7607)) ;
    inv01 ix2308 (.Y (nx2309), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_5)) ;
    inv01 ix2310 (.Y (nx2311), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_5)) ;
    mux21 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix237 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothOperand_6), .A0 (nx2313), .A1 (
          nx2315), .S0 (nx7607)) ;
    inv01 ix2312 (.Y (nx2313), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_6)) ;
    inv01 ix2314 (.Y (nx2315), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_6)) ;
    mux21 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix245 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothOperand_7), .A0 (nx2317), .A1 (
          nx2319), .S0 (nx7607)) ;
    inv01 ix2316 (.Y (nx2317), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_7)) ;
    inv01 ix2318 (.Y (nx2319), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_7)) ;
    mux21 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix253 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothOperand_8), .A0 (nx2321), .A1 (
          nx2323), .S0 (nx7607)) ;
    inv01 ix2320 (.Y (nx2321), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_8)) ;
    inv01 ix2322 (.Y (nx2323), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_8)) ;
    mux21 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix261 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothOperand_9), .A0 (nx2325), .A1 (
          nx2327), .S0 (nx7607)) ;
    inv01 ix2324 (.Y (nx2325), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_9)) ;
    inv01 ix2326 (.Y (nx2327), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_9)) ;
    mux21 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix269 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothOperand_10), .A0 (nx2329), .A1 (
          nx2331), .S0 (nx7607)) ;
    inv01 ix2328 (.Y (nx2329), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_10)) ;
    inv01 ix2330 (.Y (nx2331), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_10)) ;
    mux21 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix277 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothOperand_11), .A0 (nx2333), .A1 (
          nx2335), .S0 (nx7607)) ;
    inv01 ix2332 (.Y (nx2333), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_11)) ;
    inv01 ix2334 (.Y (nx2335), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_11)) ;
    mux21 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix285 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothOperand_12), .A0 (nx2337), .A1 (
          nx2339), .S0 (nx7609)) ;
    inv01 ix2336 (.Y (nx2337), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_12)) ;
    inv01 ix2338 (.Y (nx2339), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_12)) ;
    mux21 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix293 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothOperand_13), .A0 (nx2341), .A1 (
          nx2343), .S0 (nx7609)) ;
    inv01 ix2340 (.Y (nx2341), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_13)) ;
    inv01 ix2342 (.Y (nx2343), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_13)) ;
    mux21 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix301 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothOperand_14), .A0 (nx2345), .A1 (
          nx2347), .S0 (nx7609)) ;
    inv01 ix2344 (.Y (nx2345), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_14)) ;
    inv01 ix2346 (.Y (nx2347), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_14)) ;
    mux21 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix309 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothOperand_15), .A0 (nx2349), .A1 (
          nx2351), .S0 (nx7609)) ;
    inv01 ix2348 (.Y (nx2349), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_15)) ;
    inv01 ix2350 (.Y (nx2351), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_15)) ;
    mux21 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix317 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BoothOperand_16), .A0 (nx2353), .A1 (
          nx2355), .S0 (nx7609)) ;
    inv01 ix2352 (.Y (nx2353), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_16)) ;
    inv01 ix2354 (.Y (nx2355), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_16)) ;
    xnor2 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix321 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_AddPToBoothOperand), .A0 (nx7609), .A1 (
          nx2221)) ;
    oai32 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix393 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .A0 (
          nx8515), .A1 (RST), .A2 (nx7619), .B0 (nx2291), .B1 (nx2359)) ;
    oai32 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix403 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .A0 (
          nx8515), .A1 (RST), .A2 (nx7619), .B0 (nx2295), .B1 (nx2359)) ;
    oai32 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix413 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .A0 (
          nx8515), .A1 (RST), .A2 (nx7619), .B0 (nx2299), .B1 (nx2359)) ;
    oai32 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix423 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .A0 (
          nx8515), .A1 (RST), .A2 (nx7619), .B0 (nx2303), .B1 (nx2359)) ;
    oai32 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix433 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .A0 (
          nx8515), .A1 (RST), .A2 (nx7619), .B0 (nx2307), .B1 (nx2359)) ;
    oai32 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix443 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .A0 (
          nx8515), .A1 (RST), .A2 (nx7619), .B0 (nx2311), .B1 (nx2359)) ;
    oai32 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix453 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .A0 (
          nx8515), .A1 (RST), .A2 (nx7621), .B0 (nx2315), .B1 (nx2359)) ;
    oai32 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix463 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .A0 (
          nx8517), .A1 (RST), .A2 (nx7621), .B0 (nx2319), .B1 (nx2361)) ;
    oai32 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix473 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .A0 (
          nx8517), .A1 (RST), .A2 (nx7621), .B0 (nx2323), .B1 (nx2361)) ;
    oai32 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix483 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .A0 (
          nx2363), .A1 (RST), .A2 (nx7621), .B0 (nx2327), .B1 (nx2361)) ;
    inv01 ix2362 (.Y (nx2363), .A (CacheFilter_1__1__0)) ;
    oai32 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix493 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .A0 (
          nx2365), .A1 (RST), .A2 (nx7621), .B0 (nx2331), .B1 (nx2361)) ;
    inv01 ix2364 (.Y (nx2365), .A (CacheFilter_1__1__1)) ;
    oai32 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix503 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .A0 (
          nx2367), .A1 (RST), .A2 (nx7621), .B0 (nx2335), .B1 (nx2361)) ;
    inv01 ix2366 (.Y (nx2367), .A (CacheFilter_1__1__2)) ;
    oai32 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix513 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .A0 (
          nx2369), .A1 (RST), .A2 (nx7621), .B0 (nx2339), .B1 (nx2361)) ;
    inv01 ix2368 (.Y (nx2369), .A (CacheFilter_1__1__3)) ;
    oai32 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix523 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .A0 (
          nx2371), .A1 (RST), .A2 (nx7623), .B0 (nx2343), .B1 (nx2361)) ;
    inv01 ix2370 (.Y (nx2371), .A (CacheFilter_1__1__4)) ;
    oai32 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix533 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .A0 (
          nx2373), .A1 (RST), .A2 (nx7623), .B0 (nx2347), .B1 (nx2375)) ;
    inv01 ix2372 (.Y (nx2373), .A (CacheFilter_1__1__5)) ;
    inv01 ix2374 (.Y (nx2375), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566)) ;
    oai32 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix543 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .A0 (
          nx2377), .A1 (RST), .A2 (nx7623), .B0 (nx2351), .B1 (nx2375)) ;
    inv01 ix2376 (.Y (nx2377), .A (CacheFilter_1__1__6)) ;
    oai32 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix553 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .A0 (
          nx2379), .A1 (RST), .A2 (nx7623), .B0 (nx2355), .B1 (nx2375)) ;
    inv01 ix2378 (.Y (nx2379), .A (CacheFilter_1__1__7)) ;
    nand02_2x CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix633 (.Y (
              nx2359), .A0 (nx7347), .A1 (nx7623)) ;
    nand02_2x CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix635 (.Y (
              nx2361), .A0 (nx7347), .A1 (nx7623)) ;
    oai32 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix393 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .A0 (
          nx8517), .A1 (RST), .A2 (nx7625), .B0 (nx2289), .B1 (nx2381)) ;
    oai32 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix403 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .A0 (
          nx8517), .A1 (RST), .A2 (nx7625), .B0 (nx2293), .B1 (nx2381)) ;
    oai32 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix413 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .A0 (
          nx8517), .A1 (RST), .A2 (nx7625), .B0 (nx2297), .B1 (nx2381)) ;
    oai32 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix423 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .A0 (
          nx8517), .A1 (RST), .A2 (nx7625), .B0 (nx2301), .B1 (nx2381)) ;
    oai32 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix433 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .A0 (
          nx8517), .A1 (RST), .A2 (nx7625), .B0 (nx2305), .B1 (nx2381)) ;
    oai32 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix443 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .A0 (
          nx8519), .A1 (RST), .A2 (nx7625), .B0 (nx2309), .B1 (nx2381)) ;
    oai32 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix453 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .A0 (
          nx8519), .A1 (RST), .A2 (nx7627), .B0 (nx2313), .B1 (nx2381)) ;
    oai32 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix463 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .A0 (
          nx8519), .A1 (RST), .A2 (nx7627), .B0 (nx2317), .B1 (nx2383)) ;
    oai32 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix473 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .A0 (
          nx8519), .A1 (RST), .A2 (nx7627), .B0 (nx2321), .B1 (nx2383)) ;
    oai32 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix483 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .A0 (
          nx2363), .A1 (RST), .A2 (nx7627), .B0 (nx2325), .B1 (nx2383)) ;
    oai32 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix493 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .A0 (
          nx2385), .A1 (RST), .A2 (nx7627), .B0 (nx2329), .B1 (nx2383)) ;
    inv01 ix2384 (.Y (nx2385), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_10)) ;
    oai32 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix503 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .A0 (
          nx2387), .A1 (RST), .A2 (nx7627), .B0 (nx2333), .B1 (nx2383)) ;
    inv01 ix2386 (.Y (nx2387), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_11)) ;
    oai32 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix513 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .A0 (
          nx2389), .A1 (RST), .A2 (nx7627), .B0 (nx2337), .B1 (nx2383)) ;
    inv01 ix2388 (.Y (nx2389), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_12)) ;
    oai32 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix523 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .A0 (
          nx2391), .A1 (RST), .A2 (nx7629), .B0 (nx2341), .B1 (nx2383)) ;
    inv01 ix2390 (.Y (nx2391), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_13)) ;
    oai32 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix533 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .A0 (
          nx2393), .A1 (RST), .A2 (nx7629), .B0 (nx2345), .B1 (nx2395)) ;
    inv01 ix2392 (.Y (nx2393), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_14)) ;
    inv01 ix2394 (.Y (nx2395), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566)) ;
    oai32 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix543 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .A0 (
          nx2397), .A1 (RST), .A2 (nx7629), .B0 (nx2349), .B1 (nx2395)) ;
    inv01 ix2396 (.Y (nx2397), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_15)) ;
    oai32 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix553 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .A0 (
          nx2399), .A1 (RST), .A2 (nx7629), .B0 (nx2353), .B1 (nx2395)) ;
    inv01 ix2398 (.Y (nx2399), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_16)) ;
    nand02_2x CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix633 (.Y (
              nx2381), .A0 (nx7347), .A1 (nx7629)) ;
    nand02_2x CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix635 (.Y (
              nx2383), .A0 (nx7347), .A1 (nx7629)) ;
    oai32 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix393 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .A0 (
          nx2401), .A1 (RST), .A2 (nx7631), .B0 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx384), .B1 (nx2403)) ;
    inv01 ix2400 (.Y (nx2401), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_0)) ;
    oai32 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix403 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .A0 (
          nx2405), .A1 (RST), .A2 (nx7631), .B0 (nx2221), .B1 (nx2403)) ;
    inv01 ix2404 (.Y (nx2405), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_1)) ;
    oai32 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix413 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .A0 (
          nx2407), .A1 (RST), .A2 (nx7631), .B0 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx387), .B1 (nx2403)) ;
    inv01 ix2406 (.Y (nx2407), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_2)) ;
    oai32 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix423 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .A0 (
          nx2409), .A1 (RST), .A2 (nx7631), .B0 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx399), .B1 (nx2403)) ;
    inv01 ix2408 (.Y (nx2409), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_3)) ;
    oai32 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix433 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .A0 (
          nx2411), .A1 (RST), .A2 (nx7631), .B0 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx409), .B1 (nx2403)) ;
    inv01 ix2410 (.Y (nx2411), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_4)) ;
    oai32 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix443 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .A0 (
          nx2413), .A1 (RST), .A2 (nx7631), .B0 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx419), .B1 (nx2403)) ;
    inv01 ix2412 (.Y (nx2413), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_5)) ;
    oai32 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix453 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .A0 (
          nx2415), .A1 (RST), .A2 (nx7631), .B0 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx429), .B1 (nx2403)) ;
    inv01 ix2414 (.Y (nx2415), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_6)) ;
    oai32 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix463 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .A0 (
          nx2417), .A1 (RST), .A2 (nx7633), .B0 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx439), .B1 (nx2419)) ;
    inv01 ix2416 (.Y (nx2417), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_7)) ;
    oai32 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix473 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .A0 (
          nx2421), .A1 (RST), .A2 (nx7633), .B0 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx449), .B1 (nx2419)) ;
    inv01 ix2420 (.Y (nx2421), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_8)) ;
    oai32 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix483 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .A0 (
          nx2423), .A1 (RST), .A2 (nx7633), .B0 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx469), .B1 (nx2419)) ;
    inv01 ix2422 (.Y (nx2423), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_9)) ;
    oai32 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix493 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .A0 (
          nx2425), .A1 (RST), .A2 (nx7633), .B0 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx477), .B1 (nx2419)) ;
    inv01 ix2424 (.Y (nx2425), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_10)) ;
    oai32 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix503 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .A0 (
          nx2427), .A1 (RST), .A2 (nx7633), .B0 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx485), .B1 (nx2419)) ;
    inv01 ix2426 (.Y (nx2427), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_11)) ;
    oai32 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix513 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .A0 (
          nx2429), .A1 (RST), .A2 (nx7633), .B0 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx493), .B1 (nx2419)) ;
    inv01 ix2428 (.Y (nx2429), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_12)) ;
    oai32 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix523 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .A0 (
          nx2431), .A1 (RST), .A2 (nx7633), .B0 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx501), .B1 (nx2419)) ;
    inv01 ix2430 (.Y (nx2431), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_13)) ;
    oai32 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix533 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .A0 (
          nx2433), .A1 (RST), .A2 (nx7635), .B0 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx509), .B1 (nx2435)) ;
    inv01 ix2432 (.Y (nx2433), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_14)) ;
    inv01 ix2434 (.Y (nx2435), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566)) ;
    oai32 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix543 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .A0 (
          nx2437), .A1 (RST), .A2 (nx7635), .B0 (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_nx517), .B1 (nx2435)) ;
    inv01 ix2436 (.Y (nx2437), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_15)) ;
    oai32 CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix553 (.Y (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .A0 (
          nx2439), .A1 (RST), .A2 (nx7635), .B0 (nx2237), .B1 (nx2435)) ;
    inv01 ix2438 (.Y (nx2439), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_16)) ;
    nand02_2x CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix633 (.Y (
              nx2403), .A0 (nx7347), .A1 (nx7635)) ;
    nand02_2x CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix635 (.Y (
              nx2419), .A0 (nx7349), .A1 (nx7635)) ;
    mux21 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix404 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx403), .A0 (nx2441), .A1 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_2), .S0 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx395)) ;
    inv01 ix2440 (.Y (nx2441), .A (CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx391)) ;
    mux21 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix414 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx413), .A0 (nx2443), .A1 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_3), .S0 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx405)) ;
    inv01 ix2442 (.Y (nx2443), .A (CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx403)) ;
    mux21 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix424 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx423), .A0 (nx2445), .A1 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_4), .S0 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx415)) ;
    inv01 ix2444 (.Y (nx2445), .A (CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx413)) ;
    mux21 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix434 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx433), .A0 (nx2447), .A1 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_5), .S0 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx425)) ;
    inv01 ix2446 (.Y (nx2447), .A (CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx423)) ;
    mux21 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix444 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx443), .A0 (nx2449), .A1 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_6), .S0 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx435)) ;
    inv01 ix2448 (.Y (nx2449), .A (CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx433)) ;
    mux21 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix454 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx453), .A0 (nx2451), .A1 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_7), .S0 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx445)) ;
    inv01 ix2450 (.Y (nx2451), .A (CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx443)) ;
    mux21 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix462 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx461), .A0 (nx2453), .A1 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_8), .S0 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx455)) ;
    inv01 ix2452 (.Y (nx2453), .A (CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx453)) ;
    mux21 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix468 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx467), .A0 (nx2455), .A1 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_9), .S0 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx463)) ;
    inv01 ix2454 (.Y (nx2455), .A (CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx461)) ;
    mux21 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix476 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx475), .A0 (nx2457), .A1 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_10), .S0 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx471)) ;
    inv01 ix2456 (.Y (nx2457), .A (CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx467)) ;
    mux21 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix484 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx483), .A0 (nx2459), .A1 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_11), .S0 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx479)) ;
    inv01 ix2458 (.Y (nx2459), .A (CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx475)) ;
    mux21 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix492 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx491), .A0 (nx2461), .A1 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_12), .S0 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx487)) ;
    inv01 ix2460 (.Y (nx2461), .A (CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx483)) ;
    mux21 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix500 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx499), .A0 (nx2463), .A1 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_13), .S0 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx495)) ;
    inv01 ix2462 (.Y (nx2463), .A (CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx491)) ;
    mux21 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix508 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx507), .A0 (nx2465), .A1 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_14), .S0 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx503)) ;
    inv01 ix2464 (.Y (nx2465), .A (CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx499)) ;
    mux21 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix516 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx515), .A0 (nx2467), .A1 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_15), .S0 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx511)) ;
    inv01 ix2466 (.Y (nx2467), .A (CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx507)) ;
    mux21 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix161 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_1), .A0 (nx2469), .A1 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx379), .S0 (nx7639)) ;
    inv01 ix2468 (.Y (nx2469), .A (CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_1)) ;
    mux21 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix181 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_2), .A0 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx387), .A1 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx389), .S0 (nx7639)) ;
    mux21 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix201 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_3), .A0 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx399), .A1 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx401), .S0 (nx7639)) ;
    mux21 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix221 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_4), .A0 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx409), .A1 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx411), .S0 (nx7639)) ;
    mux21 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix241 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_5), .A0 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx419), .A1 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx421), .S0 (nx7639)) ;
    mux21 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix261 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_6), .A0 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx429), .A1 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx431), .S0 (nx7639)) ;
    mux21 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix281 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_7), .A0 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx439), .A1 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx441), .S0 (nx7639)) ;
    mux21 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix301 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_8), .A0 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx449), .A1 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx451), .S0 (nx7641)) ;
    mux21 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix321 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_9), .A0 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx469), .A1 (nx2471), .S0 (nx7641)) ;
    inv01 ix2470 (.Y (nx2471), .A (CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx316)) ;
    mux21 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix341 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_10), .A0 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx477), .A1 (nx2473), .S0 (nx7641)) ;
    inv01 ix2472 (.Y (nx2473), .A (CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx336)) ;
    mux21 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix361 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_11), .A0 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx485), .A1 (nx2475), .S0 (nx7641)) ;
    inv01 ix2474 (.Y (nx2475), .A (CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx356)) ;
    mux21 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix381 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_12), .A0 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx493), .A1 (nx2477), .S0 (nx7641)) ;
    inv01 ix2476 (.Y (nx2477), .A (CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx376)) ;
    mux21 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix401 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_13), .A0 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx501), .A1 (nx2479), .S0 (nx7641)) ;
    inv01 ix2478 (.Y (nx2479), .A (CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx396)) ;
    mux21 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix421 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_14), .A0 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx509), .A1 (nx2481), .S0 (nx7641)) ;
    inv01 ix2480 (.Y (nx2481), .A (CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx416)) ;
    mux21 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix441 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_15), .A0 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx517), .A1 (nx2483), .S0 (nx7643)) ;
    inv01 ix2482 (.Y (nx2483), .A (CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx436)) ;
    mux21 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_ix461 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_16), .A0 (nx2485), 
          .A1 (nx2487), .S0 (nx7643)) ;
    inv01 ix2484 (.Y (nx2485), .A (CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothP_16)
          ) ;
    inv01 ix2486 (.Y (nx2487), .A (CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx456)) ;
    nor02_2x CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix81 (.Y (
             CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx80), .A0 (Instr), .A1 (
             nx7309)) ;
    nor02_2x CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix319 (.Y (
             CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642), .A0 (
             CALCULATOR_Start_dup_1179), .A1 (
             CALCULATOR_CalculatingBooth_dup_1181)) ;
    nor02_2x CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix85 (.Y (
             CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_0), .A0 (
             nx7653), .A1 (nx2489)) ;
    inv01 ix2488 (.Y (nx2489), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_1)) ;
    mux21 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix125 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_1), .A0 (
          nx2491), .A1 (nx2493), .S0 (nx7653)) ;
    inv01 ix2490 (.Y (nx2491), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_2)) ;
    inv01 ix2492 (.Y (nx2493), .A (CacheWindow_1__2__0)) ;
    mux21 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix133 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_2), .A0 (
          nx2495), .A1 (nx2497), .S0 (nx7653)) ;
    inv01 ix2494 (.Y (nx2495), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_3)) ;
    inv01 ix2496 (.Y (nx2497), .A (CacheWindow_1__2__1)) ;
    mux21 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix141 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_3), .A0 (
          nx2499), .A1 (nx2501), .S0 (nx7653)) ;
    inv01 ix2498 (.Y (nx2499), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_4)) ;
    inv01 ix2500 (.Y (nx2501), .A (CacheWindow_1__2__2)) ;
    mux21 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix149 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_4), .A0 (
          nx2503), .A1 (nx2505), .S0 (nx7653)) ;
    inv01 ix2502 (.Y (nx2503), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_5)) ;
    inv01 ix2504 (.Y (nx2505), .A (CacheWindow_1__2__3)) ;
    mux21 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix157 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_5), .A0 (
          nx2507), .A1 (nx2509), .S0 (nx7653)) ;
    inv01 ix2506 (.Y (nx2507), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_6)) ;
    inv01 ix2508 (.Y (nx2509), .A (CacheWindow_1__2__4)) ;
    mux21 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix165 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_6), .A0 (
          nx2511), .A1 (nx2513), .S0 (nx7653)) ;
    inv01 ix2510 (.Y (nx2511), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_7)) ;
    inv01 ix2512 (.Y (nx2513), .A (CacheWindow_1__2__5)) ;
    mux21 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix173 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_7), .A0 (
          nx2515), .A1 (nx2517), .S0 (nx7655)) ;
    inv01 ix2514 (.Y (nx2515), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_8)) ;
    inv01 ix2516 (.Y (nx2517), .A (CacheWindow_1__2__6)) ;
    mux21 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix181 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_8), .A0 (
          nx2519), .A1 (nx2521), .S0 (nx7655)) ;
    inv01 ix2518 (.Y (nx2519), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_9)) ;
    inv01 ix2520 (.Y (nx2521), .A (CacheWindow_1__2__7)) ;
    nor02_2x CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix89 (.Y (
             CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_9), .A0 (
             nx7655), .A1 (nx2523)) ;
    inv01 ix2522 (.Y (nx2523), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_10)) ;
    nor02_2x CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix93 (.Y (
             CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_10), .A0 (
             nx7655), .A1 (nx2525)) ;
    inv01 ix2524 (.Y (nx2525), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_11)) ;
    nor02_2x CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix97 (.Y (
             CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_11), .A0 (
             nx7655), .A1 (nx2527)) ;
    inv01 ix2526 (.Y (nx2527), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_12)) ;
    nor02_2x CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix101 (.Y (
             CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_12), .A0 (
             nx7655), .A1 (nx2529)) ;
    inv01 ix2528 (.Y (nx2529), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_13)) ;
    nor02_2x CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix105 (.Y (
             CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_13), .A0 (
             nx7655), .A1 (nx2531)) ;
    inv01 ix2530 (.Y (nx2531), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_14)) ;
    nor02_2x CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix109 (.Y (
             CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_14), .A0 (
             nx7657), .A1 (nx2533)) ;
    inv01 ix2532 (.Y (nx2533), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_15)) ;
    nor02_2x CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix113 (.Y (
             CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_15), .A0 (
             nx7657), .A1 (nx2535)) ;
    inv01 ix2534 (.Y (nx2535), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_16)) ;
    nor02_2x CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix117 (.Y (
             CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_16), .A0 (
             nx7657), .A1 (nx2535)) ;
    mux21 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix189 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothOperand_0), .A0 (nx2537), .A1 (
          nx2539), .S0 (nx7645)) ;
    inv01 ix2536 (.Y (nx2537), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_0)) ;
    inv01 ix2538 (.Y (nx2539), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_0)) ;
    mux21 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix197 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothOperand_1), .A0 (nx2541), .A1 (
          nx2543), .S0 (nx7645)) ;
    inv01 ix2540 (.Y (nx2541), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_1)) ;
    inv01 ix2542 (.Y (nx2543), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_1)) ;
    mux21 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix205 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothOperand_2), .A0 (nx2545), .A1 (
          nx2547), .S0 (nx7645)) ;
    inv01 ix2544 (.Y (nx2545), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_2)) ;
    inv01 ix2546 (.Y (nx2547), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_2)) ;
    mux21 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix213 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothOperand_3), .A0 (nx2549), .A1 (
          nx2551), .S0 (nx7645)) ;
    inv01 ix2548 (.Y (nx2549), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_3)) ;
    inv01 ix2550 (.Y (nx2551), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_3)) ;
    mux21 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix221 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothOperand_4), .A0 (nx2553), .A1 (
          nx2555), .S0 (nx7645)) ;
    inv01 ix2552 (.Y (nx2553), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_4)) ;
    inv01 ix2554 (.Y (nx2555), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_4)) ;
    mux21 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix229 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothOperand_5), .A0 (nx2557), .A1 (
          nx2559), .S0 (nx7647)) ;
    inv01 ix2556 (.Y (nx2557), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_5)) ;
    inv01 ix2558 (.Y (nx2559), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_5)) ;
    mux21 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix237 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothOperand_6), .A0 (nx2561), .A1 (
          nx2563), .S0 (nx7647)) ;
    inv01 ix2560 (.Y (nx2561), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_6)) ;
    inv01 ix2562 (.Y (nx2563), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_6)) ;
    mux21 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix245 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothOperand_7), .A0 (nx2565), .A1 (
          nx2567), .S0 (nx7647)) ;
    inv01 ix2564 (.Y (nx2565), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_7)) ;
    inv01 ix2566 (.Y (nx2567), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_7)) ;
    mux21 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix253 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothOperand_8), .A0 (nx2569), .A1 (
          nx2571), .S0 (nx7647)) ;
    inv01 ix2568 (.Y (nx2569), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_8)) ;
    inv01 ix2570 (.Y (nx2571), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_8)) ;
    mux21 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix261 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothOperand_9), .A0 (nx2573), .A1 (
          nx2575), .S0 (nx7647)) ;
    inv01 ix2572 (.Y (nx2573), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_9)) ;
    inv01 ix2574 (.Y (nx2575), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_9)) ;
    mux21 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix269 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothOperand_10), .A0 (nx2577), .A1 (
          nx2579), .S0 (nx7647)) ;
    inv01 ix2576 (.Y (nx2577), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_10)) ;
    inv01 ix2578 (.Y (nx2579), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_10)) ;
    mux21 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix277 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothOperand_11), .A0 (nx2581), .A1 (
          nx2583), .S0 (nx7647)) ;
    inv01 ix2580 (.Y (nx2581), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_11)) ;
    inv01 ix2582 (.Y (nx2583), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_11)) ;
    mux21 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix285 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothOperand_12), .A0 (nx2585), .A1 (
          nx2587), .S0 (nx7649)) ;
    inv01 ix2584 (.Y (nx2585), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_12)) ;
    inv01 ix2586 (.Y (nx2587), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_12)) ;
    mux21 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix293 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothOperand_13), .A0 (nx2589), .A1 (
          nx2591), .S0 (nx7649)) ;
    inv01 ix2588 (.Y (nx2589), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_13)) ;
    inv01 ix2590 (.Y (nx2591), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_13)) ;
    mux21 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix301 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothOperand_14), .A0 (nx2593), .A1 (
          nx2595), .S0 (nx7649)) ;
    inv01 ix2592 (.Y (nx2593), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_14)) ;
    inv01 ix2594 (.Y (nx2595), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_14)) ;
    mux21 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix309 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothOperand_15), .A0 (nx2597), .A1 (
          nx2599), .S0 (nx7649)) ;
    inv01 ix2596 (.Y (nx2597), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_15)) ;
    inv01 ix2598 (.Y (nx2599), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_15)) ;
    mux21 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix317 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BoothOperand_16), .A0 (nx2601), .A1 (
          nx2603), .S0 (nx7649)) ;
    inv01 ix2600 (.Y (nx2601), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_16)) ;
    inv01 ix2602 (.Y (nx2603), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_16)) ;
    xnor2 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix321 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_AddPToBoothOperand), .A0 (nx7649), .A1 (
          nx2469)) ;
    oai32 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix393 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .A0 (
          nx8521), .A1 (RST), .A2 (nx7659), .B0 (nx2539), .B1 (nx2607)) ;
    oai32 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix403 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .A0 (
          nx8521), .A1 (RST), .A2 (nx7659), .B0 (nx2543), .B1 (nx2607)) ;
    oai32 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix413 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .A0 (
          nx8521), .A1 (RST), .A2 (nx7659), .B0 (nx2547), .B1 (nx2607)) ;
    oai32 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix423 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .A0 (
          nx8521), .A1 (RST), .A2 (nx7659), .B0 (nx2551), .B1 (nx2607)) ;
    oai32 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix433 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .A0 (
          nx8521), .A1 (RST), .A2 (nx7659), .B0 (nx2555), .B1 (nx2607)) ;
    oai32 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix443 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .A0 (
          nx8521), .A1 (RST), .A2 (nx7659), .B0 (nx2559), .B1 (nx2607)) ;
    oai32 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix453 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .A0 (
          nx8521), .A1 (RST), .A2 (nx7661), .B0 (nx2563), .B1 (nx2607)) ;
    oai32 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix463 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .A0 (
          nx8523), .A1 (RST), .A2 (nx7661), .B0 (nx2567), .B1 (nx2609)) ;
    oai32 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix473 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .A0 (
          nx8523), .A1 (RST), .A2 (nx7661), .B0 (nx2571), .B1 (nx2609)) ;
    oai32 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix483 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .A0 (
          nx2611), .A1 (RST), .A2 (nx7661), .B0 (nx2575), .B1 (nx2609)) ;
    inv01 ix2610 (.Y (nx2611), .A (CacheFilter_1__2__0)) ;
    oai32 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix493 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .A0 (
          nx2613), .A1 (RST), .A2 (nx7661), .B0 (nx2579), .B1 (nx2609)) ;
    inv01 ix2612 (.Y (nx2613), .A (CacheFilter_1__2__1)) ;
    oai32 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix503 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .A0 (
          nx2615), .A1 (RST), .A2 (nx7661), .B0 (nx2583), .B1 (nx2609)) ;
    inv01 ix2614 (.Y (nx2615), .A (CacheFilter_1__2__2)) ;
    oai32 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix513 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .A0 (
          nx2617), .A1 (RST), .A2 (nx7661), .B0 (nx2587), .B1 (nx2609)) ;
    inv01 ix2616 (.Y (nx2617), .A (CacheFilter_1__2__3)) ;
    oai32 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix523 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .A0 (
          nx2619), .A1 (RST), .A2 (nx7663), .B0 (nx2591), .B1 (nx2609)) ;
    inv01 ix2618 (.Y (nx2619), .A (CacheFilter_1__2__4)) ;
    oai32 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix533 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .A0 (
          nx2621), .A1 (RST), .A2 (nx7663), .B0 (nx2595), .B1 (nx2623)) ;
    inv01 ix2620 (.Y (nx2621), .A (CacheFilter_1__2__5)) ;
    inv01 ix2622 (.Y (nx2623), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566)) ;
    oai32 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix543 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .A0 (
          nx2625), .A1 (RST), .A2 (nx7663), .B0 (nx2599), .B1 (nx2623)) ;
    inv01 ix2624 (.Y (nx2625), .A (CacheFilter_1__2__6)) ;
    oai32 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix553 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .A0 (
          nx2627), .A1 (RST), .A2 (nx7663), .B0 (nx2603), .B1 (nx2623)) ;
    inv01 ix2626 (.Y (nx2627), .A (CacheFilter_1__2__7)) ;
    nand02_2x CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix633 (.Y (
              nx2607), .A0 (nx7349), .A1 (nx7663)) ;
    nand02_2x CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix635 (.Y (
              nx2609), .A0 (nx7349), .A1 (nx7663)) ;
    oai32 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix393 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .A0 (
          nx8523), .A1 (RST), .A2 (nx7665), .B0 (nx2537), .B1 (nx2629)) ;
    oai32 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix403 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .A0 (
          nx8523), .A1 (RST), .A2 (nx7665), .B0 (nx2541), .B1 (nx2629)) ;
    oai32 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix413 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .A0 (
          nx8523), .A1 (RST), .A2 (nx7665), .B0 (nx2545), .B1 (nx2629)) ;
    oai32 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix423 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .A0 (
          nx8523), .A1 (RST), .A2 (nx7665), .B0 (nx2549), .B1 (nx2629)) ;
    oai32 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix433 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .A0 (
          nx8523), .A1 (RST), .A2 (nx7665), .B0 (nx2553), .B1 (nx2629)) ;
    oai32 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix443 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .A0 (
          nx8525), .A1 (RST), .A2 (nx7665), .B0 (nx2557), .B1 (nx2629)) ;
    oai32 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix453 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .A0 (
          nx8525), .A1 (RST), .A2 (nx7667), .B0 (nx2561), .B1 (nx2629)) ;
    oai32 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix463 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .A0 (
          nx8525), .A1 (RST), .A2 (nx7667), .B0 (nx2565), .B1 (nx2631)) ;
    oai32 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix473 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .A0 (
          nx8525), .A1 (RST), .A2 (nx7667), .B0 (nx2569), .B1 (nx2631)) ;
    oai32 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix483 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .A0 (
          nx2611), .A1 (RST), .A2 (nx7667), .B0 (nx2573), .B1 (nx2631)) ;
    oai32 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix493 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .A0 (
          nx2633), .A1 (RST), .A2 (nx7667), .B0 (nx2577), .B1 (nx2631)) ;
    inv01 ix2632 (.Y (nx2633), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_10)) ;
    oai32 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix503 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .A0 (
          nx2635), .A1 (RST), .A2 (nx7667), .B0 (nx2581), .B1 (nx2631)) ;
    inv01 ix2634 (.Y (nx2635), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_11)) ;
    oai32 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix513 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .A0 (
          nx2637), .A1 (RST), .A2 (nx7667), .B0 (nx2585), .B1 (nx2631)) ;
    inv01 ix2636 (.Y (nx2637), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_12)) ;
    oai32 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix523 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .A0 (
          nx2639), .A1 (RST), .A2 (nx7669), .B0 (nx2589), .B1 (nx2631)) ;
    inv01 ix2638 (.Y (nx2639), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_13)) ;
    oai32 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix533 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .A0 (
          nx2641), .A1 (RST), .A2 (nx7669), .B0 (nx2593), .B1 (nx2643)) ;
    inv01 ix2640 (.Y (nx2641), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_14)) ;
    inv01 ix2642 (.Y (nx2643), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566)) ;
    oai32 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix543 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .A0 (
          nx2645), .A1 (RST), .A2 (nx7669), .B0 (nx2597), .B1 (nx2643)) ;
    inv01 ix2644 (.Y (nx2645), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_15)) ;
    oai32 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix553 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .A0 (
          nx2647), .A1 (RST), .A2 (nx7669), .B0 (nx2601), .B1 (nx2643)) ;
    inv01 ix2646 (.Y (nx2647), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_16)) ;
    nand02_2x CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix633 (.Y (
              nx2629), .A0 (nx7349), .A1 (nx7669)) ;
    nand02_2x CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix635 (.Y (
              nx2631), .A0 (nx7349), .A1 (nx7669)) ;
    oai32 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix393 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .A0 (
          nx2649), .A1 (RST), .A2 (nx7671), .B0 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx384), .B1 (nx2651)) ;
    inv01 ix2648 (.Y (nx2649), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_0)) ;
    oai32 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix403 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .A0 (
          nx2653), .A1 (RST), .A2 (nx7671), .B0 (nx2469), .B1 (nx2651)) ;
    inv01 ix2652 (.Y (nx2653), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_1)) ;
    oai32 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix413 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .A0 (
          nx2655), .A1 (RST), .A2 (nx7671), .B0 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx387), .B1 (nx2651)) ;
    inv01 ix2654 (.Y (nx2655), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_2)) ;
    oai32 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix423 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .A0 (
          nx2657), .A1 (RST), .A2 (nx7671), .B0 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx399), .B1 (nx2651)) ;
    inv01 ix2656 (.Y (nx2657), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_3)) ;
    oai32 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix433 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .A0 (
          nx2659), .A1 (RST), .A2 (nx7671), .B0 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx409), .B1 (nx2651)) ;
    inv01 ix2658 (.Y (nx2659), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_4)) ;
    oai32 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix443 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .A0 (
          nx2661), .A1 (RST), .A2 (nx7671), .B0 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx419), .B1 (nx2651)) ;
    inv01 ix2660 (.Y (nx2661), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_5)) ;
    oai32 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix453 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .A0 (
          nx2663), .A1 (RST), .A2 (nx7671), .B0 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx429), .B1 (nx2651)) ;
    inv01 ix2662 (.Y (nx2663), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_6)) ;
    oai32 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix463 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .A0 (
          nx2665), .A1 (RST), .A2 (nx7673), .B0 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx439), .B1 (nx2667)) ;
    inv01 ix2664 (.Y (nx2665), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_7)) ;
    oai32 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix473 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .A0 (
          nx2669), .A1 (RST), .A2 (nx7673), .B0 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx449), .B1 (nx2667)) ;
    inv01 ix2668 (.Y (nx2669), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_8)) ;
    oai32 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix483 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .A0 (
          nx2671), .A1 (RST), .A2 (nx7673), .B0 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx469), .B1 (nx2667)) ;
    inv01 ix2670 (.Y (nx2671), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_9)) ;
    oai32 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix493 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .A0 (
          nx2673), .A1 (RST), .A2 (nx7673), .B0 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx477), .B1 (nx2667)) ;
    inv01 ix2672 (.Y (nx2673), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_10)) ;
    oai32 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix503 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .A0 (
          nx2675), .A1 (RST), .A2 (nx7673), .B0 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx485), .B1 (nx2667)) ;
    inv01 ix2674 (.Y (nx2675), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_11)) ;
    oai32 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix513 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .A0 (
          nx2677), .A1 (RST), .A2 (nx7673), .B0 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx493), .B1 (nx2667)) ;
    inv01 ix2676 (.Y (nx2677), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_12)) ;
    oai32 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix523 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .A0 (
          nx2679), .A1 (RST), .A2 (nx7673), .B0 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx501), .B1 (nx2667)) ;
    inv01 ix2678 (.Y (nx2679), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_13)) ;
    oai32 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix533 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .A0 (
          nx2681), .A1 (RST), .A2 (nx7675), .B0 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx509), .B1 (nx2683)) ;
    inv01 ix2680 (.Y (nx2681), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_14)) ;
    inv01 ix2682 (.Y (nx2683), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566)) ;
    oai32 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix543 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .A0 (
          nx2685), .A1 (RST), .A2 (nx7675), .B0 (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_nx517), .B1 (nx2683)) ;
    inv01 ix2684 (.Y (nx2685), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_15)) ;
    oai32 CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix553 (.Y (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .A0 (
          nx2687), .A1 (RST), .A2 (nx7675), .B0 (nx2485), .B1 (nx2683)) ;
    inv01 ix2686 (.Y (nx2687), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_16)) ;
    nand02_2x CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix633 (.Y (
              nx2651), .A0 (nx7349), .A1 (nx7675)) ;
    nand02_2x CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix635 (.Y (
              nx2667), .A0 (nx7349), .A1 (nx7675)) ;
    mux21 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix404 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx403), .A0 (nx2689), .A1 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_2), .S0 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx395)) ;
    inv01 ix2688 (.Y (nx2689), .A (CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx391)) ;
    mux21 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix414 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx413), .A0 (nx2691), .A1 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_3), .S0 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx405)) ;
    inv01 ix2690 (.Y (nx2691), .A (CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx403)) ;
    mux21 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix424 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx423), .A0 (nx2693), .A1 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_4), .S0 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx415)) ;
    inv01 ix2692 (.Y (nx2693), .A (CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx413)) ;
    mux21 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix434 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx433), .A0 (nx2695), .A1 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_5), .S0 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx425)) ;
    inv01 ix2694 (.Y (nx2695), .A (CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx423)) ;
    mux21 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix444 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx443), .A0 (nx2697), .A1 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_6), .S0 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx435)) ;
    inv01 ix2696 (.Y (nx2697), .A (CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx433)) ;
    mux21 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix454 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx453), .A0 (nx2699), .A1 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_7), .S0 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx445)) ;
    inv01 ix2698 (.Y (nx2699), .A (CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx443)) ;
    mux21 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix462 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx461), .A0 (nx2701), .A1 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_8), .S0 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx455)) ;
    inv01 ix2700 (.Y (nx2701), .A (CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx453)) ;
    mux21 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix468 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx467), .A0 (nx2703), .A1 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_9), .S0 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx463)) ;
    inv01 ix2702 (.Y (nx2703), .A (CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx461)) ;
    mux21 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix476 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx475), .A0 (nx2705), .A1 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_10), .S0 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx471)) ;
    inv01 ix2704 (.Y (nx2705), .A (CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx467)) ;
    mux21 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix484 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx483), .A0 (nx2707), .A1 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_11), .S0 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx479)) ;
    inv01 ix2706 (.Y (nx2707), .A (CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx475)) ;
    mux21 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix492 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx491), .A0 (nx2709), .A1 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_12), .S0 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx487)) ;
    inv01 ix2708 (.Y (nx2709), .A (CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx483)) ;
    mux21 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix500 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx499), .A0 (nx2711), .A1 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_13), .S0 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx495)) ;
    inv01 ix2710 (.Y (nx2711), .A (CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx491)) ;
    mux21 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix508 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx507), .A0 (nx2713), .A1 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_14), .S0 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx503)) ;
    inv01 ix2712 (.Y (nx2713), .A (CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx499)) ;
    mux21 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix516 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx515), .A0 (nx2715), .A1 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_15), .S0 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx511)) ;
    inv01 ix2714 (.Y (nx2715), .A (CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx507)) ;
    mux21 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix161 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_1), .A0 (nx2717), .A1 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx379), .S0 (nx7679)) ;
    inv01 ix2716 (.Y (nx2717), .A (CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_1)) ;
    mux21 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix181 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_2), .A0 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx387), .A1 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx389), .S0 (nx7679)) ;
    mux21 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix201 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_3), .A0 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx399), .A1 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx401), .S0 (nx7679)) ;
    mux21 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix221 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_4), .A0 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx409), .A1 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx411), .S0 (nx7679)) ;
    mux21 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix241 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_5), .A0 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx419), .A1 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx421), .S0 (nx7679)) ;
    mux21 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix261 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_6), .A0 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx429), .A1 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx431), .S0 (nx7679)) ;
    mux21 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix281 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_7), .A0 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx439), .A1 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx441), .S0 (nx7679)) ;
    mux21 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix301 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_8), .A0 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx449), .A1 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx451), .S0 (nx7681)) ;
    mux21 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix321 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_9), .A0 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx469), .A1 (nx2719), .S0 (nx7681)) ;
    inv01 ix2718 (.Y (nx2719), .A (CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx316)) ;
    mux21 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix341 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_10), .A0 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx477), .A1 (nx2721), .S0 (nx7681)) ;
    inv01 ix2720 (.Y (nx2721), .A (CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx336)) ;
    mux21 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix361 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_11), .A0 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx485), .A1 (nx2723), .S0 (nx7681)) ;
    inv01 ix2722 (.Y (nx2723), .A (CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx356)) ;
    mux21 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix381 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_12), .A0 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx493), .A1 (nx2725), .S0 (nx7681)) ;
    inv01 ix2724 (.Y (nx2725), .A (CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx376)) ;
    mux21 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix401 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_13), .A0 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx501), .A1 (nx2727), .S0 (nx7681)) ;
    inv01 ix2726 (.Y (nx2727), .A (CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx396)) ;
    mux21 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix421 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_14), .A0 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx509), .A1 (nx2729), .S0 (nx7681)) ;
    inv01 ix2728 (.Y (nx2729), .A (CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx416)) ;
    mux21 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix441 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_15), .A0 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx517), .A1 (nx2731), .S0 (nx7683)) ;
    inv01 ix2730 (.Y (nx2731), .A (CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx436)) ;
    mux21 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_ix461 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_16), .A0 (nx2733), 
          .A1 (nx2735), .S0 (nx7683)) ;
    inv01 ix2732 (.Y (nx2733), .A (CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothP_16)
          ) ;
    inv01 ix2734 (.Y (nx2735), .A (CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx456)) ;
    nor02_2x CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix81 (.Y (
             CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx80), .A0 (Instr), .A1 (
             nx7309)) ;
    nor02_2x CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix319 (.Y (
             CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642), .A0 (
             CALCULATOR_Start_dup_1184), .A1 (
             CALCULATOR_CalculatingBooth_dup_1181)) ;
    nor02_2x CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix85 (.Y (
             CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_0), .A0 (
             nx7693), .A1 (nx2737)) ;
    inv01 ix2736 (.Y (nx2737), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_1)) ;
    mux21 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix125 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_1), .A0 (
          nx2739), .A1 (nx2741), .S0 (nx7693)) ;
    inv01 ix2738 (.Y (nx2739), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_2)) ;
    inv01 ix2740 (.Y (nx2741), .A (CacheWindow_1__3__0)) ;
    mux21 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix133 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_2), .A0 (
          nx2743), .A1 (nx2745), .S0 (nx7693)) ;
    inv01 ix2742 (.Y (nx2743), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_3)) ;
    inv01 ix2744 (.Y (nx2745), .A (CacheWindow_1__3__1)) ;
    mux21 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix141 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_3), .A0 (
          nx2747), .A1 (nx2749), .S0 (nx7693)) ;
    inv01 ix2746 (.Y (nx2747), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_4)) ;
    inv01 ix2748 (.Y (nx2749), .A (CacheWindow_1__3__2)) ;
    mux21 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix149 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_4), .A0 (
          nx2751), .A1 (nx2753), .S0 (nx7693)) ;
    inv01 ix2750 (.Y (nx2751), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_5)) ;
    inv01 ix2752 (.Y (nx2753), .A (CacheWindow_1__3__3)) ;
    mux21 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix157 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_5), .A0 (
          nx2755), .A1 (nx2757), .S0 (nx7693)) ;
    inv01 ix2754 (.Y (nx2755), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_6)) ;
    inv01 ix2756 (.Y (nx2757), .A (CacheWindow_1__3__4)) ;
    mux21 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix165 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_6), .A0 (
          nx2759), .A1 (nx2761), .S0 (nx7693)) ;
    inv01 ix2758 (.Y (nx2759), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_7)) ;
    inv01 ix2760 (.Y (nx2761), .A (CacheWindow_1__3__5)) ;
    mux21 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix173 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_7), .A0 (
          nx2763), .A1 (nx2765), .S0 (nx7695)) ;
    inv01 ix2762 (.Y (nx2763), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_8)) ;
    inv01 ix2764 (.Y (nx2765), .A (CacheWindow_1__3__6)) ;
    mux21 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix181 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_8), .A0 (
          nx2767), .A1 (nx2769), .S0 (nx7695)) ;
    inv01 ix2766 (.Y (nx2767), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_9)) ;
    inv01 ix2768 (.Y (nx2769), .A (CacheWindow_1__3__7)) ;
    nor02_2x CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix89 (.Y (
             CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_9), .A0 (
             nx7695), .A1 (nx2771)) ;
    inv01 ix2770 (.Y (nx2771), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_10)) ;
    nor02_2x CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix93 (.Y (
             CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_10), .A0 (
             nx7695), .A1 (nx2773)) ;
    inv01 ix2772 (.Y (nx2773), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_11)) ;
    nor02_2x CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix97 (.Y (
             CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_11), .A0 (
             nx7695), .A1 (nx2775)) ;
    inv01 ix2774 (.Y (nx2775), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_12)) ;
    nor02_2x CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix101 (.Y (
             CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_12), .A0 (
             nx7695), .A1 (nx2777)) ;
    inv01 ix2776 (.Y (nx2777), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_13)) ;
    nor02_2x CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix105 (.Y (
             CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_13), .A0 (
             nx7695), .A1 (nx2779)) ;
    inv01 ix2778 (.Y (nx2779), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_14)) ;
    nor02_2x CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix109 (.Y (
             CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_14), .A0 (
             nx7697), .A1 (nx2781)) ;
    inv01 ix2780 (.Y (nx2781), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_15)) ;
    nor02_2x CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix113 (.Y (
             CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_15), .A0 (
             nx7697), .A1 (nx2783)) ;
    inv01 ix2782 (.Y (nx2783), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_16)) ;
    nor02_2x CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix117 (.Y (
             CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_16), .A0 (
             nx7697), .A1 (nx2783)) ;
    mux21 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix189 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothOperand_0), .A0 (nx2785), .A1 (
          nx2787), .S0 (nx7685)) ;
    inv01 ix2784 (.Y (nx2785), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_0)) ;
    inv01 ix2786 (.Y (nx2787), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_0)) ;
    mux21 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix197 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothOperand_1), .A0 (nx2789), .A1 (
          nx2791), .S0 (nx7685)) ;
    inv01 ix2788 (.Y (nx2789), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_1)) ;
    inv01 ix2790 (.Y (nx2791), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_1)) ;
    mux21 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix205 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothOperand_2), .A0 (nx2793), .A1 (
          nx2795), .S0 (nx7685)) ;
    inv01 ix2792 (.Y (nx2793), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_2)) ;
    inv01 ix2794 (.Y (nx2795), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_2)) ;
    mux21 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix213 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothOperand_3), .A0 (nx2797), .A1 (
          nx2799), .S0 (nx7685)) ;
    inv01 ix2796 (.Y (nx2797), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_3)) ;
    inv01 ix2798 (.Y (nx2799), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_3)) ;
    mux21 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix221 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothOperand_4), .A0 (nx2801), .A1 (
          nx2803), .S0 (nx7685)) ;
    inv01 ix2800 (.Y (nx2801), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_4)) ;
    inv01 ix2802 (.Y (nx2803), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_4)) ;
    mux21 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix229 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothOperand_5), .A0 (nx2805), .A1 (
          nx2807), .S0 (nx7687)) ;
    inv01 ix2804 (.Y (nx2805), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_5)) ;
    inv01 ix2806 (.Y (nx2807), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_5)) ;
    mux21 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix237 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothOperand_6), .A0 (nx2809), .A1 (
          nx2811), .S0 (nx7687)) ;
    inv01 ix2808 (.Y (nx2809), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_6)) ;
    inv01 ix2810 (.Y (nx2811), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_6)) ;
    mux21 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix245 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothOperand_7), .A0 (nx2813), .A1 (
          nx2815), .S0 (nx7687)) ;
    inv01 ix2812 (.Y (nx2813), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_7)) ;
    inv01 ix2814 (.Y (nx2815), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_7)) ;
    mux21 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix253 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothOperand_8), .A0 (nx2817), .A1 (
          nx2819), .S0 (nx7687)) ;
    inv01 ix2816 (.Y (nx2817), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_8)) ;
    inv01 ix2818 (.Y (nx2819), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_8)) ;
    mux21 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix261 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothOperand_9), .A0 (nx2821), .A1 (
          nx2823), .S0 (nx7687)) ;
    inv01 ix2820 (.Y (nx2821), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_9)) ;
    inv01 ix2822 (.Y (nx2823), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_9)) ;
    mux21 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix269 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothOperand_10), .A0 (nx2825), .A1 (
          nx2827), .S0 (nx7687)) ;
    inv01 ix2824 (.Y (nx2825), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_10)) ;
    inv01 ix2826 (.Y (nx2827), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_10)) ;
    mux21 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix277 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothOperand_11), .A0 (nx2829), .A1 (
          nx2831), .S0 (nx7687)) ;
    inv01 ix2828 (.Y (nx2829), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_11)) ;
    inv01 ix2830 (.Y (nx2831), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_11)) ;
    mux21 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix285 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothOperand_12), .A0 (nx2833), .A1 (
          nx2835), .S0 (nx7689)) ;
    inv01 ix2832 (.Y (nx2833), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_12)) ;
    inv01 ix2834 (.Y (nx2835), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_12)) ;
    mux21 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix293 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothOperand_13), .A0 (nx2837), .A1 (
          nx2839), .S0 (nx7689)) ;
    inv01 ix2836 (.Y (nx2837), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_13)) ;
    inv01 ix2838 (.Y (nx2839), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_13)) ;
    mux21 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix301 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothOperand_14), .A0 (nx2841), .A1 (
          nx2843), .S0 (nx7689)) ;
    inv01 ix2840 (.Y (nx2841), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_14)) ;
    inv01 ix2842 (.Y (nx2843), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_14)) ;
    mux21 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix309 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothOperand_15), .A0 (nx2845), .A1 (
          nx2847), .S0 (nx7689)) ;
    inv01 ix2844 (.Y (nx2845), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_15)) ;
    inv01 ix2846 (.Y (nx2847), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_15)) ;
    mux21 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix317 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BoothOperand_16), .A0 (nx2849), .A1 (
          nx2851), .S0 (nx7689)) ;
    inv01 ix2848 (.Y (nx2849), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_16)) ;
    inv01 ix2850 (.Y (nx2851), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_16)) ;
    xnor2 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix321 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_AddPToBoothOperand), .A0 (nx7689), .A1 (
          nx2717)) ;
    oai32 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix393 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .A0 (
          nx8527), .A1 (RST), .A2 (nx7699), .B0 (nx2787), .B1 (nx2855)) ;
    oai32 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix403 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .A0 (
          nx8527), .A1 (RST), .A2 (nx7699), .B0 (nx2791), .B1 (nx2855)) ;
    oai32 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix413 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .A0 (
          nx8527), .A1 (RST), .A2 (nx7699), .B0 (nx2795), .B1 (nx2855)) ;
    oai32 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix423 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .A0 (
          nx8527), .A1 (RST), .A2 (nx7699), .B0 (nx2799), .B1 (nx2855)) ;
    oai32 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix433 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .A0 (
          nx8527), .A1 (RST), .A2 (nx7699), .B0 (nx2803), .B1 (nx2855)) ;
    oai32 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix443 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .A0 (
          nx8527), .A1 (RST), .A2 (nx7699), .B0 (nx2807), .B1 (nx2855)) ;
    oai32 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix453 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .A0 (
          nx8527), .A1 (RST), .A2 (nx7701), .B0 (nx2811), .B1 (nx2855)) ;
    oai32 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix463 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .A0 (
          nx8529), .A1 (RST), .A2 (nx7701), .B0 (nx2815), .B1 (nx2857)) ;
    oai32 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix473 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .A0 (
          nx8529), .A1 (RST), .A2 (nx7701), .B0 (nx2819), .B1 (nx2857)) ;
    oai32 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix483 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .A0 (
          nx2859), .A1 (RST), .A2 (nx7701), .B0 (nx2823), .B1 (nx2857)) ;
    inv01 ix2858 (.Y (nx2859), .A (CacheFilter_1__3__0)) ;
    oai32 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix493 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .A0 (
          nx2861), .A1 (RST), .A2 (nx7701), .B0 (nx2827), .B1 (nx2857)) ;
    inv01 ix2860 (.Y (nx2861), .A (CacheFilter_1__3__1)) ;
    oai32 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix503 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .A0 (
          nx2863), .A1 (RST), .A2 (nx7701), .B0 (nx2831), .B1 (nx2857)) ;
    inv01 ix2862 (.Y (nx2863), .A (CacheFilter_1__3__2)) ;
    oai32 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix513 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .A0 (
          nx2865), .A1 (RST), .A2 (nx7701), .B0 (nx2835), .B1 (nx2857)) ;
    inv01 ix2864 (.Y (nx2865), .A (CacheFilter_1__3__3)) ;
    oai32 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix523 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .A0 (
          nx2867), .A1 (RST), .A2 (nx7703), .B0 (nx2839), .B1 (nx2857)) ;
    inv01 ix2866 (.Y (nx2867), .A (CacheFilter_1__3__4)) ;
    oai32 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix533 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .A0 (
          nx2869), .A1 (RST), .A2 (nx7703), .B0 (nx2843), .B1 (nx2871)) ;
    inv01 ix2868 (.Y (nx2869), .A (CacheFilter_1__3__5)) ;
    inv01 ix2870 (.Y (nx2871), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566)) ;
    oai32 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix543 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .A0 (
          nx2873), .A1 (RST), .A2 (nx7703), .B0 (nx2847), .B1 (nx2871)) ;
    inv01 ix2872 (.Y (nx2873), .A (CacheFilter_1__3__6)) ;
    oai32 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix553 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .A0 (
          nx2875), .A1 (RST), .A2 (nx7703), .B0 (nx2851), .B1 (nx2871)) ;
    inv01 ix2874 (.Y (nx2875), .A (CacheFilter_1__3__7)) ;
    nand02_2x CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix633 (.Y (
              nx2855), .A0 (nx7351), .A1 (nx7703)) ;
    nand02_2x CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix635 (.Y (
              nx2857), .A0 (nx7351), .A1 (nx7703)) ;
    oai32 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix393 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .A0 (
          nx8529), .A1 (RST), .A2 (nx7705), .B0 (nx2785), .B1 (nx2877)) ;
    oai32 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix403 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .A0 (
          nx8529), .A1 (RST), .A2 (nx7705), .B0 (nx2789), .B1 (nx2877)) ;
    oai32 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix413 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .A0 (
          nx8529), .A1 (RST), .A2 (nx7705), .B0 (nx2793), .B1 (nx2877)) ;
    oai32 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix423 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .A0 (
          nx8529), .A1 (RST), .A2 (nx7705), .B0 (nx2797), .B1 (nx2877)) ;
    oai32 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix433 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .A0 (
          nx8529), .A1 (RST), .A2 (nx7705), .B0 (nx2801), .B1 (nx2877)) ;
    oai32 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix443 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .A0 (
          nx8531), .A1 (RST), .A2 (nx7705), .B0 (nx2805), .B1 (nx2877)) ;
    oai32 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix453 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .A0 (
          nx8531), .A1 (RST), .A2 (nx7707), .B0 (nx2809), .B1 (nx2877)) ;
    oai32 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix463 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .A0 (
          nx8531), .A1 (RST), .A2 (nx7707), .B0 (nx2813), .B1 (nx2879)) ;
    oai32 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix473 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .A0 (
          nx8531), .A1 (RST), .A2 (nx7707), .B0 (nx2817), .B1 (nx2879)) ;
    oai32 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix483 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .A0 (
          nx2859), .A1 (RST), .A2 (nx7707), .B0 (nx2821), .B1 (nx2879)) ;
    oai32 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix493 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .A0 (
          nx2881), .A1 (RST), .A2 (nx7707), .B0 (nx2825), .B1 (nx2879)) ;
    inv01 ix2880 (.Y (nx2881), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_10)) ;
    oai32 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix503 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .A0 (
          nx2883), .A1 (RST), .A2 (nx7707), .B0 (nx2829), .B1 (nx2879)) ;
    inv01 ix2882 (.Y (nx2883), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_11)) ;
    oai32 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix513 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .A0 (
          nx2885), .A1 (RST), .A2 (nx7707), .B0 (nx2833), .B1 (nx2879)) ;
    inv01 ix2884 (.Y (nx2885), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_12)) ;
    oai32 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix523 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .A0 (
          nx2887), .A1 (RST), .A2 (nx7709), .B0 (nx2837), .B1 (nx2879)) ;
    inv01 ix2886 (.Y (nx2887), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_13)) ;
    oai32 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix533 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .A0 (
          nx2889), .A1 (RST), .A2 (nx7709), .B0 (nx2841), .B1 (nx2891)) ;
    inv01 ix2888 (.Y (nx2889), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_14)) ;
    inv01 ix2890 (.Y (nx2891), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566)) ;
    oai32 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix543 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .A0 (
          nx2893), .A1 (RST), .A2 (nx7709), .B0 (nx2845), .B1 (nx2891)) ;
    inv01 ix2892 (.Y (nx2893), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_15)) ;
    oai32 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix553 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .A0 (
          nx2895), .A1 (RST), .A2 (nx7709), .B0 (nx2849), .B1 (nx2891)) ;
    inv01 ix2894 (.Y (nx2895), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_16)) ;
    nand02_2x CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix633 (.Y (
              nx2877), .A0 (nx7351), .A1 (nx7709)) ;
    nand02_2x CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix635 (.Y (
              nx2879), .A0 (nx7351), .A1 (nx7709)) ;
    oai32 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix393 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .A0 (
          nx2897), .A1 (RST), .A2 (nx7711), .B0 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx384), .B1 (nx2899)) ;
    inv01 ix2896 (.Y (nx2897), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_0)) ;
    oai32 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix403 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .A0 (
          nx2901), .A1 (RST), .A2 (nx7711), .B0 (nx2717), .B1 (nx2899)) ;
    inv01 ix2900 (.Y (nx2901), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_1)) ;
    oai32 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix413 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .A0 (
          nx2903), .A1 (RST), .A2 (nx7711), .B0 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx387), .B1 (nx2899)) ;
    inv01 ix2902 (.Y (nx2903), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_2)) ;
    oai32 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix423 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .A0 (
          nx2905), .A1 (RST), .A2 (nx7711), .B0 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx399), .B1 (nx2899)) ;
    inv01 ix2904 (.Y (nx2905), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_3)) ;
    oai32 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix433 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .A0 (
          nx2907), .A1 (RST), .A2 (nx7711), .B0 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx409), .B1 (nx2899)) ;
    inv01 ix2906 (.Y (nx2907), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_4)) ;
    oai32 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix443 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .A0 (
          nx2909), .A1 (RST), .A2 (nx7711), .B0 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx419), .B1 (nx2899)) ;
    inv01 ix2908 (.Y (nx2909), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_5)) ;
    oai32 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix453 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .A0 (
          nx2911), .A1 (RST), .A2 (nx7711), .B0 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx429), .B1 (nx2899)) ;
    inv01 ix2910 (.Y (nx2911), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_6)) ;
    oai32 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix463 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .A0 (
          nx2913), .A1 (RST), .A2 (nx7713), .B0 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx439), .B1 (nx2915)) ;
    inv01 ix2912 (.Y (nx2913), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_7)) ;
    oai32 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix473 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .A0 (
          nx2917), .A1 (RST), .A2 (nx7713), .B0 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx449), .B1 (nx2915)) ;
    inv01 ix2916 (.Y (nx2917), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_8)) ;
    oai32 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix483 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .A0 (
          nx2919), .A1 (RST), .A2 (nx7713), .B0 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx469), .B1 (nx2915)) ;
    inv01 ix2918 (.Y (nx2919), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_9)) ;
    oai32 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix493 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .A0 (
          nx2921), .A1 (RST), .A2 (nx7713), .B0 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx477), .B1 (nx2915)) ;
    inv01 ix2920 (.Y (nx2921), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_10)) ;
    oai32 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix503 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .A0 (
          nx2923), .A1 (RST), .A2 (nx7713), .B0 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx485), .B1 (nx2915)) ;
    inv01 ix2922 (.Y (nx2923), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_11)) ;
    oai32 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix513 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .A0 (
          nx2925), .A1 (RST), .A2 (nx7713), .B0 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx493), .B1 (nx2915)) ;
    inv01 ix2924 (.Y (nx2925), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_12)) ;
    oai32 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix523 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .A0 (
          nx2927), .A1 (RST), .A2 (nx7713), .B0 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx501), .B1 (nx2915)) ;
    inv01 ix2926 (.Y (nx2927), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_13)) ;
    oai32 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix533 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .A0 (
          nx2929), .A1 (RST), .A2 (nx7715), .B0 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx509), .B1 (nx2931)) ;
    inv01 ix2928 (.Y (nx2929), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_14)) ;
    inv01 ix2930 (.Y (nx2931), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566)) ;
    oai32 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix543 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .A0 (
          nx2933), .A1 (RST), .A2 (nx7715), .B0 (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_nx517), .B1 (nx2931)) ;
    inv01 ix2932 (.Y (nx2933), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_15)) ;
    oai32 CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix553 (.Y (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .A0 (
          nx2935), .A1 (RST), .A2 (nx7715), .B0 (nx2733), .B1 (nx2931)) ;
    inv01 ix2934 (.Y (nx2935), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_16)) ;
    nand02_2x CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix633 (.Y (
              nx2899), .A0 (nx7351), .A1 (nx7715)) ;
    nand02_2x CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix635 (.Y (
              nx2915), .A0 (nx7351), .A1 (nx7715)) ;
    mux21 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix404 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx403), .A0 (nx2937), .A1 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_2), .S0 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx395)) ;
    inv01 ix2936 (.Y (nx2937), .A (CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx391)) ;
    mux21 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix414 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx413), .A0 (nx2939), .A1 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_3), .S0 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx405)) ;
    inv01 ix2938 (.Y (nx2939), .A (CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx403)) ;
    mux21 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix424 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx423), .A0 (nx2941), .A1 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_4), .S0 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx415)) ;
    inv01 ix2940 (.Y (nx2941), .A (CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx413)) ;
    mux21 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix434 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx433), .A0 (nx2943), .A1 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_5), .S0 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx425)) ;
    inv01 ix2942 (.Y (nx2943), .A (CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx423)) ;
    mux21 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix444 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx443), .A0 (nx2945), .A1 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_6), .S0 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx435)) ;
    inv01 ix2944 (.Y (nx2945), .A (CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx433)) ;
    mux21 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix454 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx453), .A0 (nx2947), .A1 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_7), .S0 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx445)) ;
    inv01 ix2946 (.Y (nx2947), .A (CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx443)) ;
    mux21 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix462 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx461), .A0 (nx2949), .A1 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_8), .S0 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx455)) ;
    inv01 ix2948 (.Y (nx2949), .A (CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx453)) ;
    mux21 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix468 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx467), .A0 (nx2951), .A1 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_9), .S0 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx463)) ;
    inv01 ix2950 (.Y (nx2951), .A (CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx461)) ;
    mux21 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix476 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx475), .A0 (nx2953), .A1 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_10), .S0 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx471)) ;
    inv01 ix2952 (.Y (nx2953), .A (CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx467)) ;
    mux21 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix484 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx483), .A0 (nx2955), .A1 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_11), .S0 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx479)) ;
    inv01 ix2954 (.Y (nx2955), .A (CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx475)) ;
    mux21 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix492 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx491), .A0 (nx2957), .A1 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_12), .S0 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx487)) ;
    inv01 ix2956 (.Y (nx2957), .A (CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx483)) ;
    mux21 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix500 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx499), .A0 (nx2959), .A1 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_13), .S0 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx495)) ;
    inv01 ix2958 (.Y (nx2959), .A (CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx491)) ;
    mux21 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix508 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx507), .A0 (nx2961), .A1 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_14), .S0 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx503)) ;
    inv01 ix2960 (.Y (nx2961), .A (CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx499)) ;
    mux21 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix516 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx515), .A0 (nx2963), .A1 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_15), .S0 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx511)) ;
    inv01 ix2962 (.Y (nx2963), .A (CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx507)) ;
    mux21 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix161 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_1), .A0 (nx2965), .A1 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx379), .S0 (nx7719)) ;
    inv01 ix2964 (.Y (nx2965), .A (CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_1)) ;
    mux21 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix181 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_2), .A0 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx387), .A1 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx389), .S0 (nx7719)) ;
    mux21 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix201 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_3), .A0 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx399), .A1 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx401), .S0 (nx7719)) ;
    mux21 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix221 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_4), .A0 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx409), .A1 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx411), .S0 (nx7719)) ;
    mux21 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix241 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_5), .A0 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx419), .A1 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx421), .S0 (nx7719)) ;
    mux21 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix261 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_6), .A0 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx429), .A1 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx431), .S0 (nx7719)) ;
    mux21 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix281 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_7), .A0 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx439), .A1 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx441), .S0 (nx7719)) ;
    mux21 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix301 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_8), .A0 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx449), .A1 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx451), .S0 (nx7721)) ;
    mux21 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix321 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_9), .A0 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx469), .A1 (nx2967), .S0 (nx7721)) ;
    inv01 ix2966 (.Y (nx2967), .A (CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx316)) ;
    mux21 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix341 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_10), .A0 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx477), .A1 (nx2969), .S0 (nx7721)) ;
    inv01 ix2968 (.Y (nx2969), .A (CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx336)) ;
    mux21 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix361 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_11), .A0 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx485), .A1 (nx2971), .S0 (nx7721)) ;
    inv01 ix2970 (.Y (nx2971), .A (CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx356)) ;
    mux21 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix381 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_12), .A0 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx493), .A1 (nx2973), .S0 (nx7721)) ;
    inv01 ix2972 (.Y (nx2973), .A (CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx376)) ;
    mux21 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix401 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_13), .A0 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx501), .A1 (nx2975), .S0 (nx7721)) ;
    inv01 ix2974 (.Y (nx2975), .A (CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx396)) ;
    mux21 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix421 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_14), .A0 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx509), .A1 (nx2977), .S0 (nx7721)) ;
    inv01 ix2976 (.Y (nx2977), .A (CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx416)) ;
    mux21 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix441 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_15), .A0 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx517), .A1 (nx2979), .S0 (nx7723)) ;
    inv01 ix2978 (.Y (nx2979), .A (CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx436)) ;
    mux21 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_ix461 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_16), .A0 (nx2981), 
          .A1 (nx2983), .S0 (nx7723)) ;
    inv01 ix2980 (.Y (nx2981), .A (CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothP_16)
          ) ;
    inv01 ix2982 (.Y (nx2983), .A (CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx456)) ;
    nor02_2x CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix81 (.Y (
             CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx80), .A0 (Instr), .A1 (
             nx7309)) ;
    nor02_2x CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix319 (.Y (
             CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642), .A0 (
             CALCULATOR_Start_dup_1189), .A1 (
             CALCULATOR_CalculatingBooth_dup_1181)) ;
    nor02_2x CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix85 (.Y (
             CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_0), .A0 (
             nx7733), .A1 (nx2985)) ;
    inv01 ix2984 (.Y (nx2985), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_1)) ;
    mux21 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix125 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_1), .A0 (
          nx2987), .A1 (nx2989), .S0 (nx7733)) ;
    inv01 ix2986 (.Y (nx2987), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_2)) ;
    inv01 ix2988 (.Y (nx2989), .A (CacheWindow_1__4__0)) ;
    mux21 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix133 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_2), .A0 (
          nx2991), .A1 (nx2993), .S0 (nx7733)) ;
    inv01 ix2990 (.Y (nx2991), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_3)) ;
    inv01 ix2992 (.Y (nx2993), .A (CacheWindow_1__4__1)) ;
    mux21 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix141 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_3), .A0 (
          nx2995), .A1 (nx2997), .S0 (nx7733)) ;
    inv01 ix2994 (.Y (nx2995), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_4)) ;
    inv01 ix2996 (.Y (nx2997), .A (CacheWindow_1__4__2)) ;
    mux21 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix149 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_4), .A0 (
          nx2999), .A1 (nx3001), .S0 (nx7733)) ;
    inv01 ix2998 (.Y (nx2999), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_5)) ;
    inv01 ix3000 (.Y (nx3001), .A (CacheWindow_1__4__3)) ;
    mux21 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix157 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_5), .A0 (
          nx3003), .A1 (nx3005), .S0 (nx7733)) ;
    inv01 ix3002 (.Y (nx3003), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_6)) ;
    inv01 ix3004 (.Y (nx3005), .A (CacheWindow_1__4__4)) ;
    mux21 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix165 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_6), .A0 (
          nx3007), .A1 (nx3009), .S0 (nx7733)) ;
    inv01 ix3006 (.Y (nx3007), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_7)) ;
    inv01 ix3008 (.Y (nx3009), .A (CacheWindow_1__4__5)) ;
    mux21 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix173 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_7), .A0 (
          nx3011), .A1 (nx3013), .S0 (nx7735)) ;
    inv01 ix3010 (.Y (nx3011), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_8)) ;
    inv01 ix3012 (.Y (nx3013), .A (CacheWindow_1__4__6)) ;
    mux21 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix181 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_8), .A0 (
          nx3015), .A1 (nx3017), .S0 (nx7735)) ;
    inv01 ix3014 (.Y (nx3015), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_9)) ;
    inv01 ix3016 (.Y (nx3017), .A (CacheWindow_1__4__7)) ;
    nor02_2x CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix89 (.Y (
             CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_9), .A0 (
             nx7735), .A1 (nx3019)) ;
    inv01 ix3018 (.Y (nx3019), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_10)) ;
    nor02_2x CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix93 (.Y (
             CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_10), .A0 (
             nx7735), .A1 (nx3021)) ;
    inv01 ix3020 (.Y (nx3021), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_11)) ;
    nor02_2x CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix97 (.Y (
             CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_11), .A0 (
             nx7735), .A1 (nx3023)) ;
    inv01 ix3022 (.Y (nx3023), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_12)) ;
    nor02_2x CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix101 (.Y (
             CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_12), .A0 (
             nx7735), .A1 (nx3025)) ;
    inv01 ix3024 (.Y (nx3025), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_13)) ;
    nor02_2x CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix105 (.Y (
             CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_13), .A0 (
             nx7735), .A1 (nx3027)) ;
    inv01 ix3026 (.Y (nx3027), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_14)) ;
    nor02_2x CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix109 (.Y (
             CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_14), .A0 (
             nx7737), .A1 (nx3029)) ;
    inv01 ix3028 (.Y (nx3029), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_15)) ;
    nor02_2x CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix113 (.Y (
             CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_15), .A0 (
             nx7737), .A1 (nx3031)) ;
    inv01 ix3030 (.Y (nx3031), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_16)) ;
    nor02_2x CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix117 (.Y (
             CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_16), .A0 (
             nx7737), .A1 (nx3031)) ;
    mux21 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix189 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothOperand_0), .A0 (nx3033), .A1 (
          nx3035), .S0 (nx7725)) ;
    inv01 ix3032 (.Y (nx3033), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_0)) ;
    inv01 ix3034 (.Y (nx3035), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_0)) ;
    mux21 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix197 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothOperand_1), .A0 (nx3037), .A1 (
          nx3039), .S0 (nx7725)) ;
    inv01 ix3036 (.Y (nx3037), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_1)) ;
    inv01 ix3038 (.Y (nx3039), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_1)) ;
    mux21 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix205 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothOperand_2), .A0 (nx3041), .A1 (
          nx3043), .S0 (nx7725)) ;
    inv01 ix3040 (.Y (nx3041), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_2)) ;
    inv01 ix3042 (.Y (nx3043), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_2)) ;
    mux21 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix213 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothOperand_3), .A0 (nx3045), .A1 (
          nx3047), .S0 (nx7725)) ;
    inv01 ix3044 (.Y (nx3045), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_3)) ;
    inv01 ix3046 (.Y (nx3047), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_3)) ;
    mux21 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix221 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothOperand_4), .A0 (nx3049), .A1 (
          nx3051), .S0 (nx7725)) ;
    inv01 ix3048 (.Y (nx3049), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_4)) ;
    inv01 ix3050 (.Y (nx3051), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_4)) ;
    mux21 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix229 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothOperand_5), .A0 (nx3053), .A1 (
          nx3055), .S0 (nx7727)) ;
    inv01 ix3052 (.Y (nx3053), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_5)) ;
    inv01 ix3054 (.Y (nx3055), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_5)) ;
    mux21 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix237 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothOperand_6), .A0 (nx3057), .A1 (
          nx3059), .S0 (nx7727)) ;
    inv01 ix3056 (.Y (nx3057), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_6)) ;
    inv01 ix3058 (.Y (nx3059), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_6)) ;
    mux21 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix245 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothOperand_7), .A0 (nx3061), .A1 (
          nx3063), .S0 (nx7727)) ;
    inv01 ix3060 (.Y (nx3061), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_7)) ;
    inv01 ix3062 (.Y (nx3063), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_7)) ;
    mux21 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix253 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothOperand_8), .A0 (nx3065), .A1 (
          nx3067), .S0 (nx7727)) ;
    inv01 ix3064 (.Y (nx3065), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_8)) ;
    inv01 ix3066 (.Y (nx3067), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_8)) ;
    mux21 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix261 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothOperand_9), .A0 (nx3069), .A1 (
          nx3071), .S0 (nx7727)) ;
    inv01 ix3068 (.Y (nx3069), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_9)) ;
    inv01 ix3070 (.Y (nx3071), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_9)) ;
    mux21 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix269 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothOperand_10), .A0 (nx3073), .A1 (
          nx3075), .S0 (nx7727)) ;
    inv01 ix3072 (.Y (nx3073), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_10)) ;
    inv01 ix3074 (.Y (nx3075), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_10)) ;
    mux21 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix277 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothOperand_11), .A0 (nx3077), .A1 (
          nx3079), .S0 (nx7727)) ;
    inv01 ix3076 (.Y (nx3077), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_11)) ;
    inv01 ix3078 (.Y (nx3079), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_11)) ;
    mux21 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix285 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothOperand_12), .A0 (nx3081), .A1 (
          nx3083), .S0 (nx7729)) ;
    inv01 ix3080 (.Y (nx3081), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_12)) ;
    inv01 ix3082 (.Y (nx3083), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_12)) ;
    mux21 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix293 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothOperand_13), .A0 (nx3085), .A1 (
          nx3087), .S0 (nx7729)) ;
    inv01 ix3084 (.Y (nx3085), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_13)) ;
    inv01 ix3086 (.Y (nx3087), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_13)) ;
    mux21 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix301 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothOperand_14), .A0 (nx3089), .A1 (
          nx3091), .S0 (nx7729)) ;
    inv01 ix3088 (.Y (nx3089), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_14)) ;
    inv01 ix3090 (.Y (nx3091), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_14)) ;
    mux21 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix309 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothOperand_15), .A0 (nx3093), .A1 (
          nx3095), .S0 (nx7729)) ;
    inv01 ix3092 (.Y (nx3093), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_15)) ;
    inv01 ix3094 (.Y (nx3095), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_15)) ;
    mux21 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix317 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BoothOperand_16), .A0 (nx3097), .A1 (
          nx3099), .S0 (nx7729)) ;
    inv01 ix3096 (.Y (nx3097), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_16)) ;
    inv01 ix3098 (.Y (nx3099), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_16)) ;
    xnor2 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix321 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_AddPToBoothOperand), .A0 (nx7729), .A1 (
          nx2965)) ;
    oai32 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix393 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .A0 (
          nx8533), .A1 (RST), .A2 (nx7739), .B0 (nx3035), .B1 (nx3103)) ;
    oai32 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix403 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .A0 (
          nx8533), .A1 (RST), .A2 (nx7739), .B0 (nx3039), .B1 (nx3103)) ;
    oai32 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix413 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .A0 (
          nx8533), .A1 (RST), .A2 (nx7739), .B0 (nx3043), .B1 (nx3103)) ;
    oai32 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix423 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .A0 (
          nx8533), .A1 (RST), .A2 (nx7739), .B0 (nx3047), .B1 (nx3103)) ;
    oai32 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix433 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .A0 (
          nx8533), .A1 (RST), .A2 (nx7739), .B0 (nx3051), .B1 (nx3103)) ;
    oai32 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix443 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .A0 (
          nx8533), .A1 (RST), .A2 (nx7739), .B0 (nx3055), .B1 (nx3103)) ;
    oai32 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix453 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .A0 (
          nx8533), .A1 (RST), .A2 (nx7741), .B0 (nx3059), .B1 (nx3103)) ;
    oai32 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix463 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .A0 (
          nx8535), .A1 (RST), .A2 (nx7741), .B0 (nx3063), .B1 (nx3105)) ;
    oai32 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix473 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .A0 (
          nx8535), .A1 (RST), .A2 (nx7741), .B0 (nx3067), .B1 (nx3105)) ;
    oai32 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix483 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .A0 (
          nx3107), .A1 (RST), .A2 (nx7741), .B0 (nx3071), .B1 (nx3105)) ;
    inv01 ix3106 (.Y (nx3107), .A (CacheFilter_1__4__0)) ;
    oai32 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix493 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .A0 (
          nx3109), .A1 (RST), .A2 (nx7741), .B0 (nx3075), .B1 (nx3105)) ;
    inv01 ix3108 (.Y (nx3109), .A (CacheFilter_1__4__1)) ;
    oai32 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix503 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .A0 (
          nx3111), .A1 (RST), .A2 (nx7741), .B0 (nx3079), .B1 (nx3105)) ;
    inv01 ix3110 (.Y (nx3111), .A (CacheFilter_1__4__2)) ;
    oai32 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix513 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .A0 (
          nx3113), .A1 (RST), .A2 (nx7741), .B0 (nx3083), .B1 (nx3105)) ;
    inv01 ix3112 (.Y (nx3113), .A (CacheFilter_1__4__3)) ;
    oai32 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix523 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .A0 (
          nx3115), .A1 (RST), .A2 (nx7743), .B0 (nx3087), .B1 (nx3105)) ;
    inv01 ix3114 (.Y (nx3115), .A (CacheFilter_1__4__4)) ;
    oai32 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix533 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .A0 (
          nx3117), .A1 (RST), .A2 (nx7743), .B0 (nx3091), .B1 (nx3119)) ;
    inv01 ix3116 (.Y (nx3117), .A (CacheFilter_1__4__5)) ;
    inv01 ix3118 (.Y (nx3119), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566)) ;
    oai32 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix543 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .A0 (
          nx3121), .A1 (RST), .A2 (nx7743), .B0 (nx3095), .B1 (nx3119)) ;
    inv01 ix3120 (.Y (nx3121), .A (CacheFilter_1__4__6)) ;
    oai32 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix553 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .A0 (
          nx3123), .A1 (RST), .A2 (nx7743), .B0 (nx3099), .B1 (nx3119)) ;
    inv01 ix3122 (.Y (nx3123), .A (CacheFilter_1__4__7)) ;
    nand02_2x CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix633 (.Y (
              nx3103), .A0 (nx7351), .A1 (nx7743)) ;
    nand02_2x CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix635 (.Y (
              nx3105), .A0 (nx7353), .A1 (nx7743)) ;
    oai32 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix393 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .A0 (
          nx8535), .A1 (RST), .A2 (nx7745), .B0 (nx3033), .B1 (nx3125)) ;
    oai32 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix403 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .A0 (
          nx8535), .A1 (RST), .A2 (nx7745), .B0 (nx3037), .B1 (nx3125)) ;
    oai32 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix413 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .A0 (
          nx8535), .A1 (RST), .A2 (nx7745), .B0 (nx3041), .B1 (nx3125)) ;
    oai32 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix423 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .A0 (
          nx8535), .A1 (RST), .A2 (nx7745), .B0 (nx3045), .B1 (nx3125)) ;
    oai32 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix433 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .A0 (
          nx8535), .A1 (RST), .A2 (nx7745), .B0 (nx3049), .B1 (nx3125)) ;
    oai32 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix443 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .A0 (
          nx8537), .A1 (RST), .A2 (nx7745), .B0 (nx3053), .B1 (nx3125)) ;
    oai32 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix453 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .A0 (
          nx8537), .A1 (RST), .A2 (nx7747), .B0 (nx3057), .B1 (nx3125)) ;
    oai32 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix463 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .A0 (
          nx8537), .A1 (RST), .A2 (nx7747), .B0 (nx3061), .B1 (nx3127)) ;
    oai32 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix473 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .A0 (
          nx8537), .A1 (RST), .A2 (nx7747), .B0 (nx3065), .B1 (nx3127)) ;
    oai32 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix483 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .A0 (
          nx3107), .A1 (RST), .A2 (nx7747), .B0 (nx3069), .B1 (nx3127)) ;
    oai32 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix493 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .A0 (
          nx3129), .A1 (RST), .A2 (nx7747), .B0 (nx3073), .B1 (nx3127)) ;
    inv01 ix3128 (.Y (nx3129), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_10)) ;
    oai32 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix503 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .A0 (
          nx3131), .A1 (RST), .A2 (nx7747), .B0 (nx3077), .B1 (nx3127)) ;
    inv01 ix3130 (.Y (nx3131), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_11)) ;
    oai32 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix513 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .A0 (
          nx3133), .A1 (RST), .A2 (nx7747), .B0 (nx3081), .B1 (nx3127)) ;
    inv01 ix3132 (.Y (nx3133), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_12)) ;
    oai32 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix523 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .A0 (
          nx3135), .A1 (RST), .A2 (nx7749), .B0 (nx3085), .B1 (nx3127)) ;
    inv01 ix3134 (.Y (nx3135), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_13)) ;
    oai32 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix533 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .A0 (
          nx3137), .A1 (RST), .A2 (nx7749), .B0 (nx3089), .B1 (nx3139)) ;
    inv01 ix3136 (.Y (nx3137), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_14)) ;
    inv01 ix3138 (.Y (nx3139), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566)) ;
    oai32 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix543 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .A0 (
          nx3141), .A1 (RST), .A2 (nx7749), .B0 (nx3093), .B1 (nx3139)) ;
    inv01 ix3140 (.Y (nx3141), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_15)) ;
    oai32 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix553 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .A0 (
          nx3143), .A1 (RST), .A2 (nx7749), .B0 (nx3097), .B1 (nx3139)) ;
    inv01 ix3142 (.Y (nx3143), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_16)) ;
    nand02_2x CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix633 (.Y (
              nx3125), .A0 (nx7353), .A1 (nx7749)) ;
    nand02_2x CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix635 (.Y (
              nx3127), .A0 (nx7353), .A1 (nx7749)) ;
    oai32 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix393 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .A0 (
          nx3145), .A1 (RST), .A2 (nx7751), .B0 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx384), .B1 (nx3147)) ;
    inv01 ix3144 (.Y (nx3145), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_0)) ;
    oai32 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix403 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .A0 (
          nx3149), .A1 (RST), .A2 (nx7751), .B0 (nx2965), .B1 (nx3147)) ;
    inv01 ix3148 (.Y (nx3149), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_1)) ;
    oai32 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix413 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .A0 (
          nx3151), .A1 (RST), .A2 (nx7751), .B0 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx387), .B1 (nx3147)) ;
    inv01 ix3150 (.Y (nx3151), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_2)) ;
    oai32 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix423 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .A0 (
          nx3153), .A1 (RST), .A2 (nx7751), .B0 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx399), .B1 (nx3147)) ;
    inv01 ix3152 (.Y (nx3153), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_3)) ;
    oai32 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix433 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .A0 (
          nx3155), .A1 (RST), .A2 (nx7751), .B0 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx409), .B1 (nx3147)) ;
    inv01 ix3154 (.Y (nx3155), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_4)) ;
    oai32 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix443 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .A0 (
          nx3157), .A1 (RST), .A2 (nx7751), .B0 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx419), .B1 (nx3147)) ;
    inv01 ix3156 (.Y (nx3157), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_5)) ;
    oai32 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix453 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .A0 (
          nx3159), .A1 (RST), .A2 (nx7751), .B0 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx429), .B1 (nx3147)) ;
    inv01 ix3158 (.Y (nx3159), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_6)) ;
    oai32 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix463 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .A0 (
          nx3161), .A1 (RST), .A2 (nx7753), .B0 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx439), .B1 (nx3163)) ;
    inv01 ix3160 (.Y (nx3161), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_7)) ;
    oai32 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix473 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .A0 (
          nx3165), .A1 (RST), .A2 (nx7753), .B0 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx449), .B1 (nx3163)) ;
    inv01 ix3164 (.Y (nx3165), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_8)) ;
    oai32 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix483 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .A0 (
          nx3167), .A1 (RST), .A2 (nx7753), .B0 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx469), .B1 (nx3163)) ;
    inv01 ix3166 (.Y (nx3167), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_9)) ;
    oai32 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix493 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .A0 (
          nx3169), .A1 (RST), .A2 (nx7753), .B0 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx477), .B1 (nx3163)) ;
    inv01 ix3168 (.Y (nx3169), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_10)) ;
    oai32 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix503 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .A0 (
          nx3171), .A1 (RST), .A2 (nx7753), .B0 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx485), .B1 (nx3163)) ;
    inv01 ix3170 (.Y (nx3171), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_11)) ;
    oai32 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix513 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .A0 (
          nx3173), .A1 (RST), .A2 (nx7753), .B0 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx493), .B1 (nx3163)) ;
    inv01 ix3172 (.Y (nx3173), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_12)) ;
    oai32 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix523 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .A0 (
          nx3175), .A1 (RST), .A2 (nx7753), .B0 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx501), .B1 (nx3163)) ;
    inv01 ix3174 (.Y (nx3175), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_13)) ;
    oai32 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix533 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .A0 (
          nx3177), .A1 (RST), .A2 (nx7755), .B0 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx509), .B1 (nx3179)) ;
    inv01 ix3176 (.Y (nx3177), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_14)) ;
    inv01 ix3178 (.Y (nx3179), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566)) ;
    oai32 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix543 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .A0 (
          nx3181), .A1 (RST), .A2 (nx7755), .B0 (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_nx517), .B1 (nx3179)) ;
    inv01 ix3180 (.Y (nx3181), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_15)) ;
    oai32 CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix553 (.Y (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .A0 (
          nx3183), .A1 (RST), .A2 (nx7755), .B0 (nx2981), .B1 (nx3179)) ;
    inv01 ix3182 (.Y (nx3183), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_16)) ;
    nand02_2x CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix633 (.Y (
              nx3147), .A0 (nx7353), .A1 (nx7755)) ;
    nand02_2x CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix635 (.Y (
              nx3163), .A0 (nx7353), .A1 (nx7755)) ;
    mux21 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix404 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx403), .A0 (nx3185), .A1 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_2), .S0 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx395)) ;
    inv01 ix3184 (.Y (nx3185), .A (CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx391)) ;
    mux21 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix414 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx413), .A0 (nx3187), .A1 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_3), .S0 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx405)) ;
    inv01 ix3186 (.Y (nx3187), .A (CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx403)) ;
    mux21 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix424 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx423), .A0 (nx3189), .A1 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_4), .S0 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx415)) ;
    inv01 ix3188 (.Y (nx3189), .A (CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx413)) ;
    mux21 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix434 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx433), .A0 (nx3191), .A1 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_5), .S0 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx425)) ;
    inv01 ix3190 (.Y (nx3191), .A (CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx423)) ;
    mux21 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix444 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx443), .A0 (nx3193), .A1 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_6), .S0 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx435)) ;
    inv01 ix3192 (.Y (nx3193), .A (CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx433)) ;
    mux21 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix454 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx453), .A0 (nx3195), .A1 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_7), .S0 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx445)) ;
    inv01 ix3194 (.Y (nx3195), .A (CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx443)) ;
    mux21 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix462 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx461), .A0 (nx3197), .A1 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_8), .S0 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx455)) ;
    inv01 ix3196 (.Y (nx3197), .A (CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx453)) ;
    mux21 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix468 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx467), .A0 (nx3199), .A1 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_9), .S0 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx463)) ;
    inv01 ix3198 (.Y (nx3199), .A (CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx461)) ;
    mux21 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix476 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx475), .A0 (nx3201), .A1 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_10), .S0 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx471)) ;
    inv01 ix3200 (.Y (nx3201), .A (CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx467)) ;
    mux21 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix484 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx483), .A0 (nx3203), .A1 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_11), .S0 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx479)) ;
    inv01 ix3202 (.Y (nx3203), .A (CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx475)) ;
    mux21 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix492 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx491), .A0 (nx3205), .A1 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_12), .S0 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx487)) ;
    inv01 ix3204 (.Y (nx3205), .A (CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx483)) ;
    mux21 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix500 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx499), .A0 (nx3207), .A1 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_13), .S0 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx495)) ;
    inv01 ix3206 (.Y (nx3207), .A (CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx491)) ;
    mux21 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix508 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx507), .A0 (nx3209), .A1 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_14), .S0 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx503)) ;
    inv01 ix3208 (.Y (nx3209), .A (CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx499)) ;
    mux21 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix516 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx515), .A0 (nx3211), .A1 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_15), .S0 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx511)) ;
    inv01 ix3210 (.Y (nx3211), .A (CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx507)) ;
    mux21 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix161 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_1), .A0 (nx3213), .A1 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx379), .S0 (nx7759)) ;
    inv01 ix3212 (.Y (nx3213), .A (CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_1)) ;
    mux21 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix181 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_2), .A0 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx387), .A1 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx389), .S0 (nx7759)) ;
    mux21 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix201 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_3), .A0 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx399), .A1 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx401), .S0 (nx7759)) ;
    mux21 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix221 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_4), .A0 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx409), .A1 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx411), .S0 (nx7759)) ;
    mux21 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix241 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_5), .A0 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx419), .A1 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx421), .S0 (nx7759)) ;
    mux21 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix261 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_6), .A0 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx429), .A1 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx431), .S0 (nx7759)) ;
    mux21 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix281 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_7), .A0 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx439), .A1 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx441), .S0 (nx7759)) ;
    mux21 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix301 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_8), .A0 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx449), .A1 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx451), .S0 (nx7761)) ;
    mux21 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix321 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_9), .A0 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx469), .A1 (nx3215), .S0 (nx7761)) ;
    inv01 ix3214 (.Y (nx3215), .A (CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx316)) ;
    mux21 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix341 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_10), .A0 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx477), .A1 (nx3217), .S0 (nx7761)) ;
    inv01 ix3216 (.Y (nx3217), .A (CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx336)) ;
    mux21 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix361 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_11), .A0 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx485), .A1 (nx3219), .S0 (nx7761)) ;
    inv01 ix3218 (.Y (nx3219), .A (CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx356)) ;
    mux21 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix381 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_12), .A0 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx493), .A1 (nx3221), .S0 (nx7761)) ;
    inv01 ix3220 (.Y (nx3221), .A (CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx376)) ;
    mux21 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix401 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_13), .A0 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx501), .A1 (nx3223), .S0 (nx7761)) ;
    inv01 ix3222 (.Y (nx3223), .A (CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx396)) ;
    mux21 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix421 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_14), .A0 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx509), .A1 (nx3225), .S0 (nx7761)) ;
    inv01 ix3224 (.Y (nx3225), .A (CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx416)) ;
    mux21 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix441 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_15), .A0 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx517), .A1 (nx3227), .S0 (nx7763)) ;
    inv01 ix3226 (.Y (nx3227), .A (CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx436)) ;
    mux21 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_ix461 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_16), .A0 (nx3229), 
          .A1 (nx3231), .S0 (nx7763)) ;
    inv01 ix3228 (.Y (nx3229), .A (CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothP_16)
          ) ;
    inv01 ix3230 (.Y (nx3231), .A (CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx456)) ;
    nor02_2x CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix81 (.Y (
             CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx80), .A0 (Instr), .A1 (
             nx7309)) ;
    nor02_2x CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix319 (.Y (
             CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642), .A0 (
             CALCULATOR_Start_dup_1194), .A1 (
             CALCULATOR_CalculatingBooth_dup_1181)) ;
    nor02_2x CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix85 (.Y (
             CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_0), .A0 (
             nx7773), .A1 (nx3233)) ;
    inv01 ix3232 (.Y (nx3233), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_1)) ;
    mux21 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix125 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_1), .A0 (
          nx3235), .A1 (nx3237), .S0 (nx7773)) ;
    inv01 ix3234 (.Y (nx3235), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_2)) ;
    inv01 ix3236 (.Y (nx3237), .A (CacheWindow_2__0__0)) ;
    mux21 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix133 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_2), .A0 (
          nx3239), .A1 (nx3241), .S0 (nx7773)) ;
    inv01 ix3238 (.Y (nx3239), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_3)) ;
    inv01 ix3240 (.Y (nx3241), .A (CacheWindow_2__0__1)) ;
    mux21 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix141 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_3), .A0 (
          nx3243), .A1 (nx3245), .S0 (nx7773)) ;
    inv01 ix3242 (.Y (nx3243), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_4)) ;
    inv01 ix3244 (.Y (nx3245), .A (CacheWindow_2__0__2)) ;
    mux21 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix149 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_4), .A0 (
          nx3247), .A1 (nx3249), .S0 (nx7773)) ;
    inv01 ix3246 (.Y (nx3247), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_5)) ;
    inv01 ix3248 (.Y (nx3249), .A (CacheWindow_2__0__3)) ;
    mux21 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix157 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_5), .A0 (
          nx3251), .A1 (nx3253), .S0 (nx7773)) ;
    inv01 ix3250 (.Y (nx3251), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_6)) ;
    inv01 ix3252 (.Y (nx3253), .A (CacheWindow_2__0__4)) ;
    mux21 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix165 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_6), .A0 (
          nx3255), .A1 (nx3257), .S0 (nx7773)) ;
    inv01 ix3254 (.Y (nx3255), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_7)) ;
    inv01 ix3256 (.Y (nx3257), .A (CacheWindow_2__0__5)) ;
    mux21 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix173 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_7), .A0 (
          nx3259), .A1 (nx3261), .S0 (nx7775)) ;
    inv01 ix3258 (.Y (nx3259), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_8)) ;
    inv01 ix3260 (.Y (nx3261), .A (CacheWindow_2__0__6)) ;
    mux21 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix181 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_8), .A0 (
          nx3263), .A1 (nx3265), .S0 (nx7775)) ;
    inv01 ix3262 (.Y (nx3263), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_9)) ;
    inv01 ix3264 (.Y (nx3265), .A (CacheWindow_2__0__7)) ;
    nor02_2x CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix89 (.Y (
             CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_9), .A0 (
             nx7775), .A1 (nx3267)) ;
    inv01 ix3266 (.Y (nx3267), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_10)) ;
    nor02_2x CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix93 (.Y (
             CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_10), .A0 (
             nx7775), .A1 (nx3269)) ;
    inv01 ix3268 (.Y (nx3269), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_11)) ;
    nor02_2x CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix97 (.Y (
             CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_11), .A0 (
             nx7775), .A1 (nx3271)) ;
    inv01 ix3270 (.Y (nx3271), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_12)) ;
    nor02_2x CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix101 (.Y (
             CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_12), .A0 (
             nx7775), .A1 (nx3273)) ;
    inv01 ix3272 (.Y (nx3273), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_13)) ;
    nor02_2x CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix105 (.Y (
             CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_13), .A0 (
             nx7775), .A1 (nx3275)) ;
    inv01 ix3274 (.Y (nx3275), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_14)) ;
    nor02_2x CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix109 (.Y (
             CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_14), .A0 (
             nx7777), .A1 (nx3277)) ;
    inv01 ix3276 (.Y (nx3277), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_15)) ;
    nor02_2x CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix113 (.Y (
             CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_15), .A0 (
             nx7777), .A1 (nx3279)) ;
    inv01 ix3278 (.Y (nx3279), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_16)) ;
    nor02_2x CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix117 (.Y (
             CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_16), .A0 (
             nx7777), .A1 (nx3279)) ;
    mux21 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix189 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothOperand_0), .A0 (nx3281), .A1 (
          nx3283), .S0 (nx7765)) ;
    inv01 ix3280 (.Y (nx3281), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_0)) ;
    inv01 ix3282 (.Y (nx3283), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_0)) ;
    mux21 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix197 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothOperand_1), .A0 (nx3285), .A1 (
          nx3287), .S0 (nx7765)) ;
    inv01 ix3284 (.Y (nx3285), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_1)) ;
    inv01 ix3286 (.Y (nx3287), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_1)) ;
    mux21 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix205 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothOperand_2), .A0 (nx3289), .A1 (
          nx3291), .S0 (nx7765)) ;
    inv01 ix3288 (.Y (nx3289), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_2)) ;
    inv01 ix3290 (.Y (nx3291), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_2)) ;
    mux21 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix213 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothOperand_3), .A0 (nx3293), .A1 (
          nx3295), .S0 (nx7765)) ;
    inv01 ix3292 (.Y (nx3293), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_3)) ;
    inv01 ix3294 (.Y (nx3295), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_3)) ;
    mux21 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix221 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothOperand_4), .A0 (nx3297), .A1 (
          nx3299), .S0 (nx7765)) ;
    inv01 ix3296 (.Y (nx3297), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_4)) ;
    inv01 ix3298 (.Y (nx3299), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_4)) ;
    mux21 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix229 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothOperand_5), .A0 (nx3301), .A1 (
          nx3303), .S0 (nx7767)) ;
    inv01 ix3300 (.Y (nx3301), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_5)) ;
    inv01 ix3302 (.Y (nx3303), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_5)) ;
    mux21 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix237 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothOperand_6), .A0 (nx3305), .A1 (
          nx3307), .S0 (nx7767)) ;
    inv01 ix3304 (.Y (nx3305), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_6)) ;
    inv01 ix3306 (.Y (nx3307), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_6)) ;
    mux21 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix245 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothOperand_7), .A0 (nx3309), .A1 (
          nx3311), .S0 (nx7767)) ;
    inv01 ix3308 (.Y (nx3309), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_7)) ;
    inv01 ix3310 (.Y (nx3311), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_7)) ;
    mux21 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix253 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothOperand_8), .A0 (nx3313), .A1 (
          nx3315), .S0 (nx7767)) ;
    inv01 ix3312 (.Y (nx3313), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_8)) ;
    inv01 ix3314 (.Y (nx3315), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_8)) ;
    mux21 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix261 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothOperand_9), .A0 (nx3317), .A1 (
          nx3319), .S0 (nx7767)) ;
    inv01 ix3316 (.Y (nx3317), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_9)) ;
    inv01 ix3318 (.Y (nx3319), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_9)) ;
    mux21 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix269 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothOperand_10), .A0 (nx3321), .A1 (
          nx3323), .S0 (nx7767)) ;
    inv01 ix3320 (.Y (nx3321), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_10)) ;
    inv01 ix3322 (.Y (nx3323), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_10)) ;
    mux21 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix277 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothOperand_11), .A0 (nx3325), .A1 (
          nx3327), .S0 (nx7767)) ;
    inv01 ix3324 (.Y (nx3325), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_11)) ;
    inv01 ix3326 (.Y (nx3327), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_11)) ;
    mux21 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix285 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothOperand_12), .A0 (nx3329), .A1 (
          nx3331), .S0 (nx7769)) ;
    inv01 ix3328 (.Y (nx3329), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_12)) ;
    inv01 ix3330 (.Y (nx3331), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_12)) ;
    mux21 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix293 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothOperand_13), .A0 (nx3333), .A1 (
          nx3335), .S0 (nx7769)) ;
    inv01 ix3332 (.Y (nx3333), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_13)) ;
    inv01 ix3334 (.Y (nx3335), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_13)) ;
    mux21 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix301 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothOperand_14), .A0 (nx3337), .A1 (
          nx3339), .S0 (nx7769)) ;
    inv01 ix3336 (.Y (nx3337), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_14)) ;
    inv01 ix3338 (.Y (nx3339), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_14)) ;
    mux21 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix309 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothOperand_15), .A0 (nx3341), .A1 (
          nx3343), .S0 (nx7769)) ;
    inv01 ix3340 (.Y (nx3341), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_15)) ;
    inv01 ix3342 (.Y (nx3343), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_15)) ;
    mux21 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix317 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BoothOperand_16), .A0 (nx3345), .A1 (
          nx3347), .S0 (nx7769)) ;
    inv01 ix3344 (.Y (nx3345), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_16)) ;
    inv01 ix3346 (.Y (nx3347), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_16)) ;
    xnor2 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix321 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_AddPToBoothOperand), .A0 (nx7769), .A1 (
          nx3213)) ;
    oai32 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix393 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .A0 (
          nx8539), .A1 (RST), .A2 (nx7779), .B0 (nx3283), .B1 (nx3351)) ;
    oai32 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix403 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .A0 (
          nx8539), .A1 (RST), .A2 (nx7779), .B0 (nx3287), .B1 (nx3351)) ;
    oai32 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix413 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .A0 (
          nx8539), .A1 (RST), .A2 (nx7779), .B0 (nx3291), .B1 (nx3351)) ;
    oai32 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix423 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .A0 (
          nx8539), .A1 (RST), .A2 (nx7779), .B0 (nx3295), .B1 (nx3351)) ;
    oai32 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix433 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .A0 (
          nx8539), .A1 (RST), .A2 (nx7779), .B0 (nx3299), .B1 (nx3351)) ;
    oai32 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix443 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .A0 (
          nx8539), .A1 (RST), .A2 (nx7779), .B0 (nx3303), .B1 (nx3351)) ;
    oai32 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix453 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .A0 (
          nx8539), .A1 (RST), .A2 (nx7781), .B0 (nx3307), .B1 (nx3351)) ;
    oai32 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix463 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .A0 (
          nx8541), .A1 (RST), .A2 (nx7781), .B0 (nx3311), .B1 (nx3353)) ;
    oai32 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix473 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .A0 (
          nx8541), .A1 (RST), .A2 (nx7781), .B0 (nx3315), .B1 (nx3353)) ;
    oai32 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix483 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .A0 (
          nx3355), .A1 (RST), .A2 (nx7781), .B0 (nx3319), .B1 (nx3353)) ;
    inv01 ix3354 (.Y (nx3355), .A (CacheFilter_2__0__0)) ;
    oai32 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix493 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .A0 (
          nx3357), .A1 (RST), .A2 (nx7781), .B0 (nx3323), .B1 (nx3353)) ;
    inv01 ix3356 (.Y (nx3357), .A (CacheFilter_2__0__1)) ;
    oai32 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix503 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .A0 (
          nx3359), .A1 (RST), .A2 (nx7781), .B0 (nx3327), .B1 (nx3353)) ;
    inv01 ix3358 (.Y (nx3359), .A (CacheFilter_2__0__2)) ;
    oai32 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix513 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .A0 (
          nx3361), .A1 (RST), .A2 (nx7781), .B0 (nx3331), .B1 (nx3353)) ;
    inv01 ix3360 (.Y (nx3361), .A (CacheFilter_2__0__3)) ;
    oai32 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix523 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .A0 (
          nx3363), .A1 (RST), .A2 (nx7783), .B0 (nx3335), .B1 (nx3353)) ;
    inv01 ix3362 (.Y (nx3363), .A (CacheFilter_2__0__4)) ;
    oai32 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix533 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .A0 (
          nx3365), .A1 (RST), .A2 (nx7783), .B0 (nx3339), .B1 (nx3367)) ;
    inv01 ix3364 (.Y (nx3365), .A (CacheFilter_2__0__5)) ;
    inv01 ix3366 (.Y (nx3367), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566)) ;
    oai32 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix543 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .A0 (
          nx3369), .A1 (RST), .A2 (nx7783), .B0 (nx3343), .B1 (nx3367)) ;
    inv01 ix3368 (.Y (nx3369), .A (CacheFilter_2__0__6)) ;
    oai32 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix553 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .A0 (
          nx3371), .A1 (RST), .A2 (nx7783), .B0 (nx3347), .B1 (nx3367)) ;
    inv01 ix3370 (.Y (nx3371), .A (CacheFilter_2__0__7)) ;
    nand02_2x CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix633 (.Y (
              nx3351), .A0 (nx7353), .A1 (nx7783)) ;
    nand02_2x CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix635 (.Y (
              nx3353), .A0 (nx7353), .A1 (nx7783)) ;
    oai32 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix393 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .A0 (
          nx8541), .A1 (RST), .A2 (nx7785), .B0 (nx3281), .B1 (nx3373)) ;
    oai32 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix403 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .A0 (
          nx8541), .A1 (RST), .A2 (nx7785), .B0 (nx3285), .B1 (nx3373)) ;
    oai32 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix413 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .A0 (
          nx8541), .A1 (RST), .A2 (nx7785), .B0 (nx3289), .B1 (nx3373)) ;
    oai32 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix423 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .A0 (
          nx8541), .A1 (RST), .A2 (nx7785), .B0 (nx3293), .B1 (nx3373)) ;
    oai32 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix433 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .A0 (
          nx8541), .A1 (RST), .A2 (nx7785), .B0 (nx3297), .B1 (nx3373)) ;
    oai32 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix443 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .A0 (
          nx8543), .A1 (RST), .A2 (nx7785), .B0 (nx3301), .B1 (nx3373)) ;
    oai32 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix453 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .A0 (
          nx8543), .A1 (RST), .A2 (nx7787), .B0 (nx3305), .B1 (nx3373)) ;
    oai32 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix463 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .A0 (
          nx8543), .A1 (RST), .A2 (nx7787), .B0 (nx3309), .B1 (nx3375)) ;
    oai32 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix473 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .A0 (
          nx8543), .A1 (RST), .A2 (nx7787), .B0 (nx3313), .B1 (nx3375)) ;
    oai32 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix483 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .A0 (
          nx3355), .A1 (RST), .A2 (nx7787), .B0 (nx3317), .B1 (nx3375)) ;
    oai32 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix493 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .A0 (
          nx3377), .A1 (RST), .A2 (nx7787), .B0 (nx3321), .B1 (nx3375)) ;
    inv01 ix3376 (.Y (nx3377), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_10)) ;
    oai32 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix503 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .A0 (
          nx3379), .A1 (RST), .A2 (nx7787), .B0 (nx3325), .B1 (nx3375)) ;
    inv01 ix3378 (.Y (nx3379), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_11)) ;
    oai32 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix513 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .A0 (
          nx3381), .A1 (RST), .A2 (nx7787), .B0 (nx3329), .B1 (nx3375)) ;
    inv01 ix3380 (.Y (nx3381), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_12)) ;
    oai32 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix523 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .A0 (
          nx3383), .A1 (RST), .A2 (nx7789), .B0 (nx3333), .B1 (nx3375)) ;
    inv01 ix3382 (.Y (nx3383), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_13)) ;
    oai32 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix533 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .A0 (
          nx3385), .A1 (RST), .A2 (nx7789), .B0 (nx3337), .B1 (nx3387)) ;
    inv01 ix3384 (.Y (nx3385), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_14)) ;
    inv01 ix3386 (.Y (nx3387), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566)) ;
    oai32 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix543 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .A0 (
          nx3389), .A1 (RST), .A2 (nx7789), .B0 (nx3341), .B1 (nx3387)) ;
    inv01 ix3388 (.Y (nx3389), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_15)) ;
    oai32 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix553 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .A0 (
          nx3391), .A1 (RST), .A2 (nx7789), .B0 (nx3345), .B1 (nx3387)) ;
    inv01 ix3390 (.Y (nx3391), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_16)) ;
    nand02_2x CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix633 (.Y (
              nx3373), .A0 (nx7355), .A1 (nx7789)) ;
    nand02_2x CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix635 (.Y (
              nx3375), .A0 (nx7355), .A1 (nx7789)) ;
    oai32 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix393 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .A0 (
          nx3393), .A1 (RST), .A2 (nx7791), .B0 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx384), .B1 (nx3395)) ;
    inv01 ix3392 (.Y (nx3393), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_0)) ;
    oai32 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix403 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .A0 (
          nx3397), .A1 (RST), .A2 (nx7791), .B0 (nx3213), .B1 (nx3395)) ;
    inv01 ix3396 (.Y (nx3397), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_1)) ;
    oai32 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix413 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .A0 (
          nx3399), .A1 (RST), .A2 (nx7791), .B0 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx387), .B1 (nx3395)) ;
    inv01 ix3398 (.Y (nx3399), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_2)) ;
    oai32 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix423 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .A0 (
          nx3401), .A1 (RST), .A2 (nx7791), .B0 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx399), .B1 (nx3395)) ;
    inv01 ix3400 (.Y (nx3401), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_3)) ;
    oai32 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix433 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .A0 (
          nx3403), .A1 (RST), .A2 (nx7791), .B0 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx409), .B1 (nx3395)) ;
    inv01 ix3402 (.Y (nx3403), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_4)) ;
    oai32 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix443 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .A0 (
          nx3405), .A1 (RST), .A2 (nx7791), .B0 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx419), .B1 (nx3395)) ;
    inv01 ix3404 (.Y (nx3405), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_5)) ;
    oai32 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix453 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .A0 (
          nx3407), .A1 (RST), .A2 (nx7791), .B0 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx429), .B1 (nx3395)) ;
    inv01 ix3406 (.Y (nx3407), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_6)) ;
    oai32 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix463 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .A0 (
          nx3409), .A1 (RST), .A2 (nx7793), .B0 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx439), .B1 (nx3411)) ;
    inv01 ix3408 (.Y (nx3409), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_7)) ;
    oai32 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix473 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .A0 (
          nx3413), .A1 (RST), .A2 (nx7793), .B0 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx449), .B1 (nx3411)) ;
    inv01 ix3412 (.Y (nx3413), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_8)) ;
    oai32 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix483 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .A0 (
          nx3415), .A1 (RST), .A2 (nx7793), .B0 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx469), .B1 (nx3411)) ;
    inv01 ix3414 (.Y (nx3415), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_9)) ;
    oai32 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix493 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .A0 (
          nx3417), .A1 (RST), .A2 (nx7793), .B0 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx477), .B1 (nx3411)) ;
    inv01 ix3416 (.Y (nx3417), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_10)) ;
    oai32 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix503 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .A0 (
          nx3419), .A1 (RST), .A2 (nx7793), .B0 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx485), .B1 (nx3411)) ;
    inv01 ix3418 (.Y (nx3419), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_11)) ;
    oai32 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix513 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .A0 (
          nx3421), .A1 (RST), .A2 (nx7793), .B0 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx493), .B1 (nx3411)) ;
    inv01 ix3420 (.Y (nx3421), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_12)) ;
    oai32 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix523 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .A0 (
          nx3423), .A1 (RST), .A2 (nx7793), .B0 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx501), .B1 (nx3411)) ;
    inv01 ix3422 (.Y (nx3423), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_13)) ;
    oai32 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix533 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .A0 (
          nx3425), .A1 (RST), .A2 (nx7795), .B0 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx509), .B1 (nx3427)) ;
    inv01 ix3424 (.Y (nx3425), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_14)) ;
    inv01 ix3426 (.Y (nx3427), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566)) ;
    oai32 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix543 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .A0 (
          nx3429), .A1 (RST), .A2 (nx7795), .B0 (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_nx517), .B1 (nx3427)) ;
    inv01 ix3428 (.Y (nx3429), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_15)) ;
    oai32 CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix553 (.Y (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .A0 (
          nx3431), .A1 (RST), .A2 (nx7795), .B0 (nx3229), .B1 (nx3427)) ;
    inv01 ix3430 (.Y (nx3431), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_16)) ;
    nand02_2x CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix633 (.Y (
              nx3395), .A0 (nx7355), .A1 (nx7795)) ;
    nand02_2x CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix635 (.Y (
              nx3411), .A0 (nx7355), .A1 (nx7795)) ;
    mux21 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix404 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx403), .A0 (nx3433), .A1 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_2), .S0 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx395)) ;
    inv01 ix3432 (.Y (nx3433), .A (CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx391)) ;
    mux21 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix414 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx413), .A0 (nx3435), .A1 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_3), .S0 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx405)) ;
    inv01 ix3434 (.Y (nx3435), .A (CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx403)) ;
    mux21 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix424 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx423), .A0 (nx3437), .A1 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_4), .S0 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx415)) ;
    inv01 ix3436 (.Y (nx3437), .A (CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx413)) ;
    mux21 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix434 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx433), .A0 (nx3439), .A1 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_5), .S0 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx425)) ;
    inv01 ix3438 (.Y (nx3439), .A (CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx423)) ;
    mux21 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix444 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx443), .A0 (nx3441), .A1 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_6), .S0 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx435)) ;
    inv01 ix3440 (.Y (nx3441), .A (CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx433)) ;
    mux21 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix454 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx453), .A0 (nx3443), .A1 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_7), .S0 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx445)) ;
    inv01 ix3442 (.Y (nx3443), .A (CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx443)) ;
    mux21 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix462 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx461), .A0 (nx3445), .A1 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_8), .S0 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx455)) ;
    inv01 ix3444 (.Y (nx3445), .A (CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx453)) ;
    mux21 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix468 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx467), .A0 (nx3447), .A1 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_9), .S0 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx463)) ;
    inv01 ix3446 (.Y (nx3447), .A (CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx461)) ;
    mux21 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix476 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx475), .A0 (nx3449), .A1 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_10), .S0 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx471)) ;
    inv01 ix3448 (.Y (nx3449), .A (CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx467)) ;
    mux21 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix484 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx483), .A0 (nx3451), .A1 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_11), .S0 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx479)) ;
    inv01 ix3450 (.Y (nx3451), .A (CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx475)) ;
    mux21 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix492 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx491), .A0 (nx3453), .A1 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_12), .S0 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx487)) ;
    inv01 ix3452 (.Y (nx3453), .A (CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx483)) ;
    mux21 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix500 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx499), .A0 (nx3455), .A1 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_13), .S0 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx495)) ;
    inv01 ix3454 (.Y (nx3455), .A (CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx491)) ;
    mux21 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix508 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx507), .A0 (nx3457), .A1 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_14), .S0 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx503)) ;
    inv01 ix3456 (.Y (nx3457), .A (CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx499)) ;
    mux21 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix516 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx515), .A0 (nx3459), .A1 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_15), .S0 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx511)) ;
    inv01 ix3458 (.Y (nx3459), .A (CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx507)) ;
    mux21 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix161 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_1), .A0 (nx3461), .A1 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx379), .S0 (nx7799)) ;
    inv01 ix3460 (.Y (nx3461), .A (CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_1)) ;
    mux21 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix181 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_2), .A0 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx387), .A1 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx389), .S0 (nx7799)) ;
    mux21 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix201 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_3), .A0 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx399), .A1 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx401), .S0 (nx7799)) ;
    mux21 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix221 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_4), .A0 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx409), .A1 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx411), .S0 (nx7799)) ;
    mux21 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix241 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_5), .A0 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx419), .A1 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx421), .S0 (nx7799)) ;
    mux21 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix261 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_6), .A0 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx429), .A1 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx431), .S0 (nx7799)) ;
    mux21 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix281 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_7), .A0 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx439), .A1 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx441), .S0 (nx7799)) ;
    mux21 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix301 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_8), .A0 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx449), .A1 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx451), .S0 (nx7801)) ;
    mux21 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix321 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_9), .A0 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx469), .A1 (nx3463), .S0 (nx7801)) ;
    inv01 ix3462 (.Y (nx3463), .A (CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx316)) ;
    mux21 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix341 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_10), .A0 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx477), .A1 (nx3465), .S0 (nx7801)) ;
    inv01 ix3464 (.Y (nx3465), .A (CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx336)) ;
    mux21 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix361 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_11), .A0 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx485), .A1 (nx3467), .S0 (nx7801)) ;
    inv01 ix3466 (.Y (nx3467), .A (CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx356)) ;
    mux21 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix381 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_12), .A0 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx493), .A1 (nx3469), .S0 (nx7801)) ;
    inv01 ix3468 (.Y (nx3469), .A (CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx376)) ;
    mux21 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix401 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_13), .A0 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx501), .A1 (nx3471), .S0 (nx7801)) ;
    inv01 ix3470 (.Y (nx3471), .A (CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx396)) ;
    mux21 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix421 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_14), .A0 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx509), .A1 (nx3473), .S0 (nx7801)) ;
    inv01 ix3472 (.Y (nx3473), .A (CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx416)) ;
    mux21 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix441 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_15), .A0 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx517), .A1 (nx3475), .S0 (nx7803)) ;
    inv01 ix3474 (.Y (nx3475), .A (CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx436)) ;
    mux21 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_ix461 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_16), .A0 (nx3477), 
          .A1 (nx3479), .S0 (nx7803)) ;
    inv01 ix3476 (.Y (nx3477), .A (CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothP_16)
          ) ;
    inv01 ix3478 (.Y (nx3479), .A (CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx456)) ;
    nor02_2x CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix81 (.Y (
             CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx80), .A0 (Instr), .A1 (
             nx7309)) ;
    nor02_2x CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix319 (.Y (
             CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642), .A0 (
             CALCULATOR_Start_dup_1199), .A1 (
             CALCULATOR_CalculatingBooth_dup_1181)) ;
    nor02_2x CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix85 (.Y (
             CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_0), .A0 (
             nx7813), .A1 (nx3481)) ;
    inv01 ix3480 (.Y (nx3481), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_1)) ;
    mux21 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix125 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_1), .A0 (
          nx3483), .A1 (nx3485), .S0 (nx7813)) ;
    inv01 ix3482 (.Y (nx3483), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_2)) ;
    inv01 ix3484 (.Y (nx3485), .A (CacheWindow_2__1__0)) ;
    mux21 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix133 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_2), .A0 (
          nx3487), .A1 (nx3489), .S0 (nx7813)) ;
    inv01 ix3486 (.Y (nx3487), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_3)) ;
    inv01 ix3488 (.Y (nx3489), .A (CacheWindow_2__1__1)) ;
    mux21 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix141 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_3), .A0 (
          nx3491), .A1 (nx3493), .S0 (nx7813)) ;
    inv01 ix3490 (.Y (nx3491), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_4)) ;
    inv01 ix3492 (.Y (nx3493), .A (CacheWindow_2__1__2)) ;
    mux21 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix149 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_4), .A0 (
          nx3495), .A1 (nx3497), .S0 (nx7813)) ;
    inv01 ix3494 (.Y (nx3495), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_5)) ;
    inv01 ix3496 (.Y (nx3497), .A (CacheWindow_2__1__3)) ;
    mux21 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix157 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_5), .A0 (
          nx3499), .A1 (nx3501), .S0 (nx7813)) ;
    inv01 ix3498 (.Y (nx3499), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_6)) ;
    inv01 ix3500 (.Y (nx3501), .A (CacheWindow_2__1__4)) ;
    mux21 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix165 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_6), .A0 (
          nx3503), .A1 (nx3505), .S0 (nx7813)) ;
    inv01 ix3502 (.Y (nx3503), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_7)) ;
    inv01 ix3504 (.Y (nx3505), .A (CacheWindow_2__1__5)) ;
    mux21 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix173 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_7), .A0 (
          nx3507), .A1 (nx3509), .S0 (nx7815)) ;
    inv01 ix3506 (.Y (nx3507), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_8)) ;
    inv01 ix3508 (.Y (nx3509), .A (CacheWindow_2__1__6)) ;
    mux21 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix181 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_8), .A0 (
          nx3511), .A1 (nx3513), .S0 (nx7815)) ;
    inv01 ix3510 (.Y (nx3511), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_9)) ;
    inv01 ix3512 (.Y (nx3513), .A (CacheWindow_2__1__7)) ;
    nor02_2x CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix89 (.Y (
             CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_9), .A0 (
             nx7815), .A1 (nx3515)) ;
    inv01 ix3514 (.Y (nx3515), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_10)) ;
    nor02_2x CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix93 (.Y (
             CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_10), .A0 (
             nx7815), .A1 (nx3517)) ;
    inv01 ix3516 (.Y (nx3517), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_11)) ;
    nor02_2x CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix97 (.Y (
             CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_11), .A0 (
             nx7815), .A1 (nx3519)) ;
    inv01 ix3518 (.Y (nx3519), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_12)) ;
    nor02_2x CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix101 (.Y (
             CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_12), .A0 (
             nx7815), .A1 (nx3521)) ;
    inv01 ix3520 (.Y (nx3521), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_13)) ;
    nor02_2x CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix105 (.Y (
             CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_13), .A0 (
             nx7815), .A1 (nx3523)) ;
    inv01 ix3522 (.Y (nx3523), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_14)) ;
    nor02_2x CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix109 (.Y (
             CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_14), .A0 (
             nx7817), .A1 (nx3525)) ;
    inv01 ix3524 (.Y (nx3525), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_15)) ;
    nor02_2x CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix113 (.Y (
             CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_15), .A0 (
             nx7817), .A1 (nx3527)) ;
    inv01 ix3526 (.Y (nx3527), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_16)) ;
    nor02_2x CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix117 (.Y (
             CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_16), .A0 (
             nx7817), .A1 (nx3527)) ;
    mux21 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix189 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothOperand_0), .A0 (nx3529), .A1 (
          nx3531), .S0 (nx7805)) ;
    inv01 ix3528 (.Y (nx3529), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_0)) ;
    inv01 ix3530 (.Y (nx3531), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_0)) ;
    mux21 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix197 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothOperand_1), .A0 (nx3533), .A1 (
          nx3535), .S0 (nx7805)) ;
    inv01 ix3532 (.Y (nx3533), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_1)) ;
    inv01 ix3534 (.Y (nx3535), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_1)) ;
    mux21 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix205 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothOperand_2), .A0 (nx3537), .A1 (
          nx3539), .S0 (nx7805)) ;
    inv01 ix3536 (.Y (nx3537), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_2)) ;
    inv01 ix3538 (.Y (nx3539), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_2)) ;
    mux21 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix213 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothOperand_3), .A0 (nx3541), .A1 (
          nx3543), .S0 (nx7805)) ;
    inv01 ix3540 (.Y (nx3541), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_3)) ;
    inv01 ix3542 (.Y (nx3543), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_3)) ;
    mux21 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix221 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothOperand_4), .A0 (nx3545), .A1 (
          nx3547), .S0 (nx7805)) ;
    inv01 ix3544 (.Y (nx3545), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_4)) ;
    inv01 ix3546 (.Y (nx3547), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_4)) ;
    mux21 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix229 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothOperand_5), .A0 (nx3549), .A1 (
          nx3551), .S0 (nx7807)) ;
    inv01 ix3548 (.Y (nx3549), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_5)) ;
    inv01 ix3550 (.Y (nx3551), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_5)) ;
    mux21 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix237 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothOperand_6), .A0 (nx3553), .A1 (
          nx3555), .S0 (nx7807)) ;
    inv01 ix3552 (.Y (nx3553), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_6)) ;
    inv01 ix3554 (.Y (nx3555), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_6)) ;
    mux21 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix245 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothOperand_7), .A0 (nx3557), .A1 (
          nx3559), .S0 (nx7807)) ;
    inv01 ix3556 (.Y (nx3557), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_7)) ;
    inv01 ix3558 (.Y (nx3559), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_7)) ;
    mux21 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix253 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothOperand_8), .A0 (nx3561), .A1 (
          nx3563), .S0 (nx7807)) ;
    inv01 ix3560 (.Y (nx3561), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_8)) ;
    inv01 ix3562 (.Y (nx3563), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_8)) ;
    mux21 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix261 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothOperand_9), .A0 (nx3565), .A1 (
          nx3567), .S0 (nx7807)) ;
    inv01 ix3564 (.Y (nx3565), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_9)) ;
    inv01 ix3566 (.Y (nx3567), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_9)) ;
    mux21 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix269 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothOperand_10), .A0 (nx3569), .A1 (
          nx3571), .S0 (nx7807)) ;
    inv01 ix3568 (.Y (nx3569), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_10)) ;
    inv01 ix3570 (.Y (nx3571), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_10)) ;
    mux21 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix277 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothOperand_11), .A0 (nx3573), .A1 (
          nx3575), .S0 (nx7807)) ;
    inv01 ix3572 (.Y (nx3573), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_11)) ;
    inv01 ix3574 (.Y (nx3575), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_11)) ;
    mux21 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix285 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothOperand_12), .A0 (nx3577), .A1 (
          nx3579), .S0 (nx7809)) ;
    inv01 ix3576 (.Y (nx3577), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_12)) ;
    inv01 ix3578 (.Y (nx3579), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_12)) ;
    mux21 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix293 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothOperand_13), .A0 (nx3581), .A1 (
          nx3583), .S0 (nx7809)) ;
    inv01 ix3580 (.Y (nx3581), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_13)) ;
    inv01 ix3582 (.Y (nx3583), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_13)) ;
    mux21 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix301 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothOperand_14), .A0 (nx3585), .A1 (
          nx3587), .S0 (nx7809)) ;
    inv01 ix3584 (.Y (nx3585), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_14)) ;
    inv01 ix3586 (.Y (nx3587), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_14)) ;
    mux21 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix309 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothOperand_15), .A0 (nx3589), .A1 (
          nx3591), .S0 (nx7809)) ;
    inv01 ix3588 (.Y (nx3589), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_15)) ;
    inv01 ix3590 (.Y (nx3591), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_15)) ;
    mux21 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix317 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BoothOperand_16), .A0 (nx3593), .A1 (
          nx3595), .S0 (nx7809)) ;
    inv01 ix3592 (.Y (nx3593), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_16)) ;
    inv01 ix3594 (.Y (nx3595), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_16)) ;
    xnor2 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix321 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_AddPToBoothOperand), .A0 (nx7809), .A1 (
          nx3461)) ;
    oai32 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix393 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .A0 (
          nx8545), .A1 (RST), .A2 (nx7819), .B0 (nx3531), .B1 (nx3599)) ;
    oai32 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix403 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .A0 (
          nx8545), .A1 (RST), .A2 (nx7819), .B0 (nx3535), .B1 (nx3599)) ;
    oai32 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix413 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .A0 (
          nx8545), .A1 (RST), .A2 (nx7819), .B0 (nx3539), .B1 (nx3599)) ;
    oai32 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix423 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .A0 (
          nx8545), .A1 (RST), .A2 (nx7819), .B0 (nx3543), .B1 (nx3599)) ;
    oai32 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix433 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .A0 (
          nx8545), .A1 (RST), .A2 (nx7819), .B0 (nx3547), .B1 (nx3599)) ;
    oai32 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix443 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .A0 (
          nx8545), .A1 (RST), .A2 (nx7819), .B0 (nx3551), .B1 (nx3599)) ;
    oai32 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix453 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .A0 (
          nx8545), .A1 (RST), .A2 (nx7821), .B0 (nx3555), .B1 (nx3599)) ;
    oai32 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix463 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .A0 (
          nx8547), .A1 (RST), .A2 (nx7821), .B0 (nx3559), .B1 (nx3601)) ;
    oai32 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix473 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .A0 (
          nx8547), .A1 (RST), .A2 (nx7821), .B0 (nx3563), .B1 (nx3601)) ;
    oai32 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix483 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .A0 (
          nx3603), .A1 (RST), .A2 (nx7821), .B0 (nx3567), .B1 (nx3601)) ;
    inv01 ix3602 (.Y (nx3603), .A (CacheFilter_2__1__0)) ;
    oai32 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix493 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .A0 (
          nx3605), .A1 (RST), .A2 (nx7821), .B0 (nx3571), .B1 (nx3601)) ;
    inv01 ix3604 (.Y (nx3605), .A (CacheFilter_2__1__1)) ;
    oai32 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix503 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .A0 (
          nx3607), .A1 (RST), .A2 (nx7821), .B0 (nx3575), .B1 (nx3601)) ;
    inv01 ix3606 (.Y (nx3607), .A (CacheFilter_2__1__2)) ;
    oai32 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix513 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .A0 (
          nx3609), .A1 (RST), .A2 (nx7821), .B0 (nx3579), .B1 (nx3601)) ;
    inv01 ix3608 (.Y (nx3609), .A (CacheFilter_2__1__3)) ;
    oai32 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix523 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .A0 (
          nx3611), .A1 (RST), .A2 (nx7823), .B0 (nx3583), .B1 (nx3601)) ;
    inv01 ix3610 (.Y (nx3611), .A (CacheFilter_2__1__4)) ;
    oai32 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix533 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .A0 (
          nx3613), .A1 (RST), .A2 (nx7823), .B0 (nx3587), .B1 (nx3615)) ;
    inv01 ix3612 (.Y (nx3613), .A (CacheFilter_2__1__5)) ;
    inv01 ix3614 (.Y (nx3615), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566)) ;
    oai32 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix543 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .A0 (
          nx3617), .A1 (RST), .A2 (nx7823), .B0 (nx3591), .B1 (nx3615)) ;
    inv01 ix3616 (.Y (nx3617), .A (CacheFilter_2__1__6)) ;
    oai32 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix553 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .A0 (
          nx3619), .A1 (RST), .A2 (nx7823), .B0 (nx3595), .B1 (nx3615)) ;
    inv01 ix3618 (.Y (nx3619), .A (CacheFilter_2__1__7)) ;
    nand02_2x CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix633 (.Y (
              nx3599), .A0 (nx7355), .A1 (nx7823)) ;
    nand02_2x CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix635 (.Y (
              nx3601), .A0 (nx7355), .A1 (nx7823)) ;
    oai32 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix393 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .A0 (
          nx8547), .A1 (RST), .A2 (nx7825), .B0 (nx3529), .B1 (nx3621)) ;
    oai32 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix403 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .A0 (
          nx8547), .A1 (RST), .A2 (nx7825), .B0 (nx3533), .B1 (nx3621)) ;
    oai32 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix413 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .A0 (
          nx8547), .A1 (RST), .A2 (nx7825), .B0 (nx3537), .B1 (nx3621)) ;
    oai32 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix423 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .A0 (
          nx8547), .A1 (RST), .A2 (nx7825), .B0 (nx3541), .B1 (nx3621)) ;
    oai32 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix433 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .A0 (
          nx8547), .A1 (RST), .A2 (nx7825), .B0 (nx3545), .B1 (nx3621)) ;
    oai32 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix443 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .A0 (
          nx8549), .A1 (RST), .A2 (nx7825), .B0 (nx3549), .B1 (nx3621)) ;
    oai32 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix453 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .A0 (
          nx8549), .A1 (RST), .A2 (nx7827), .B0 (nx3553), .B1 (nx3621)) ;
    oai32 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix463 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .A0 (
          nx8549), .A1 (RST), .A2 (nx7827), .B0 (nx3557), .B1 (nx3623)) ;
    oai32 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix473 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .A0 (
          nx8549), .A1 (RST), .A2 (nx7827), .B0 (nx3561), .B1 (nx3623)) ;
    oai32 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix483 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .A0 (
          nx3603), .A1 (RST), .A2 (nx7827), .B0 (nx3565), .B1 (nx3623)) ;
    oai32 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix493 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .A0 (
          nx3625), .A1 (RST), .A2 (nx7827), .B0 (nx3569), .B1 (nx3623)) ;
    inv01 ix3624 (.Y (nx3625), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_10)) ;
    oai32 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix503 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .A0 (
          nx3627), .A1 (RST), .A2 (nx7827), .B0 (nx3573), .B1 (nx3623)) ;
    inv01 ix3626 (.Y (nx3627), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_11)) ;
    oai32 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix513 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .A0 (
          nx3629), .A1 (RST), .A2 (nx7827), .B0 (nx3577), .B1 (nx3623)) ;
    inv01 ix3628 (.Y (nx3629), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_12)) ;
    oai32 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix523 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .A0 (
          nx3631), .A1 (RST), .A2 (nx7829), .B0 (nx3581), .B1 (nx3623)) ;
    inv01 ix3630 (.Y (nx3631), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_13)) ;
    oai32 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix533 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .A0 (
          nx3633), .A1 (RST), .A2 (nx7829), .B0 (nx3585), .B1 (nx3635)) ;
    inv01 ix3632 (.Y (nx3633), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_14)) ;
    inv01 ix3634 (.Y (nx3635), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566)) ;
    oai32 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix543 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .A0 (
          nx3637), .A1 (RST), .A2 (nx7829), .B0 (nx3589), .B1 (nx3635)) ;
    inv01 ix3636 (.Y (nx3637), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_15)) ;
    oai32 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix553 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .A0 (
          nx3639), .A1 (RST), .A2 (nx7829), .B0 (nx3593), .B1 (nx3635)) ;
    inv01 ix3638 (.Y (nx3639), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_16)) ;
    nand02_2x CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix633 (.Y (
              nx3621), .A0 (nx7355), .A1 (nx7829)) ;
    nand02_2x CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix635 (.Y (
              nx3623), .A0 (nx7357), .A1 (nx7829)) ;
    oai32 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix393 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .A0 (
          nx3641), .A1 (RST), .A2 (nx7831), .B0 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx384), .B1 (nx3643)) ;
    inv01 ix3640 (.Y (nx3641), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_0)) ;
    oai32 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix403 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .A0 (
          nx3645), .A1 (RST), .A2 (nx7831), .B0 (nx3461), .B1 (nx3643)) ;
    inv01 ix3644 (.Y (nx3645), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_1)) ;
    oai32 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix413 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .A0 (
          nx3647), .A1 (RST), .A2 (nx7831), .B0 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx387), .B1 (nx3643)) ;
    inv01 ix3646 (.Y (nx3647), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_2)) ;
    oai32 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix423 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .A0 (
          nx3649), .A1 (RST), .A2 (nx7831), .B0 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx399), .B1 (nx3643)) ;
    inv01 ix3648 (.Y (nx3649), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_3)) ;
    oai32 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix433 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .A0 (
          nx3651), .A1 (RST), .A2 (nx7831), .B0 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx409), .B1 (nx3643)) ;
    inv01 ix3650 (.Y (nx3651), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_4)) ;
    oai32 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix443 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .A0 (
          nx3653), .A1 (RST), .A2 (nx7831), .B0 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx419), .B1 (nx3643)) ;
    inv01 ix3652 (.Y (nx3653), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_5)) ;
    oai32 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix453 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .A0 (
          nx3655), .A1 (RST), .A2 (nx7831), .B0 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx429), .B1 (nx3643)) ;
    inv01 ix3654 (.Y (nx3655), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_6)) ;
    oai32 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix463 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .A0 (
          nx3657), .A1 (RST), .A2 (nx7833), .B0 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx439), .B1 (nx3659)) ;
    inv01 ix3656 (.Y (nx3657), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_7)) ;
    oai32 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix473 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .A0 (
          nx3661), .A1 (RST), .A2 (nx7833), .B0 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx449), .B1 (nx3659)) ;
    inv01 ix3660 (.Y (nx3661), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_8)) ;
    oai32 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix483 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .A0 (
          nx3663), .A1 (RST), .A2 (nx7833), .B0 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx469), .B1 (nx3659)) ;
    inv01 ix3662 (.Y (nx3663), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_9)) ;
    oai32 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix493 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .A0 (
          nx3665), .A1 (RST), .A2 (nx7833), .B0 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx477), .B1 (nx3659)) ;
    inv01 ix3664 (.Y (nx3665), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_10)) ;
    oai32 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix503 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .A0 (
          nx3667), .A1 (RST), .A2 (nx7833), .B0 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx485), .B1 (nx3659)) ;
    inv01 ix3666 (.Y (nx3667), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_11)) ;
    oai32 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix513 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .A0 (
          nx3669), .A1 (RST), .A2 (nx7833), .B0 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx493), .B1 (nx3659)) ;
    inv01 ix3668 (.Y (nx3669), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_12)) ;
    oai32 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix523 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .A0 (
          nx3671), .A1 (RST), .A2 (nx7833), .B0 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx501), .B1 (nx3659)) ;
    inv01 ix3670 (.Y (nx3671), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_13)) ;
    oai32 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix533 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .A0 (
          nx3673), .A1 (RST), .A2 (nx7835), .B0 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx509), .B1 (nx3675)) ;
    inv01 ix3672 (.Y (nx3673), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_14)) ;
    inv01 ix3674 (.Y (nx3675), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566)) ;
    oai32 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix543 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .A0 (
          nx3677), .A1 (RST), .A2 (nx7835), .B0 (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_nx517), .B1 (nx3675)) ;
    inv01 ix3676 (.Y (nx3677), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_15)) ;
    oai32 CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix553 (.Y (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .A0 (
          nx3679), .A1 (RST), .A2 (nx7835), .B0 (nx3477), .B1 (nx3675)) ;
    inv01 ix3678 (.Y (nx3679), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_16)) ;
    nand02_2x CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix633 (.Y (
              nx3643), .A0 (nx7357), .A1 (nx7835)) ;
    nand02_2x CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix635 (.Y (
              nx3659), .A0 (nx7357), .A1 (nx7835)) ;
    mux21 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix404 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx403), .A0 (nx3681), .A1 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_2), .S0 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx395)) ;
    inv01 ix3680 (.Y (nx3681), .A (CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx391)) ;
    mux21 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix414 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx413), .A0 (nx3683), .A1 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_3), .S0 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx405)) ;
    inv01 ix3682 (.Y (nx3683), .A (CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx403)) ;
    mux21 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix424 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx423), .A0 (nx3685), .A1 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_4), .S0 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx415)) ;
    inv01 ix3684 (.Y (nx3685), .A (CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx413)) ;
    mux21 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix434 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx433), .A0 (nx3687), .A1 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_5), .S0 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx425)) ;
    inv01 ix3686 (.Y (nx3687), .A (CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx423)) ;
    mux21 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix444 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx443), .A0 (nx3689), .A1 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_6), .S0 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx435)) ;
    inv01 ix3688 (.Y (nx3689), .A (CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx433)) ;
    mux21 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix454 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx453), .A0 (nx3691), .A1 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_7), .S0 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx445)) ;
    inv01 ix3690 (.Y (nx3691), .A (CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx443)) ;
    mux21 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix462 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx461), .A0 (nx3693), .A1 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_8), .S0 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx455)) ;
    inv01 ix3692 (.Y (nx3693), .A (CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx453)) ;
    mux21 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix468 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx467), .A0 (nx3695), .A1 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_9), .S0 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx463)) ;
    inv01 ix3694 (.Y (nx3695), .A (CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx461)) ;
    mux21 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix476 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx475), .A0 (nx3697), .A1 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_10), .S0 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx471)) ;
    inv01 ix3696 (.Y (nx3697), .A (CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx467)) ;
    mux21 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix484 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx483), .A0 (nx3699), .A1 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_11), .S0 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx479)) ;
    inv01 ix3698 (.Y (nx3699), .A (CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx475)) ;
    mux21 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix492 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx491), .A0 (nx3701), .A1 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_12), .S0 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx487)) ;
    inv01 ix3700 (.Y (nx3701), .A (CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx483)) ;
    mux21 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix500 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx499), .A0 (nx3703), .A1 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_13), .S0 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx495)) ;
    inv01 ix3702 (.Y (nx3703), .A (CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx491)) ;
    mux21 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix508 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx507), .A0 (nx3705), .A1 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_14), .S0 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx503)) ;
    inv01 ix3704 (.Y (nx3705), .A (CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx499)) ;
    mux21 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix516 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx515), .A0 (nx3707), .A1 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_15), .S0 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx511)) ;
    inv01 ix3706 (.Y (nx3707), .A (CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx507)) ;
    mux21 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix161 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_1), .A0 (nx3709), .A1 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx379), .S0 (nx7839)) ;
    inv01 ix3708 (.Y (nx3709), .A (CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_1)) ;
    mux21 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix181 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_2), .A0 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx387), .A1 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx389), .S0 (nx7839)) ;
    mux21 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix201 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_3), .A0 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx399), .A1 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx401), .S0 (nx7839)) ;
    mux21 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix221 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_4), .A0 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx409), .A1 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx411), .S0 (nx7839)) ;
    mux21 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix241 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_5), .A0 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx419), .A1 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx421), .S0 (nx7839)) ;
    mux21 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix261 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_6), .A0 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx429), .A1 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx431), .S0 (nx7839)) ;
    mux21 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix281 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_7), .A0 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx439), .A1 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx441), .S0 (nx7839)) ;
    mux21 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix301 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_8), .A0 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx449), .A1 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx451), .S0 (nx7841)) ;
    mux21 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix321 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_9), .A0 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx469), .A1 (nx3711), .S0 (nx7841)) ;
    inv01 ix3710 (.Y (nx3711), .A (CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx316)) ;
    mux21 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix341 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_10), .A0 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx477), .A1 (nx3713), .S0 (nx7841)) ;
    inv01 ix3712 (.Y (nx3713), .A (CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx336)) ;
    mux21 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix361 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_11), .A0 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx485), .A1 (nx3715), .S0 (nx7841)) ;
    inv01 ix3714 (.Y (nx3715), .A (CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx356)) ;
    mux21 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix381 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_12), .A0 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx493), .A1 (nx3717), .S0 (nx7841)) ;
    inv01 ix3716 (.Y (nx3717), .A (CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx376)) ;
    mux21 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix401 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_13), .A0 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx501), .A1 (nx3719), .S0 (nx7841)) ;
    inv01 ix3718 (.Y (nx3719), .A (CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx396)) ;
    mux21 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix421 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_14), .A0 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx509), .A1 (nx3721), .S0 (nx7841)) ;
    inv01 ix3720 (.Y (nx3721), .A (CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx416)) ;
    mux21 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix441 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_15), .A0 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx517), .A1 (nx3723), .S0 (nx7843)) ;
    inv01 ix3722 (.Y (nx3723), .A (CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx436)) ;
    mux21 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_ix461 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_16), .A0 (nx3725), 
          .A1 (nx3727), .S0 (nx7843)) ;
    inv01 ix3724 (.Y (nx3725), .A (CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothP_16)
          ) ;
    inv01 ix3726 (.Y (nx3727), .A (CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx456)) ;
    nor02_2x CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix81 (.Y (
             CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx80), .A0 (Instr), .A1 (
             nx7309)) ;
    nor02_2x CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix319 (.Y (
             CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642), .A0 (
             CALCULATOR_Start_dup_1204), .A1 (
             CALCULATOR_CalculatingBooth_dup_1181)) ;
    nor02_2x CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix85 (.Y (
             CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_0), .A0 (
             nx7853), .A1 (nx3729)) ;
    inv01 ix3728 (.Y (nx3729), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_1)) ;
    mux21 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix125 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_1), .A0 (
          nx3731), .A1 (nx3733), .S0 (nx7853)) ;
    inv01 ix3730 (.Y (nx3731), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_2)) ;
    inv01 ix3732 (.Y (nx3733), .A (CacheWindow_2__2__0)) ;
    mux21 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix133 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_2), .A0 (
          nx3735), .A1 (nx3737), .S0 (nx7853)) ;
    inv01 ix3734 (.Y (nx3735), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_3)) ;
    inv01 ix3736 (.Y (nx3737), .A (CacheWindow_2__2__1)) ;
    mux21 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix141 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_3), .A0 (
          nx3739), .A1 (nx3741), .S0 (nx7853)) ;
    inv01 ix3738 (.Y (nx3739), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_4)) ;
    inv01 ix3740 (.Y (nx3741), .A (CacheWindow_2__2__2)) ;
    mux21 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix149 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_4), .A0 (
          nx3743), .A1 (nx3745), .S0 (nx7853)) ;
    inv01 ix3742 (.Y (nx3743), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_5)) ;
    inv01 ix3744 (.Y (nx3745), .A (CacheWindow_2__2__3)) ;
    mux21 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix157 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_5), .A0 (
          nx3747), .A1 (nx3749), .S0 (nx7853)) ;
    inv01 ix3746 (.Y (nx3747), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_6)) ;
    inv01 ix3748 (.Y (nx3749), .A (CacheWindow_2__2__4)) ;
    mux21 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix165 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_6), .A0 (
          nx3751), .A1 (nx3753), .S0 (nx7853)) ;
    inv01 ix3750 (.Y (nx3751), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_7)) ;
    inv01 ix3752 (.Y (nx3753), .A (CacheWindow_2__2__5)) ;
    mux21 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix173 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_7), .A0 (
          nx3755), .A1 (nx3757), .S0 (nx7855)) ;
    inv01 ix3754 (.Y (nx3755), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_8)) ;
    inv01 ix3756 (.Y (nx3757), .A (CacheWindow_2__2__6)) ;
    mux21 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix181 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_8), .A0 (
          nx3759), .A1 (nx3761), .S0 (nx7855)) ;
    inv01 ix3758 (.Y (nx3759), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_9)) ;
    inv01 ix3760 (.Y (nx3761), .A (CacheWindow_2__2__7)) ;
    nor02_2x CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix89 (.Y (
             CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_9), .A0 (
             nx7855), .A1 (nx3763)) ;
    inv01 ix3762 (.Y (nx3763), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_10)) ;
    nor02_2x CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix93 (.Y (
             CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_10), .A0 (
             nx7855), .A1 (nx3765)) ;
    inv01 ix3764 (.Y (nx3765), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_11)) ;
    nor02_2x CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix97 (.Y (
             CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_11), .A0 (
             nx7855), .A1 (nx3767)) ;
    inv01 ix3766 (.Y (nx3767), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_12)) ;
    nor02_2x CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix101 (.Y (
             CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_12), .A0 (
             nx7855), .A1 (nx3769)) ;
    inv01 ix3768 (.Y (nx3769), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_13)) ;
    nor02_2x CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix105 (.Y (
             CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_13), .A0 (
             nx7855), .A1 (nx3771)) ;
    inv01 ix3770 (.Y (nx3771), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_14)) ;
    nor02_2x CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix109 (.Y (
             CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_14), .A0 (
             nx7857), .A1 (nx3773)) ;
    inv01 ix3772 (.Y (nx3773), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_15)) ;
    nor02_2x CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix113 (.Y (
             CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_15), .A0 (
             nx7857), .A1 (nx3775)) ;
    inv01 ix3774 (.Y (nx3775), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_16)) ;
    nor02_2x CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix117 (.Y (
             CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_16), .A0 (
             nx7857), .A1 (nx3775)) ;
    mux21 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix189 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothOperand_0), .A0 (nx3777), .A1 (
          nx3779), .S0 (nx7845)) ;
    inv01 ix3776 (.Y (nx3777), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_0)) ;
    inv01 ix3778 (.Y (nx3779), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_0)) ;
    mux21 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix197 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothOperand_1), .A0 (nx3781), .A1 (
          nx3783), .S0 (nx7845)) ;
    inv01 ix3780 (.Y (nx3781), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_1)) ;
    inv01 ix3782 (.Y (nx3783), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_1)) ;
    mux21 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix205 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothOperand_2), .A0 (nx3785), .A1 (
          nx3787), .S0 (nx7845)) ;
    inv01 ix3784 (.Y (nx3785), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_2)) ;
    inv01 ix3786 (.Y (nx3787), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_2)) ;
    mux21 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix213 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothOperand_3), .A0 (nx3789), .A1 (
          nx3791), .S0 (nx7845)) ;
    inv01 ix3788 (.Y (nx3789), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_3)) ;
    inv01 ix3790 (.Y (nx3791), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_3)) ;
    mux21 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix221 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothOperand_4), .A0 (nx3793), .A1 (
          nx3795), .S0 (nx7845)) ;
    inv01 ix3792 (.Y (nx3793), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_4)) ;
    inv01 ix3794 (.Y (nx3795), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_4)) ;
    mux21 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix229 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothOperand_5), .A0 (nx3797), .A1 (
          nx3799), .S0 (nx7847)) ;
    inv01 ix3796 (.Y (nx3797), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_5)) ;
    inv01 ix3798 (.Y (nx3799), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_5)) ;
    mux21 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix237 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothOperand_6), .A0 (nx3801), .A1 (
          nx3803), .S0 (nx7847)) ;
    inv01 ix3800 (.Y (nx3801), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_6)) ;
    inv01 ix3802 (.Y (nx3803), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_6)) ;
    mux21 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix245 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothOperand_7), .A0 (nx3805), .A1 (
          nx3807), .S0 (nx7847)) ;
    inv01 ix3804 (.Y (nx3805), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_7)) ;
    inv01 ix3806 (.Y (nx3807), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_7)) ;
    mux21 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix253 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothOperand_8), .A0 (nx3809), .A1 (
          nx3811), .S0 (nx7847)) ;
    inv01 ix3808 (.Y (nx3809), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_8)) ;
    inv01 ix3810 (.Y (nx3811), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_8)) ;
    mux21 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix261 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothOperand_9), .A0 (nx3813), .A1 (
          nx3815), .S0 (nx7847)) ;
    inv01 ix3812 (.Y (nx3813), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_9)) ;
    inv01 ix3814 (.Y (nx3815), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_9)) ;
    mux21 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix269 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothOperand_10), .A0 (nx3817), .A1 (
          nx3819), .S0 (nx7847)) ;
    inv01 ix3816 (.Y (nx3817), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_10)) ;
    inv01 ix3818 (.Y (nx3819), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_10)) ;
    mux21 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix277 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothOperand_11), .A0 (nx3821), .A1 (
          nx3823), .S0 (nx7847)) ;
    inv01 ix3820 (.Y (nx3821), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_11)) ;
    inv01 ix3822 (.Y (nx3823), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_11)) ;
    mux21 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix285 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothOperand_12), .A0 (nx3825), .A1 (
          nx3827), .S0 (nx7849)) ;
    inv01 ix3824 (.Y (nx3825), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_12)) ;
    inv01 ix3826 (.Y (nx3827), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_12)) ;
    mux21 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix293 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothOperand_13), .A0 (nx3829), .A1 (
          nx3831), .S0 (nx7849)) ;
    inv01 ix3828 (.Y (nx3829), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_13)) ;
    inv01 ix3830 (.Y (nx3831), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_13)) ;
    mux21 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix301 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothOperand_14), .A0 (nx3833), .A1 (
          nx3835), .S0 (nx7849)) ;
    inv01 ix3832 (.Y (nx3833), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_14)) ;
    inv01 ix3834 (.Y (nx3835), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_14)) ;
    mux21 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix309 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothOperand_15), .A0 (nx3837), .A1 (
          nx3839), .S0 (nx7849)) ;
    inv01 ix3836 (.Y (nx3837), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_15)) ;
    inv01 ix3838 (.Y (nx3839), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_15)) ;
    mux21 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix317 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BoothOperand_16), .A0 (nx3841), .A1 (
          nx3843), .S0 (nx7849)) ;
    inv01 ix3840 (.Y (nx3841), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_16)) ;
    inv01 ix3842 (.Y (nx3843), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_16)) ;
    xnor2 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix321 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_AddPToBoothOperand), .A0 (nx7849), .A1 (
          nx3709)) ;
    oai32 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix393 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .A0 (
          nx8551), .A1 (RST), .A2 (nx7859), .B0 (nx3779), .B1 (nx3847)) ;
    oai32 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix403 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .A0 (
          nx8551), .A1 (RST), .A2 (nx7859), .B0 (nx3783), .B1 (nx3847)) ;
    oai32 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix413 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .A0 (
          nx8551), .A1 (RST), .A2 (nx7859), .B0 (nx3787), .B1 (nx3847)) ;
    oai32 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix423 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .A0 (
          nx8551), .A1 (RST), .A2 (nx7859), .B0 (nx3791), .B1 (nx3847)) ;
    oai32 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix433 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .A0 (
          nx8551), .A1 (RST), .A2 (nx7859), .B0 (nx3795), .B1 (nx3847)) ;
    oai32 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix443 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .A0 (
          nx8551), .A1 (RST), .A2 (nx7859), .B0 (nx3799), .B1 (nx3847)) ;
    oai32 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix453 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .A0 (
          nx8551), .A1 (RST), .A2 (nx7861), .B0 (nx3803), .B1 (nx3847)) ;
    oai32 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix463 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .A0 (
          nx8553), .A1 (RST), .A2 (nx7861), .B0 (nx3807), .B1 (nx3849)) ;
    oai32 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix473 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .A0 (
          nx8553), .A1 (RST), .A2 (nx7861), .B0 (nx3811), .B1 (nx3849)) ;
    oai32 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix483 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .A0 (
          nx3851), .A1 (RST), .A2 (nx7861), .B0 (nx3815), .B1 (nx3849)) ;
    inv01 ix3850 (.Y (nx3851), .A (CacheFilter_2__2__0)) ;
    oai32 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix493 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .A0 (
          nx3853), .A1 (RST), .A2 (nx7861), .B0 (nx3819), .B1 (nx3849)) ;
    inv01 ix3852 (.Y (nx3853), .A (CacheFilter_2__2__1)) ;
    oai32 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix503 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .A0 (
          nx3855), .A1 (RST), .A2 (nx7861), .B0 (nx3823), .B1 (nx3849)) ;
    inv01 ix3854 (.Y (nx3855), .A (CacheFilter_2__2__2)) ;
    oai32 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix513 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .A0 (
          nx3857), .A1 (RST), .A2 (nx7861), .B0 (nx3827), .B1 (nx3849)) ;
    inv01 ix3856 (.Y (nx3857), .A (CacheFilter_2__2__3)) ;
    oai32 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix523 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .A0 (
          nx3859), .A1 (RST), .A2 (nx7863), .B0 (nx3831), .B1 (nx3849)) ;
    inv01 ix3858 (.Y (nx3859), .A (CacheFilter_2__2__4)) ;
    oai32 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix533 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .A0 (
          nx3861), .A1 (RST), .A2 (nx7863), .B0 (nx3835), .B1 (nx3863)) ;
    inv01 ix3860 (.Y (nx3861), .A (CacheFilter_2__2__5)) ;
    inv01 ix3862 (.Y (nx3863), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566)) ;
    oai32 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix543 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .A0 (
          nx3865), .A1 (RST), .A2 (nx7863), .B0 (nx3839), .B1 (nx3863)) ;
    inv01 ix3864 (.Y (nx3865), .A (CacheFilter_2__2__6)) ;
    oai32 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix553 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .A0 (
          nx3867), .A1 (RST), .A2 (nx7863), .B0 (nx3843), .B1 (nx3863)) ;
    inv01 ix3866 (.Y (nx3867), .A (CacheFilter_2__2__7)) ;
    nand02_2x CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix633 (.Y (
              nx3847), .A0 (nx7357), .A1 (nx7863)) ;
    nand02_2x CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix635 (.Y (
              nx3849), .A0 (nx7357), .A1 (nx7863)) ;
    oai32 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix393 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .A0 (
          nx8553), .A1 (RST), .A2 (nx7865), .B0 (nx3777), .B1 (nx3869)) ;
    oai32 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix403 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .A0 (
          nx8553), .A1 (RST), .A2 (nx7865), .B0 (nx3781), .B1 (nx3869)) ;
    oai32 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix413 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .A0 (
          nx8553), .A1 (RST), .A2 (nx7865), .B0 (nx3785), .B1 (nx3869)) ;
    oai32 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix423 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .A0 (
          nx8553), .A1 (RST), .A2 (nx7865), .B0 (nx3789), .B1 (nx3869)) ;
    oai32 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix433 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .A0 (
          nx8553), .A1 (RST), .A2 (nx7865), .B0 (nx3793), .B1 (nx3869)) ;
    oai32 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix443 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .A0 (
          nx8555), .A1 (RST), .A2 (nx7865), .B0 (nx3797), .B1 (nx3869)) ;
    oai32 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix453 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .A0 (
          nx8555), .A1 (RST), .A2 (nx7867), .B0 (nx3801), .B1 (nx3869)) ;
    oai32 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix463 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .A0 (
          nx8555), .A1 (RST), .A2 (nx7867), .B0 (nx3805), .B1 (nx3871)) ;
    oai32 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix473 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .A0 (
          nx8555), .A1 (RST), .A2 (nx7867), .B0 (nx3809), .B1 (nx3871)) ;
    oai32 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix483 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .A0 (
          nx3851), .A1 (RST), .A2 (nx7867), .B0 (nx3813), .B1 (nx3871)) ;
    oai32 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix493 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .A0 (
          nx3873), .A1 (RST), .A2 (nx7867), .B0 (nx3817), .B1 (nx3871)) ;
    inv01 ix3872 (.Y (nx3873), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_10)) ;
    oai32 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix503 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .A0 (
          nx3875), .A1 (RST), .A2 (nx7867), .B0 (nx3821), .B1 (nx3871)) ;
    inv01 ix3874 (.Y (nx3875), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_11)) ;
    oai32 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix513 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .A0 (
          nx3877), .A1 (RST), .A2 (nx7867), .B0 (nx3825), .B1 (nx3871)) ;
    inv01 ix3876 (.Y (nx3877), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_12)) ;
    oai32 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix523 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .A0 (
          nx3879), .A1 (RST), .A2 (nx7869), .B0 (nx3829), .B1 (nx3871)) ;
    inv01 ix3878 (.Y (nx3879), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_13)) ;
    oai32 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix533 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .A0 (
          nx3881), .A1 (RST), .A2 (nx7869), .B0 (nx3833), .B1 (nx3883)) ;
    inv01 ix3880 (.Y (nx3881), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_14)) ;
    inv01 ix3882 (.Y (nx3883), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566)) ;
    oai32 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix543 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .A0 (
          nx3885), .A1 (RST), .A2 (nx7869), .B0 (nx3837), .B1 (nx3883)) ;
    inv01 ix3884 (.Y (nx3885), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_15)) ;
    oai32 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix553 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .A0 (
          nx3887), .A1 (RST), .A2 (nx7869), .B0 (nx3841), .B1 (nx3883)) ;
    inv01 ix3886 (.Y (nx3887), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_16)) ;
    nand02_2x CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix633 (.Y (
              nx3869), .A0 (nx7357), .A1 (nx7869)) ;
    nand02_2x CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix635 (.Y (
              nx3871), .A0 (nx7357), .A1 (nx7869)) ;
    oai32 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix393 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .A0 (
          nx3889), .A1 (RST), .A2 (nx7871), .B0 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx384), .B1 (nx3891)) ;
    inv01 ix3888 (.Y (nx3889), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_0)) ;
    oai32 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix403 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .A0 (
          nx3893), .A1 (RST), .A2 (nx7871), .B0 (nx3709), .B1 (nx3891)) ;
    inv01 ix3892 (.Y (nx3893), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_1)) ;
    oai32 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix413 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .A0 (
          nx3895), .A1 (RST), .A2 (nx7871), .B0 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx387), .B1 (nx3891)) ;
    inv01 ix3894 (.Y (nx3895), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_2)) ;
    oai32 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix423 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .A0 (
          nx3897), .A1 (RST), .A2 (nx7871), .B0 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx399), .B1 (nx3891)) ;
    inv01 ix3896 (.Y (nx3897), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_3)) ;
    oai32 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix433 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .A0 (
          nx3899), .A1 (RST), .A2 (nx7871), .B0 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx409), .B1 (nx3891)) ;
    inv01 ix3898 (.Y (nx3899), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_4)) ;
    oai32 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix443 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .A0 (
          nx3901), .A1 (RST), .A2 (nx7871), .B0 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx419), .B1 (nx3891)) ;
    inv01 ix3900 (.Y (nx3901), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_5)) ;
    oai32 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix453 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .A0 (
          nx3903), .A1 (RST), .A2 (nx7871), .B0 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx429), .B1 (nx3891)) ;
    inv01 ix3902 (.Y (nx3903), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_6)) ;
    oai32 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix463 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .A0 (
          nx3905), .A1 (RST), .A2 (nx7873), .B0 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx439), .B1 (nx3907)) ;
    inv01 ix3904 (.Y (nx3905), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_7)) ;
    oai32 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix473 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .A0 (
          nx3909), .A1 (RST), .A2 (nx7873), .B0 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx449), .B1 (nx3907)) ;
    inv01 ix3908 (.Y (nx3909), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_8)) ;
    oai32 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix483 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .A0 (
          nx3911), .A1 (RST), .A2 (nx7873), .B0 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx469), .B1 (nx3907)) ;
    inv01 ix3910 (.Y (nx3911), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_9)) ;
    oai32 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix493 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .A0 (
          nx3913), .A1 (RST), .A2 (nx7873), .B0 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx477), .B1 (nx3907)) ;
    inv01 ix3912 (.Y (nx3913), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_10)) ;
    oai32 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix503 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .A0 (
          nx3915), .A1 (RST), .A2 (nx7873), .B0 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx485), .B1 (nx3907)) ;
    inv01 ix3914 (.Y (nx3915), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_11)) ;
    oai32 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix513 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .A0 (
          nx3917), .A1 (RST), .A2 (nx7873), .B0 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx493), .B1 (nx3907)) ;
    inv01 ix3916 (.Y (nx3917), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_12)) ;
    oai32 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix523 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .A0 (
          nx3919), .A1 (RST), .A2 (nx7873), .B0 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx501), .B1 (nx3907)) ;
    inv01 ix3918 (.Y (nx3919), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_13)) ;
    oai32 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix533 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .A0 (
          nx3921), .A1 (RST), .A2 (nx7875), .B0 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx509), .B1 (nx3923)) ;
    inv01 ix3920 (.Y (nx3921), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_14)) ;
    inv01 ix3922 (.Y (nx3923), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566)) ;
    oai32 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix543 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .A0 (
          nx3925), .A1 (RST), .A2 (nx7875), .B0 (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_nx517), .B1 (nx3923)) ;
    inv01 ix3924 (.Y (nx3925), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_15)) ;
    oai32 CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix553 (.Y (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .A0 (
          nx3927), .A1 (RST), .A2 (nx7875), .B0 (nx3725), .B1 (nx3923)) ;
    inv01 ix3926 (.Y (nx3927), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_16)) ;
    nand02_2x CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix633 (.Y (
              nx3891), .A0 (nx7359), .A1 (nx7875)) ;
    nand02_2x CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix635 (.Y (
              nx3907), .A0 (nx7359), .A1 (nx7875)) ;
    mux21 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix404 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx403), .A0 (nx3929), .A1 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_2), .S0 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx395)) ;
    inv01 ix3928 (.Y (nx3929), .A (CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx391)) ;
    mux21 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix414 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx413), .A0 (nx3931), .A1 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_3), .S0 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx405)) ;
    inv01 ix3930 (.Y (nx3931), .A (CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx403)) ;
    mux21 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix424 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx423), .A0 (nx3933), .A1 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_4), .S0 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx415)) ;
    inv01 ix3932 (.Y (nx3933), .A (CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx413)) ;
    mux21 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix434 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx433), .A0 (nx3935), .A1 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_5), .S0 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx425)) ;
    inv01 ix3934 (.Y (nx3935), .A (CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx423)) ;
    mux21 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix444 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx443), .A0 (nx3937), .A1 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_6), .S0 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx435)) ;
    inv01 ix3936 (.Y (nx3937), .A (CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx433)) ;
    mux21 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix454 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx453), .A0 (nx3939), .A1 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_7), .S0 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx445)) ;
    inv01 ix3938 (.Y (nx3939), .A (CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx443)) ;
    mux21 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix462 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx461), .A0 (nx3941), .A1 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_8), .S0 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx455)) ;
    inv01 ix3940 (.Y (nx3941), .A (CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx453)) ;
    mux21 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix468 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx467), .A0 (nx3943), .A1 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_9), .S0 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx463)) ;
    inv01 ix3942 (.Y (nx3943), .A (CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx461)) ;
    mux21 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix476 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx475), .A0 (nx3945), .A1 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_10), .S0 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx471)) ;
    inv01 ix3944 (.Y (nx3945), .A (CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx467)) ;
    mux21 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix484 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx483), .A0 (nx3947), .A1 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_11), .S0 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx479)) ;
    inv01 ix3946 (.Y (nx3947), .A (CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx475)) ;
    mux21 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix492 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx491), .A0 (nx3949), .A1 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_12), .S0 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx487)) ;
    inv01 ix3948 (.Y (nx3949), .A (CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx483)) ;
    mux21 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix500 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx499), .A0 (nx3951), .A1 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_13), .S0 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx495)) ;
    inv01 ix3950 (.Y (nx3951), .A (CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx491)) ;
    mux21 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix508 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx507), .A0 (nx3953), .A1 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_14), .S0 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx503)) ;
    inv01 ix3952 (.Y (nx3953), .A (CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx499)) ;
    mux21 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix516 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx515), .A0 (nx3955), .A1 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_15), .S0 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx511)) ;
    inv01 ix3954 (.Y (nx3955), .A (CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx507)) ;
    mux21 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix161 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_1), .A0 (nx3957), .A1 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx379), .S0 (nx7879)) ;
    inv01 ix3956 (.Y (nx3957), .A (CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_1)) ;
    mux21 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix181 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_2), .A0 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx387), .A1 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx389), .S0 (nx7879)) ;
    mux21 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix201 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_3), .A0 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx399), .A1 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx401), .S0 (nx7879)) ;
    mux21 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix221 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_4), .A0 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx409), .A1 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx411), .S0 (nx7879)) ;
    mux21 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix241 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_5), .A0 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx419), .A1 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx421), .S0 (nx7879)) ;
    mux21 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix261 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_6), .A0 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx429), .A1 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx431), .S0 (nx7879)) ;
    mux21 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix281 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_7), .A0 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx439), .A1 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx441), .S0 (nx7879)) ;
    mux21 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix301 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_8), .A0 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx449), .A1 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx451), .S0 (nx7881)) ;
    mux21 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix321 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_9), .A0 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx469), .A1 (nx3959), .S0 (nx7881)) ;
    inv01 ix3958 (.Y (nx3959), .A (CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx316)) ;
    mux21 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix341 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_10), .A0 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx477), .A1 (nx3961), .S0 (nx7881)) ;
    inv01 ix3960 (.Y (nx3961), .A (CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx336)) ;
    mux21 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix361 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_11), .A0 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx485), .A1 (nx3963), .S0 (nx7881)) ;
    inv01 ix3962 (.Y (nx3963), .A (CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx356)) ;
    mux21 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix381 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_12), .A0 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx493), .A1 (nx3965), .S0 (nx7881)) ;
    inv01 ix3964 (.Y (nx3965), .A (CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx376)) ;
    mux21 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix401 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_13), .A0 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx501), .A1 (nx3967), .S0 (nx7881)) ;
    inv01 ix3966 (.Y (nx3967), .A (CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx396)) ;
    mux21 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix421 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_14), .A0 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx509), .A1 (nx3969), .S0 (nx7881)) ;
    inv01 ix3968 (.Y (nx3969), .A (CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx416)) ;
    mux21 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix441 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_15), .A0 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx517), .A1 (nx3971), .S0 (nx7883)) ;
    inv01 ix3970 (.Y (nx3971), .A (CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx436)) ;
    mux21 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_ix461 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_16), .A0 (nx3973), 
          .A1 (nx3975), .S0 (nx7883)) ;
    inv01 ix3972 (.Y (nx3973), .A (CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothP_16)
          ) ;
    inv01 ix3974 (.Y (nx3975), .A (CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx456)) ;
    nor02_2x CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix81 (.Y (
             CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx80), .A0 (Instr), .A1 (
             nx7309)) ;
    nor02_2x CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix319 (.Y (
             CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642), .A0 (
             CALCULATOR_Start_dup_1209), .A1 (
             CALCULATOR_CalculatingBooth_dup_1181)) ;
    nor02_2x CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix85 (.Y (
             CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_0), .A0 (
             nx7893), .A1 (nx3977)) ;
    inv01 ix3976 (.Y (nx3977), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_1)) ;
    mux21 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix125 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_1), .A0 (
          nx3979), .A1 (nx3981), .S0 (nx7893)) ;
    inv01 ix3978 (.Y (nx3979), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_2)) ;
    inv01 ix3980 (.Y (nx3981), .A (CacheWindow_2__3__0)) ;
    mux21 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix133 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_2), .A0 (
          nx3983), .A1 (nx3985), .S0 (nx7893)) ;
    inv01 ix3982 (.Y (nx3983), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_3)) ;
    inv01 ix3984 (.Y (nx3985), .A (CacheWindow_2__3__1)) ;
    mux21 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix141 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_3), .A0 (
          nx3987), .A1 (nx3989), .S0 (nx7893)) ;
    inv01 ix3986 (.Y (nx3987), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_4)) ;
    inv01 ix3988 (.Y (nx3989), .A (CacheWindow_2__3__2)) ;
    mux21 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix149 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_4), .A0 (
          nx3991), .A1 (nx3993), .S0 (nx7893)) ;
    inv01 ix3990 (.Y (nx3991), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_5)) ;
    inv01 ix3992 (.Y (nx3993), .A (CacheWindow_2__3__3)) ;
    mux21 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix157 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_5), .A0 (
          nx3995), .A1 (nx3997), .S0 (nx7893)) ;
    inv01 ix3994 (.Y (nx3995), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_6)) ;
    inv01 ix3996 (.Y (nx3997), .A (CacheWindow_2__3__4)) ;
    mux21 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix165 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_6), .A0 (
          nx3999), .A1 (nx4001), .S0 (nx7893)) ;
    inv01 ix3998 (.Y (nx3999), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_7)) ;
    inv01 ix4000 (.Y (nx4001), .A (CacheWindow_2__3__5)) ;
    mux21 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix173 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_7), .A0 (
          nx4003), .A1 (nx4005), .S0 (nx7895)) ;
    inv01 ix4002 (.Y (nx4003), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_8)) ;
    inv01 ix4004 (.Y (nx4005), .A (CacheWindow_2__3__6)) ;
    mux21 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix181 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_8), .A0 (
          nx4007), .A1 (nx4009), .S0 (nx7895)) ;
    inv01 ix4006 (.Y (nx4007), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_9)) ;
    inv01 ix4008 (.Y (nx4009), .A (CacheWindow_2__3__7)) ;
    nor02_2x CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix89 (.Y (
             CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_9), .A0 (
             nx7895), .A1 (nx4011)) ;
    inv01 ix4010 (.Y (nx4011), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_10)) ;
    nor02_2x CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix93 (.Y (
             CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_10), .A0 (
             nx7895), .A1 (nx4013)) ;
    inv01 ix4012 (.Y (nx4013), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_11)) ;
    nor02_2x CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix97 (.Y (
             CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_11), .A0 (
             nx7895), .A1 (nx4015)) ;
    inv01 ix4014 (.Y (nx4015), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_12)) ;
    nor02_2x CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix101 (.Y (
             CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_12), .A0 (
             nx7895), .A1 (nx4017)) ;
    inv01 ix4016 (.Y (nx4017), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_13)) ;
    nor02_2x CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix105 (.Y (
             CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_13), .A0 (
             nx7895), .A1 (nx4019)) ;
    inv01 ix4018 (.Y (nx4019), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_14)) ;
    nor02_2x CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix109 (.Y (
             CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_14), .A0 (
             nx7897), .A1 (nx4021)) ;
    inv01 ix4020 (.Y (nx4021), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_15)) ;
    nor02_2x CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix113 (.Y (
             CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_15), .A0 (
             nx7897), .A1 (nx4023)) ;
    inv01 ix4022 (.Y (nx4023), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_16)) ;
    nor02_2x CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix117 (.Y (
             CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_16), .A0 (
             nx7897), .A1 (nx4023)) ;
    mux21 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix189 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothOperand_0), .A0 (nx4025), .A1 (
          nx4027), .S0 (nx7885)) ;
    inv01 ix4024 (.Y (nx4025), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_0)) ;
    inv01 ix4026 (.Y (nx4027), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_0)) ;
    mux21 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix197 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothOperand_1), .A0 (nx4029), .A1 (
          nx4031), .S0 (nx7885)) ;
    inv01 ix4028 (.Y (nx4029), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_1)) ;
    inv01 ix4030 (.Y (nx4031), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_1)) ;
    mux21 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix205 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothOperand_2), .A0 (nx4033), .A1 (
          nx4035), .S0 (nx7885)) ;
    inv01 ix4032 (.Y (nx4033), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_2)) ;
    inv01 ix4034 (.Y (nx4035), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_2)) ;
    mux21 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix213 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothOperand_3), .A0 (nx4037), .A1 (
          nx4039), .S0 (nx7885)) ;
    inv01 ix4036 (.Y (nx4037), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_3)) ;
    inv01 ix4038 (.Y (nx4039), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_3)) ;
    mux21 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix221 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothOperand_4), .A0 (nx4041), .A1 (
          nx4043), .S0 (nx7885)) ;
    inv01 ix4040 (.Y (nx4041), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_4)) ;
    inv01 ix4042 (.Y (nx4043), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_4)) ;
    mux21 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix229 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothOperand_5), .A0 (nx4045), .A1 (
          nx4047), .S0 (nx7887)) ;
    inv01 ix4044 (.Y (nx4045), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_5)) ;
    inv01 ix4046 (.Y (nx4047), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_5)) ;
    mux21 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix237 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothOperand_6), .A0 (nx4049), .A1 (
          nx4051), .S0 (nx7887)) ;
    inv01 ix4048 (.Y (nx4049), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_6)) ;
    inv01 ix4050 (.Y (nx4051), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_6)) ;
    mux21 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix245 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothOperand_7), .A0 (nx4053), .A1 (
          nx4055), .S0 (nx7887)) ;
    inv01 ix4052 (.Y (nx4053), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_7)) ;
    inv01 ix4054 (.Y (nx4055), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_7)) ;
    mux21 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix253 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothOperand_8), .A0 (nx4057), .A1 (
          nx4059), .S0 (nx7887)) ;
    inv01 ix4056 (.Y (nx4057), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_8)) ;
    inv01 ix4058 (.Y (nx4059), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_8)) ;
    mux21 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix261 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothOperand_9), .A0 (nx4061), .A1 (
          nx4063), .S0 (nx7887)) ;
    inv01 ix4060 (.Y (nx4061), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_9)) ;
    inv01 ix4062 (.Y (nx4063), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_9)) ;
    mux21 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix269 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothOperand_10), .A0 (nx4065), .A1 (
          nx4067), .S0 (nx7887)) ;
    inv01 ix4064 (.Y (nx4065), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_10)) ;
    inv01 ix4066 (.Y (nx4067), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_10)) ;
    mux21 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix277 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothOperand_11), .A0 (nx4069), .A1 (
          nx4071), .S0 (nx7887)) ;
    inv01 ix4068 (.Y (nx4069), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_11)) ;
    inv01 ix4070 (.Y (nx4071), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_11)) ;
    mux21 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix285 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothOperand_12), .A0 (nx4073), .A1 (
          nx4075), .S0 (nx7889)) ;
    inv01 ix4072 (.Y (nx4073), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_12)) ;
    inv01 ix4074 (.Y (nx4075), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_12)) ;
    mux21 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix293 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothOperand_13), .A0 (nx4077), .A1 (
          nx4079), .S0 (nx7889)) ;
    inv01 ix4076 (.Y (nx4077), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_13)) ;
    inv01 ix4078 (.Y (nx4079), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_13)) ;
    mux21 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix301 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothOperand_14), .A0 (nx4081), .A1 (
          nx4083), .S0 (nx7889)) ;
    inv01 ix4080 (.Y (nx4081), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_14)) ;
    inv01 ix4082 (.Y (nx4083), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_14)) ;
    mux21 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix309 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothOperand_15), .A0 (nx4085), .A1 (
          nx4087), .S0 (nx7889)) ;
    inv01 ix4084 (.Y (nx4085), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_15)) ;
    inv01 ix4086 (.Y (nx4087), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_15)) ;
    mux21 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix317 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BoothOperand_16), .A0 (nx4089), .A1 (
          nx4091), .S0 (nx7889)) ;
    inv01 ix4088 (.Y (nx4089), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_16)) ;
    inv01 ix4090 (.Y (nx4091), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_16)) ;
    xnor2 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix321 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_AddPToBoothOperand), .A0 (nx7889), .A1 (
          nx3957)) ;
    oai32 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix393 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .A0 (
          nx8557), .A1 (RST), .A2 (nx7899), .B0 (nx4027), .B1 (nx4095)) ;
    oai32 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix403 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .A0 (
          nx8557), .A1 (RST), .A2 (nx7899), .B0 (nx4031), .B1 (nx4095)) ;
    oai32 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix413 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .A0 (
          nx8557), .A1 (RST), .A2 (nx7899), .B0 (nx4035), .B1 (nx4095)) ;
    oai32 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix423 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .A0 (
          nx8557), .A1 (RST), .A2 (nx7899), .B0 (nx4039), .B1 (nx4095)) ;
    oai32 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix433 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .A0 (
          nx8557), .A1 (RST), .A2 (nx7899), .B0 (nx4043), .B1 (nx4095)) ;
    oai32 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix443 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .A0 (
          nx8557), .A1 (RST), .A2 (nx7899), .B0 (nx4047), .B1 (nx4095)) ;
    oai32 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix453 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .A0 (
          nx8557), .A1 (RST), .A2 (nx7901), .B0 (nx4051), .B1 (nx4095)) ;
    oai32 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix463 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .A0 (
          nx8559), .A1 (RST), .A2 (nx7901), .B0 (nx4055), .B1 (nx4097)) ;
    oai32 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix473 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .A0 (
          nx8559), .A1 (RST), .A2 (nx7901), .B0 (nx4059), .B1 (nx4097)) ;
    oai32 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix483 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .A0 (
          nx4099), .A1 (RST), .A2 (nx7901), .B0 (nx4063), .B1 (nx4097)) ;
    inv01 ix4098 (.Y (nx4099), .A (CacheFilter_2__3__0)) ;
    oai32 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix493 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .A0 (
          nx4101), .A1 (RST), .A2 (nx7901), .B0 (nx4067), .B1 (nx4097)) ;
    inv01 ix4100 (.Y (nx4101), .A (CacheFilter_2__3__1)) ;
    oai32 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix503 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .A0 (
          nx4103), .A1 (RST), .A2 (nx7901), .B0 (nx4071), .B1 (nx4097)) ;
    inv01 ix4102 (.Y (nx4103), .A (CacheFilter_2__3__2)) ;
    oai32 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix513 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .A0 (
          nx4105), .A1 (RST), .A2 (nx7901), .B0 (nx4075), .B1 (nx4097)) ;
    inv01 ix4104 (.Y (nx4105), .A (CacheFilter_2__3__3)) ;
    oai32 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix523 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .A0 (
          nx4107), .A1 (RST), .A2 (nx7903), .B0 (nx4079), .B1 (nx4097)) ;
    inv01 ix4106 (.Y (nx4107), .A (CacheFilter_2__3__4)) ;
    oai32 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix533 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .A0 (
          nx4109), .A1 (RST), .A2 (nx7903), .B0 (nx4083), .B1 (nx4111)) ;
    inv01 ix4108 (.Y (nx4109), .A (CacheFilter_2__3__5)) ;
    inv01 ix4110 (.Y (nx4111), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566)) ;
    oai32 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix543 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .A0 (
          nx4113), .A1 (RST), .A2 (nx7903), .B0 (nx4087), .B1 (nx4111)) ;
    inv01 ix4112 (.Y (nx4113), .A (CacheFilter_2__3__6)) ;
    oai32 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix553 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .A0 (
          nx4115), .A1 (RST), .A2 (nx7903), .B0 (nx4091), .B1 (nx4111)) ;
    inv01 ix4114 (.Y (nx4115), .A (CacheFilter_2__3__7)) ;
    nand02_2x CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix633 (.Y (
              nx4095), .A0 (nx7359), .A1 (nx7903)) ;
    nand02_2x CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix635 (.Y (
              nx4097), .A0 (nx7359), .A1 (nx7903)) ;
    oai32 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix393 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .A0 (
          nx8559), .A1 (RST), .A2 (nx7905), .B0 (nx4025), .B1 (nx4117)) ;
    oai32 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix403 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .A0 (
          nx8559), .A1 (RST), .A2 (nx7905), .B0 (nx4029), .B1 (nx4117)) ;
    oai32 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix413 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .A0 (
          nx8559), .A1 (RST), .A2 (nx7905), .B0 (nx4033), .B1 (nx4117)) ;
    oai32 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix423 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .A0 (
          nx8559), .A1 (RST), .A2 (nx7905), .B0 (nx4037), .B1 (nx4117)) ;
    oai32 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix433 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .A0 (
          nx8559), .A1 (RST), .A2 (nx7905), .B0 (nx4041), .B1 (nx4117)) ;
    oai32 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix443 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .A0 (
          nx8561), .A1 (RST), .A2 (nx7905), .B0 (nx4045), .B1 (nx4117)) ;
    oai32 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix453 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .A0 (
          nx8561), .A1 (RST), .A2 (nx7907), .B0 (nx4049), .B1 (nx4117)) ;
    oai32 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix463 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .A0 (
          nx8561), .A1 (RST), .A2 (nx7907), .B0 (nx4053), .B1 (nx4119)) ;
    oai32 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix473 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .A0 (
          nx8561), .A1 (RST), .A2 (nx7907), .B0 (nx4057), .B1 (nx4119)) ;
    oai32 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix483 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .A0 (
          nx4099), .A1 (RST), .A2 (nx7907), .B0 (nx4061), .B1 (nx4119)) ;
    oai32 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix493 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .A0 (
          nx4121), .A1 (RST), .A2 (nx7907), .B0 (nx4065), .B1 (nx4119)) ;
    inv01 ix4120 (.Y (nx4121), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_10)) ;
    oai32 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix503 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .A0 (
          nx4123), .A1 (RST), .A2 (nx7907), .B0 (nx4069), .B1 (nx4119)) ;
    inv01 ix4122 (.Y (nx4123), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_11)) ;
    oai32 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix513 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .A0 (
          nx4125), .A1 (RST), .A2 (nx7907), .B0 (nx4073), .B1 (nx4119)) ;
    inv01 ix4124 (.Y (nx4125), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_12)) ;
    oai32 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix523 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .A0 (
          nx4127), .A1 (RST), .A2 (nx7909), .B0 (nx4077), .B1 (nx4119)) ;
    inv01 ix4126 (.Y (nx4127), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_13)) ;
    oai32 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix533 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .A0 (
          nx4129), .A1 (RST), .A2 (nx7909), .B0 (nx4081), .B1 (nx4131)) ;
    inv01 ix4128 (.Y (nx4129), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_14)) ;
    inv01 ix4130 (.Y (nx4131), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566)) ;
    oai32 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix543 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .A0 (
          nx4133), .A1 (RST), .A2 (nx7909), .B0 (nx4085), .B1 (nx4131)) ;
    inv01 ix4132 (.Y (nx4133), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_15)) ;
    oai32 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix553 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .A0 (
          nx4135), .A1 (RST), .A2 (nx7909), .B0 (nx4089), .B1 (nx4131)) ;
    inv01 ix4134 (.Y (nx4135), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_16)) ;
    nand02_2x CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix633 (.Y (
              nx4117), .A0 (nx7359), .A1 (nx7909)) ;
    nand02_2x CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix635 (.Y (
              nx4119), .A0 (nx7359), .A1 (nx7909)) ;
    oai32 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix393 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .A0 (
          nx4137), .A1 (RST), .A2 (nx7911), .B0 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx384), .B1 (nx4139)) ;
    inv01 ix4136 (.Y (nx4137), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_0)) ;
    oai32 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix403 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .A0 (
          nx4141), .A1 (RST), .A2 (nx7911), .B0 (nx3957), .B1 (nx4139)) ;
    inv01 ix4140 (.Y (nx4141), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_1)) ;
    oai32 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix413 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .A0 (
          nx4143), .A1 (RST), .A2 (nx7911), .B0 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx387), .B1 (nx4139)) ;
    inv01 ix4142 (.Y (nx4143), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_2)) ;
    oai32 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix423 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .A0 (
          nx4145), .A1 (RST), .A2 (nx7911), .B0 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx399), .B1 (nx4139)) ;
    inv01 ix4144 (.Y (nx4145), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_3)) ;
    oai32 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix433 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .A0 (
          nx4147), .A1 (RST), .A2 (nx7911), .B0 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx409), .B1 (nx4139)) ;
    inv01 ix4146 (.Y (nx4147), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_4)) ;
    oai32 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix443 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .A0 (
          nx4149), .A1 (RST), .A2 (nx7911), .B0 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx419), .B1 (nx4139)) ;
    inv01 ix4148 (.Y (nx4149), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_5)) ;
    oai32 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix453 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .A0 (
          nx4151), .A1 (RST), .A2 (nx7911), .B0 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx429), .B1 (nx4139)) ;
    inv01 ix4150 (.Y (nx4151), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_6)) ;
    oai32 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix463 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .A0 (
          nx4153), .A1 (RST), .A2 (nx7913), .B0 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx439), .B1 (nx4155)) ;
    inv01 ix4152 (.Y (nx4153), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_7)) ;
    oai32 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix473 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .A0 (
          nx4157), .A1 (RST), .A2 (nx7913), .B0 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx449), .B1 (nx4155)) ;
    inv01 ix4156 (.Y (nx4157), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_8)) ;
    oai32 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix483 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .A0 (
          nx4159), .A1 (RST), .A2 (nx7913), .B0 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx469), .B1 (nx4155)) ;
    inv01 ix4158 (.Y (nx4159), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_9)) ;
    oai32 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix493 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .A0 (
          nx4161), .A1 (RST), .A2 (nx7913), .B0 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx477), .B1 (nx4155)) ;
    inv01 ix4160 (.Y (nx4161), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_10)) ;
    oai32 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix503 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .A0 (
          nx4163), .A1 (RST), .A2 (nx7913), .B0 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx485), .B1 (nx4155)) ;
    inv01 ix4162 (.Y (nx4163), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_11)) ;
    oai32 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix513 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .A0 (
          nx4165), .A1 (RST), .A2 (nx7913), .B0 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx493), .B1 (nx4155)) ;
    inv01 ix4164 (.Y (nx4165), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_12)) ;
    oai32 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix523 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .A0 (
          nx4167), .A1 (RST), .A2 (nx7913), .B0 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx501), .B1 (nx4155)) ;
    inv01 ix4166 (.Y (nx4167), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_13)) ;
    oai32 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix533 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .A0 (
          nx4169), .A1 (RST), .A2 (nx7915), .B0 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx509), .B1 (nx4171)) ;
    inv01 ix4168 (.Y (nx4169), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_14)) ;
    inv01 ix4170 (.Y (nx4171), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566)) ;
    oai32 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix543 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .A0 (
          nx4173), .A1 (RST), .A2 (nx7915), .B0 (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_nx517), .B1 (nx4171)) ;
    inv01 ix4172 (.Y (nx4173), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_15)) ;
    oai32 CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix553 (.Y (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .A0 (
          nx4175), .A1 (RST), .A2 (nx7915), .B0 (nx3973), .B1 (nx4171)) ;
    inv01 ix4174 (.Y (nx4175), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_16)) ;
    nand02_2x CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix633 (.Y (
              nx4139), .A0 (nx7359), .A1 (nx7915)) ;
    nand02_2x CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix635 (.Y (
              nx4155), .A0 (nx7361), .A1 (nx7915)) ;
    mux21 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix404 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx403), .A0 (nx4177), .A1 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_2), .S0 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx395)) ;
    inv01 ix4176 (.Y (nx4177), .A (CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx391)) ;
    mux21 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix414 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx413), .A0 (nx4179), .A1 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_3), .S0 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx405)) ;
    inv01 ix4178 (.Y (nx4179), .A (CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx403)) ;
    mux21 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix424 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx423), .A0 (nx4181), .A1 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_4), .S0 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx415)) ;
    inv01 ix4180 (.Y (nx4181), .A (CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx413)) ;
    mux21 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix434 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx433), .A0 (nx4183), .A1 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_5), .S0 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx425)) ;
    inv01 ix4182 (.Y (nx4183), .A (CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx423)) ;
    mux21 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix444 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx443), .A0 (nx4185), .A1 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_6), .S0 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx435)) ;
    inv01 ix4184 (.Y (nx4185), .A (CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx433)) ;
    mux21 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix454 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx453), .A0 (nx4187), .A1 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_7), .S0 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx445)) ;
    inv01 ix4186 (.Y (nx4187), .A (CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx443)) ;
    mux21 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix462 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx461), .A0 (nx4189), .A1 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_8), .S0 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx455)) ;
    inv01 ix4188 (.Y (nx4189), .A (CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx453)) ;
    mux21 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix468 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx467), .A0 (nx4191), .A1 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_9), .S0 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx463)) ;
    inv01 ix4190 (.Y (nx4191), .A (CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx461)) ;
    mux21 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix476 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx475), .A0 (nx4193), .A1 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_10), .S0 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx471)) ;
    inv01 ix4192 (.Y (nx4193), .A (CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx467)) ;
    mux21 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix484 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx483), .A0 (nx4195), .A1 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_11), .S0 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx479)) ;
    inv01 ix4194 (.Y (nx4195), .A (CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx475)) ;
    mux21 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix492 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx491), .A0 (nx4197), .A1 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_12), .S0 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx487)) ;
    inv01 ix4196 (.Y (nx4197), .A (CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx483)) ;
    mux21 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix500 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx499), .A0 (nx4199), .A1 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_13), .S0 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx495)) ;
    inv01 ix4198 (.Y (nx4199), .A (CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx491)) ;
    mux21 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix508 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx507), .A0 (nx4201), .A1 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_14), .S0 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx503)) ;
    inv01 ix4200 (.Y (nx4201), .A (CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx499)) ;
    mux21 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix516 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx515), .A0 (nx4203), .A1 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_15), .S0 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx511)) ;
    inv01 ix4202 (.Y (nx4203), .A (CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx507)) ;
    mux21 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix161 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_1), .A0 (nx4205), .A1 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx379), .S0 (nx7919)) ;
    inv01 ix4204 (.Y (nx4205), .A (CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_1)) ;
    mux21 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix181 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_2), .A0 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx387), .A1 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx389), .S0 (nx7919)) ;
    mux21 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix201 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_3), .A0 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx399), .A1 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx401), .S0 (nx7919)) ;
    mux21 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix221 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_4), .A0 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx409), .A1 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx411), .S0 (nx7919)) ;
    mux21 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix241 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_5), .A0 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx419), .A1 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx421), .S0 (nx7919)) ;
    mux21 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix261 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_6), .A0 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx429), .A1 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx431), .S0 (nx7919)) ;
    mux21 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix281 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_7), .A0 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx439), .A1 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx441), .S0 (nx7919)) ;
    mux21 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix301 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_8), .A0 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx449), .A1 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx451), .S0 (nx7921)) ;
    mux21 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix321 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_9), .A0 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx469), .A1 (nx4207), .S0 (nx7921)) ;
    inv01 ix4206 (.Y (nx4207), .A (CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx316)) ;
    mux21 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix341 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_10), .A0 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx477), .A1 (nx4209), .S0 (nx7921)) ;
    inv01 ix4208 (.Y (nx4209), .A (CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx336)) ;
    mux21 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix361 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_11), .A0 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx485), .A1 (nx4211), .S0 (nx7921)) ;
    inv01 ix4210 (.Y (nx4211), .A (CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx356)) ;
    mux21 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix381 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_12), .A0 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx493), .A1 (nx4213), .S0 (nx7921)) ;
    inv01 ix4212 (.Y (nx4213), .A (CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx376)) ;
    mux21 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix401 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_13), .A0 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx501), .A1 (nx4215), .S0 (nx7921)) ;
    inv01 ix4214 (.Y (nx4215), .A (CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx396)) ;
    mux21 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix421 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_14), .A0 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx509), .A1 (nx4217), .S0 (nx7921)) ;
    inv01 ix4216 (.Y (nx4217), .A (CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx416)) ;
    mux21 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix441 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_15), .A0 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx517), .A1 (nx4219), .S0 (nx7923)) ;
    inv01 ix4218 (.Y (nx4219), .A (CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx436)) ;
    mux21 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_ix461 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_16), .A0 (nx4221), 
          .A1 (nx4223), .S0 (nx7923)) ;
    inv01 ix4220 (.Y (nx4221), .A (CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothP_16)
          ) ;
    inv01 ix4222 (.Y (nx4223), .A (CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx456)) ;
    nor02_2x CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix81 (.Y (
             CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_nx80), .A0 (Instr), .A1 (
             nx7313)) ;
    nor02_2x CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix319 (.Y (
             CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642), .A0 (
             CALCULATOR_Start_dup_1222), .A1 (
             CALCULATOR_CalculatingBooth_dup_1224)) ;
    nor02_2x CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix85 (.Y (
             CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_0), .A0 (
             nx7933), .A1 (nx4225)) ;
    inv01 ix4224 (.Y (nx4225), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_1)) ;
    mux21 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix125 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_1), .A0 (
          nx4227), .A1 (nx4229), .S0 (nx7933)) ;
    inv01 ix4226 (.Y (nx4227), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_2)) ;
    inv01 ix4228 (.Y (nx4229), .A (CacheWindow_2__4__0)) ;
    mux21 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix133 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_2), .A0 (
          nx4231), .A1 (nx4233), .S0 (nx7933)) ;
    inv01 ix4230 (.Y (nx4231), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_3)) ;
    inv01 ix4232 (.Y (nx4233), .A (CacheWindow_2__4__1)) ;
    mux21 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix141 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_3), .A0 (
          nx4235), .A1 (nx4237), .S0 (nx7933)) ;
    inv01 ix4234 (.Y (nx4235), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_4)) ;
    inv01 ix4236 (.Y (nx4237), .A (CacheWindow_2__4__2)) ;
    mux21 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix149 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_4), .A0 (
          nx4239), .A1 (nx4241), .S0 (nx7933)) ;
    inv01 ix4238 (.Y (nx4239), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_5)) ;
    inv01 ix4240 (.Y (nx4241), .A (CacheWindow_2__4__3)) ;
    mux21 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix157 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_5), .A0 (
          nx4243), .A1 (nx4245), .S0 (nx7933)) ;
    inv01 ix4242 (.Y (nx4243), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_6)) ;
    inv01 ix4244 (.Y (nx4245), .A (CacheWindow_2__4__4)) ;
    mux21 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix165 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_6), .A0 (
          nx4247), .A1 (nx4249), .S0 (nx7933)) ;
    inv01 ix4246 (.Y (nx4247), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_7)) ;
    inv01 ix4248 (.Y (nx4249), .A (CacheWindow_2__4__5)) ;
    mux21 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix173 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_7), .A0 (
          nx4251), .A1 (nx4253), .S0 (nx7935)) ;
    inv01 ix4250 (.Y (nx4251), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_8)) ;
    inv01 ix4252 (.Y (nx4253), .A (CacheWindow_2__4__6)) ;
    mux21 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix181 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_8), .A0 (
          nx4255), .A1 (nx4257), .S0 (nx7935)) ;
    inv01 ix4254 (.Y (nx4255), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_9)) ;
    inv01 ix4256 (.Y (nx4257), .A (CacheWindow_2__4__7)) ;
    nor02_2x CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix89 (.Y (
             CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_9), .A0 (
             nx7935), .A1 (nx4259)) ;
    inv01 ix4258 (.Y (nx4259), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_10)) ;
    nor02_2x CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix93 (.Y (
             CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_10), .A0 (
             nx7935), .A1 (nx4261)) ;
    inv01 ix4260 (.Y (nx4261), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_11)) ;
    nor02_2x CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix97 (.Y (
             CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_11), .A0 (
             nx7935), .A1 (nx4263)) ;
    inv01 ix4262 (.Y (nx4263), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_12)) ;
    nor02_2x CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix101 (.Y (
             CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_12), .A0 (
             nx7935), .A1 (nx4265)) ;
    inv01 ix4264 (.Y (nx4265), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_13)) ;
    nor02_2x CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix105 (.Y (
             CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_13), .A0 (
             nx7935), .A1 (nx4267)) ;
    inv01 ix4266 (.Y (nx4267), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_14)) ;
    nor02_2x CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix109 (.Y (
             CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_14), .A0 (
             nx7937), .A1 (nx4269)) ;
    inv01 ix4268 (.Y (nx4269), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_15)) ;
    nor02_2x CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix113 (.Y (
             CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_15), .A0 (
             nx7937), .A1 (nx4271)) ;
    inv01 ix4270 (.Y (nx4271), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_16)) ;
    nor02_2x CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix117 (.Y (
             CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_16), .A0 (
             nx7937), .A1 (nx4271)) ;
    mux21 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix189 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothOperand_0), .A0 (nx4273), .A1 (
          nx4275), .S0 (nx7925)) ;
    inv01 ix4272 (.Y (nx4273), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_0)) ;
    inv01 ix4274 (.Y (nx4275), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_0)) ;
    mux21 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix197 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothOperand_1), .A0 (nx4277), .A1 (
          nx4279), .S0 (nx7925)) ;
    inv01 ix4276 (.Y (nx4277), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_1)) ;
    inv01 ix4278 (.Y (nx4279), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_1)) ;
    mux21 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix205 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothOperand_2), .A0 (nx4281), .A1 (
          nx4283), .S0 (nx7925)) ;
    inv01 ix4280 (.Y (nx4281), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_2)) ;
    inv01 ix4282 (.Y (nx4283), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_2)) ;
    mux21 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix213 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothOperand_3), .A0 (nx4285), .A1 (
          nx4287), .S0 (nx7925)) ;
    inv01 ix4284 (.Y (nx4285), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_3)) ;
    inv01 ix4286 (.Y (nx4287), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_3)) ;
    mux21 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix221 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothOperand_4), .A0 (nx4289), .A1 (
          nx4291), .S0 (nx7925)) ;
    inv01 ix4288 (.Y (nx4289), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_4)) ;
    inv01 ix4290 (.Y (nx4291), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_4)) ;
    mux21 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix229 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothOperand_5), .A0 (nx4293), .A1 (
          nx4295), .S0 (nx7927)) ;
    inv01 ix4292 (.Y (nx4293), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_5)) ;
    inv01 ix4294 (.Y (nx4295), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_5)) ;
    mux21 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix237 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothOperand_6), .A0 (nx4297), .A1 (
          nx4299), .S0 (nx7927)) ;
    inv01 ix4296 (.Y (nx4297), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_6)) ;
    inv01 ix4298 (.Y (nx4299), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_6)) ;
    mux21 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix245 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothOperand_7), .A0 (nx4301), .A1 (
          nx4303), .S0 (nx7927)) ;
    inv01 ix4300 (.Y (nx4301), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_7)) ;
    inv01 ix4302 (.Y (nx4303), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_7)) ;
    mux21 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix253 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothOperand_8), .A0 (nx4305), .A1 (
          nx4307), .S0 (nx7927)) ;
    inv01 ix4304 (.Y (nx4305), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_8)) ;
    inv01 ix4306 (.Y (nx4307), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_8)) ;
    mux21 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix261 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothOperand_9), .A0 (nx4309), .A1 (
          nx4311), .S0 (nx7927)) ;
    inv01 ix4308 (.Y (nx4309), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_9)) ;
    inv01 ix4310 (.Y (nx4311), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_9)) ;
    mux21 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix269 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothOperand_10), .A0 (nx4313), .A1 (
          nx4315), .S0 (nx7927)) ;
    inv01 ix4312 (.Y (nx4313), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_10)) ;
    inv01 ix4314 (.Y (nx4315), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_10)) ;
    mux21 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix277 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothOperand_11), .A0 (nx4317), .A1 (
          nx4319), .S0 (nx7927)) ;
    inv01 ix4316 (.Y (nx4317), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_11)) ;
    inv01 ix4318 (.Y (nx4319), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_11)) ;
    mux21 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix285 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothOperand_12), .A0 (nx4321), .A1 (
          nx4323), .S0 (nx7929)) ;
    inv01 ix4320 (.Y (nx4321), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_12)) ;
    inv01 ix4322 (.Y (nx4323), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_12)) ;
    mux21 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix293 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothOperand_13), .A0 (nx4325), .A1 (
          nx4327), .S0 (nx7929)) ;
    inv01 ix4324 (.Y (nx4325), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_13)) ;
    inv01 ix4326 (.Y (nx4327), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_13)) ;
    mux21 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix301 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothOperand_14), .A0 (nx4329), .A1 (
          nx4331), .S0 (nx7929)) ;
    inv01 ix4328 (.Y (nx4329), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_14)) ;
    inv01 ix4330 (.Y (nx4331), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_14)) ;
    mux21 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix309 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothOperand_15), .A0 (nx4333), .A1 (
          nx4335), .S0 (nx7929)) ;
    inv01 ix4332 (.Y (nx4333), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_15)) ;
    inv01 ix4334 (.Y (nx4335), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_15)) ;
    mux21 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix317 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BoothOperand_16), .A0 (nx4337), .A1 (
          nx4339), .S0 (nx7929)) ;
    inv01 ix4336 (.Y (nx4337), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_16)) ;
    inv01 ix4338 (.Y (nx4339), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_16)) ;
    xnor2 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix321 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_AddPToBoothOperand), .A0 (nx7929), .A1 (
          nx4205)) ;
    oai32 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix393 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .A0 (
          nx8563), .A1 (RST), .A2 (nx7939), .B0 (nx4275), .B1 (nx4343)) ;
    oai32 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix403 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .A0 (
          nx8563), .A1 (RST), .A2 (nx7939), .B0 (nx4279), .B1 (nx4343)) ;
    oai32 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix413 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .A0 (
          nx8563), .A1 (RST), .A2 (nx7939), .B0 (nx4283), .B1 (nx4343)) ;
    oai32 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix423 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .A0 (
          nx8563), .A1 (RST), .A2 (nx7939), .B0 (nx4287), .B1 (nx4343)) ;
    oai32 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix433 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .A0 (
          nx8563), .A1 (RST), .A2 (nx7939), .B0 (nx4291), .B1 (nx4343)) ;
    oai32 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix443 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .A0 (
          nx8563), .A1 (RST), .A2 (nx7939), .B0 (nx4295), .B1 (nx4343)) ;
    oai32 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix453 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .A0 (
          nx8563), .A1 (RST), .A2 (nx7941), .B0 (nx4299), .B1 (nx4343)) ;
    oai32 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix463 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .A0 (
          nx8565), .A1 (RST), .A2 (nx7941), .B0 (nx4303), .B1 (nx4345)) ;
    oai32 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix473 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .A0 (
          nx8565), .A1 (RST), .A2 (nx7941), .B0 (nx4307), .B1 (nx4345)) ;
    oai32 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix483 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .A0 (
          nx4347), .A1 (RST), .A2 (nx7941), .B0 (nx4311), .B1 (nx4345)) ;
    inv01 ix4346 (.Y (nx4347), .A (CacheFilter_2__4__0)) ;
    oai32 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix493 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .A0 (
          nx4349), .A1 (RST), .A2 (nx7941), .B0 (nx4315), .B1 (nx4345)) ;
    inv01 ix4348 (.Y (nx4349), .A (CacheFilter_2__4__1)) ;
    oai32 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix503 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .A0 (
          nx4351), .A1 (RST), .A2 (nx7941), .B0 (nx4319), .B1 (nx4345)) ;
    inv01 ix4350 (.Y (nx4351), .A (CacheFilter_2__4__2)) ;
    oai32 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix513 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .A0 (
          nx4353), .A1 (RST), .A2 (nx7941), .B0 (nx4323), .B1 (nx4345)) ;
    inv01 ix4352 (.Y (nx4353), .A (CacheFilter_2__4__3)) ;
    oai32 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix523 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .A0 (
          nx4355), .A1 (RST), .A2 (nx7943), .B0 (nx4327), .B1 (nx4345)) ;
    inv01 ix4354 (.Y (nx4355), .A (CacheFilter_2__4__4)) ;
    oai32 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix533 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .A0 (
          nx4357), .A1 (RST), .A2 (nx7943), .B0 (nx4331), .B1 (nx4359)) ;
    inv01 ix4356 (.Y (nx4357), .A (CacheFilter_2__4__5)) ;
    inv01 ix4358 (.Y (nx4359), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566)) ;
    oai32 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix543 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .A0 (
          nx4361), .A1 (RST), .A2 (nx7943), .B0 (nx4335), .B1 (nx4359)) ;
    inv01 ix4360 (.Y (nx4361), .A (CacheFilter_2__4__6)) ;
    oai32 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix553 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .A0 (
          nx4363), .A1 (RST), .A2 (nx7943), .B0 (nx4339), .B1 (nx4359)) ;
    inv01 ix4362 (.Y (nx4363), .A (CacheFilter_2__4__7)) ;
    nand02_2x CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix633 (.Y (
              nx4343), .A0 (nx7361), .A1 (nx7943)) ;
    nand02_2x CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix635 (.Y (
              nx4345), .A0 (nx7361), .A1 (nx7943)) ;
    oai32 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix393 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .A0 (
          nx8565), .A1 (RST), .A2 (nx7945), .B0 (nx4273), .B1 (nx4365)) ;
    oai32 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix403 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .A0 (
          nx8565), .A1 (RST), .A2 (nx7945), .B0 (nx4277), .B1 (nx4365)) ;
    oai32 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix413 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .A0 (
          nx8565), .A1 (RST), .A2 (nx7945), .B0 (nx4281), .B1 (nx4365)) ;
    oai32 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix423 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .A0 (
          nx8565), .A1 (RST), .A2 (nx7945), .B0 (nx4285), .B1 (nx4365)) ;
    oai32 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix433 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .A0 (
          nx8565), .A1 (RST), .A2 (nx7945), .B0 (nx4289), .B1 (nx4365)) ;
    oai32 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix443 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .A0 (
          nx8567), .A1 (RST), .A2 (nx7945), .B0 (nx4293), .B1 (nx4365)) ;
    oai32 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix453 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .A0 (
          nx8567), .A1 (RST), .A2 (nx7947), .B0 (nx4297), .B1 (nx4365)) ;
    oai32 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix463 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .A0 (
          nx8567), .A1 (RST), .A2 (nx7947), .B0 (nx4301), .B1 (nx4367)) ;
    oai32 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix473 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .A0 (
          nx8567), .A1 (RST), .A2 (nx7947), .B0 (nx4305), .B1 (nx4367)) ;
    oai32 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix483 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .A0 (
          nx4347), .A1 (RST), .A2 (nx7947), .B0 (nx4309), .B1 (nx4367)) ;
    oai32 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix493 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .A0 (
          nx4369), .A1 (RST), .A2 (nx7947), .B0 (nx4313), .B1 (nx4367)) ;
    inv01 ix4368 (.Y (nx4369), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_10)) ;
    oai32 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix503 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .A0 (
          nx4371), .A1 (RST), .A2 (nx7947), .B0 (nx4317), .B1 (nx4367)) ;
    inv01 ix4370 (.Y (nx4371), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_11)) ;
    oai32 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix513 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .A0 (
          nx4373), .A1 (RST), .A2 (nx7947), .B0 (nx4321), .B1 (nx4367)) ;
    inv01 ix4372 (.Y (nx4373), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_12)) ;
    oai32 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix523 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .A0 (
          nx4375), .A1 (RST), .A2 (nx7949), .B0 (nx4325), .B1 (nx4367)) ;
    inv01 ix4374 (.Y (nx4375), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_13)) ;
    oai32 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix533 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .A0 (
          nx4377), .A1 (RST), .A2 (nx7949), .B0 (nx4329), .B1 (nx4379)) ;
    inv01 ix4376 (.Y (nx4377), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_14)) ;
    inv01 ix4378 (.Y (nx4379), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566)) ;
    oai32 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix543 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .A0 (
          nx4381), .A1 (RST), .A2 (nx7949), .B0 (nx4333), .B1 (nx4379)) ;
    inv01 ix4380 (.Y (nx4381), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_15)) ;
    oai32 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix553 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .A0 (
          nx4383), .A1 (RST), .A2 (nx7949), .B0 (nx4337), .B1 (nx4379)) ;
    inv01 ix4382 (.Y (nx4383), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_16)) ;
    nand02_2x CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix633 (.Y (
              nx4365), .A0 (nx7361), .A1 (nx7949)) ;
    nand02_2x CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix635 (.Y (
              nx4367), .A0 (nx7361), .A1 (nx7949)) ;
    oai32 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix393 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .A0 (
          nx4385), .A1 (RST), .A2 (nx7951), .B0 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_nx384), .B1 (nx4387)) ;
    inv01 ix4384 (.Y (nx4385), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_0)) ;
    oai32 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix403 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .A0 (
          nx4389), .A1 (RST), .A2 (nx7951), .B0 (nx4205), .B1 (nx4387)) ;
    inv01 ix4388 (.Y (nx4389), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_1)) ;
    oai32 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix413 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .A0 (
          nx4391), .A1 (RST), .A2 (nx7951), .B0 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx387), .B1 (nx4387)) ;
    inv01 ix4390 (.Y (nx4391), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_2)) ;
    oai32 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix423 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .A0 (
          nx4393), .A1 (RST), .A2 (nx7951), .B0 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx399), .B1 (nx4387)) ;
    inv01 ix4392 (.Y (nx4393), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_3)) ;
    oai32 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix433 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .A0 (
          nx4395), .A1 (RST), .A2 (nx7951), .B0 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx409), .B1 (nx4387)) ;
    inv01 ix4394 (.Y (nx4395), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_4)) ;
    oai32 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix443 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .A0 (
          nx4397), .A1 (RST), .A2 (nx7951), .B0 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx419), .B1 (nx4387)) ;
    inv01 ix4396 (.Y (nx4397), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_5)) ;
    oai32 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix453 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .A0 (
          nx4399), .A1 (RST), .A2 (nx7951), .B0 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx429), .B1 (nx4387)) ;
    inv01 ix4398 (.Y (nx4399), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_6)) ;
    oai32 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix463 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .A0 (
          nx4401), .A1 (RST), .A2 (nx7953), .B0 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx439), .B1 (nx4403)) ;
    inv01 ix4400 (.Y (nx4401), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_7)) ;
    oai32 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix473 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .A0 (
          nx4405), .A1 (RST), .A2 (nx7953), .B0 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx449), .B1 (nx4403)) ;
    inv01 ix4404 (.Y (nx4405), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_8)) ;
    oai32 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix483 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .A0 (
          nx4407), .A1 (RST), .A2 (nx7953), .B0 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx469), .B1 (nx4403)) ;
    inv01 ix4406 (.Y (nx4407), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_9)) ;
    oai32 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix493 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .A0 (
          nx4409), .A1 (RST), .A2 (nx7953), .B0 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx477), .B1 (nx4403)) ;
    inv01 ix4408 (.Y (nx4409), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_10)) ;
    oai32 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix503 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .A0 (
          nx4411), .A1 (RST), .A2 (nx7953), .B0 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx485), .B1 (nx4403)) ;
    inv01 ix4410 (.Y (nx4411), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_11)) ;
    oai32 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix513 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .A0 (
          nx4413), .A1 (RST), .A2 (nx7953), .B0 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx493), .B1 (nx4403)) ;
    inv01 ix4412 (.Y (nx4413), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_12)) ;
    oai32 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix523 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .A0 (
          nx4415), .A1 (RST), .A2 (nx7953), .B0 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx501), .B1 (nx4403)) ;
    inv01 ix4414 (.Y (nx4415), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_13)) ;
    oai32 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix533 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .A0 (
          nx4417), .A1 (RST), .A2 (nx7955), .B0 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx509), .B1 (nx4419)) ;
    inv01 ix4416 (.Y (nx4417), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_14)) ;
    inv01 ix4418 (.Y (nx4419), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566)) ;
    oai32 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix543 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .A0 (
          nx4421), .A1 (RST), .A2 (nx7955), .B0 (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_nx517), .B1 (nx4419)) ;
    inv01 ix4420 (.Y (nx4421), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_15)) ;
    oai32 CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix553 (.Y (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .A0 (
          nx4423), .A1 (RST), .A2 (nx7955), .B0 (nx4221), .B1 (nx4419)) ;
    inv01 ix4422 (.Y (nx4423), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_16)) ;
    nand02_2x CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix633 (.Y (
              nx4387), .A0 (nx7361), .A1 (nx7955)) ;
    nand02_2x CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix635 (.Y (
              nx4403), .A0 (nx7361), .A1 (nx7955)) ;
    mux21 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix404 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx403), .A0 (nx4425), .A1 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_2), .S0 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx395)) ;
    inv01 ix4424 (.Y (nx4425), .A (CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx391)) ;
    mux21 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix414 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx413), .A0 (nx4427), .A1 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_3), .S0 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx405)) ;
    inv01 ix4426 (.Y (nx4427), .A (CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx403)) ;
    mux21 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix424 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx423), .A0 (nx4429), .A1 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_4), .S0 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx415)) ;
    inv01 ix4428 (.Y (nx4429), .A (CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx413)) ;
    mux21 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix434 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx433), .A0 (nx4431), .A1 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_5), .S0 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx425)) ;
    inv01 ix4430 (.Y (nx4431), .A (CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx423)) ;
    mux21 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix444 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx443), .A0 (nx4433), .A1 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_6), .S0 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx435)) ;
    inv01 ix4432 (.Y (nx4433), .A (CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx433)) ;
    mux21 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix454 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx453), .A0 (nx4435), .A1 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_7), .S0 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx445)) ;
    inv01 ix4434 (.Y (nx4435), .A (CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx443)) ;
    mux21 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix462 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx461), .A0 (nx4437), .A1 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_8), .S0 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx455)) ;
    inv01 ix4436 (.Y (nx4437), .A (CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx453)) ;
    mux21 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix468 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx467), .A0 (nx4439), .A1 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_9), .S0 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx463)) ;
    inv01 ix4438 (.Y (nx4439), .A (CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx461)) ;
    mux21 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix476 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx475), .A0 (nx4441), .A1 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_10), .S0 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx471)) ;
    inv01 ix4440 (.Y (nx4441), .A (CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx467)) ;
    mux21 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix484 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx483), .A0 (nx4443), .A1 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_11), .S0 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx479)) ;
    inv01 ix4442 (.Y (nx4443), .A (CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx475)) ;
    mux21 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix492 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx491), .A0 (nx4445), .A1 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_12), .S0 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx487)) ;
    inv01 ix4444 (.Y (nx4445), .A (CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx483)) ;
    mux21 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix500 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx499), .A0 (nx4447), .A1 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_13), .S0 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx495)) ;
    inv01 ix4446 (.Y (nx4447), .A (CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx491)) ;
    mux21 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix508 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx507), .A0 (nx4449), .A1 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_14), .S0 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx503)) ;
    inv01 ix4448 (.Y (nx4449), .A (CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx499)) ;
    mux21 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix516 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx515), .A0 (nx4451), .A1 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_15), .S0 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx511)) ;
    inv01 ix4450 (.Y (nx4451), .A (CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx507)) ;
    mux21 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix161 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_1), .A0 (nx4453), .A1 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx379), .S0 (nx7959)) ;
    inv01 ix4452 (.Y (nx4453), .A (CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_1)) ;
    mux21 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix181 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_2), .A0 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx387), .A1 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx389), .S0 (nx7959)) ;
    mux21 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix201 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_3), .A0 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx399), .A1 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx401), .S0 (nx7959)) ;
    mux21 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix221 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_4), .A0 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx409), .A1 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx411), .S0 (nx7959)) ;
    mux21 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix241 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_5), .A0 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx419), .A1 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx421), .S0 (nx7959)) ;
    mux21 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix261 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_6), .A0 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx429), .A1 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx431), .S0 (nx7959)) ;
    mux21 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix281 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_7), .A0 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx439), .A1 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx441), .S0 (nx7959)) ;
    mux21 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix301 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_8), .A0 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx449), .A1 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx451), .S0 (nx7961)) ;
    mux21 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix321 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_9), .A0 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx469), .A1 (nx4455), .S0 (nx7961)) ;
    inv01 ix4454 (.Y (nx4455), .A (CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx316)) ;
    mux21 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix341 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_10), .A0 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx477), .A1 (nx4457), .S0 (nx7961)) ;
    inv01 ix4456 (.Y (nx4457), .A (CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx336)) ;
    mux21 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix361 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_11), .A0 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx485), .A1 (nx4459), .S0 (nx7961)) ;
    inv01 ix4458 (.Y (nx4459), .A (CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx356)) ;
    mux21 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix381 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_12), .A0 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx493), .A1 (nx4461), .S0 (nx7961)) ;
    inv01 ix4460 (.Y (nx4461), .A (CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx376)) ;
    mux21 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix401 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_13), .A0 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx501), .A1 (nx4463), .S0 (nx7961)) ;
    inv01 ix4462 (.Y (nx4463), .A (CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx396)) ;
    mux21 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix421 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_14), .A0 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx509), .A1 (nx4465), .S0 (nx7961)) ;
    inv01 ix4464 (.Y (nx4465), .A (CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx416)) ;
    mux21 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix441 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_15), .A0 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx517), .A1 (nx4467), .S0 (nx7963)) ;
    inv01 ix4466 (.Y (nx4467), .A (CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx436)) ;
    mux21 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_ix461 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_16), .A0 (nx4469), 
          .A1 (nx4471), .S0 (nx7963)) ;
    inv01 ix4468 (.Y (nx4469), .A (CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothP_16)
          ) ;
    inv01 ix4470 (.Y (nx4471), .A (CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx456)) ;
    nor02_2x CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix81 (.Y (
             CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_nx80), .A0 (Instr), .A1 (
             nx7313)) ;
    nor02_2x CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix319 (.Y (
             CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642), .A0 (
             CALCULATOR_Start_dup_1235), .A1 (
             CALCULATOR_CalculatingBooth_dup_1224)) ;
    nor02_2x CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix85 (.Y (
             CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_0), .A0 (
             nx7973), .A1 (nx4473)) ;
    inv01 ix4472 (.Y (nx4473), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_1)) ;
    mux21 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix125 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_1), .A0 (
          nx4475), .A1 (nx4477), .S0 (nx7973)) ;
    inv01 ix4474 (.Y (nx4475), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_2)) ;
    inv01 ix4476 (.Y (nx4477), .A (CacheWindow_3__0__0)) ;
    mux21 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix133 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_2), .A0 (
          nx4479), .A1 (nx4481), .S0 (nx7973)) ;
    inv01 ix4478 (.Y (nx4479), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_3)) ;
    inv01 ix4480 (.Y (nx4481), .A (CacheWindow_3__0__1)) ;
    mux21 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix141 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_3), .A0 (
          nx4483), .A1 (nx4485), .S0 (nx7973)) ;
    inv01 ix4482 (.Y (nx4483), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_4)) ;
    inv01 ix4484 (.Y (nx4485), .A (CacheWindow_3__0__2)) ;
    mux21 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix149 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_4), .A0 (
          nx4487), .A1 (nx4489), .S0 (nx7973)) ;
    inv01 ix4486 (.Y (nx4487), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_5)) ;
    inv01 ix4488 (.Y (nx4489), .A (CacheWindow_3__0__3)) ;
    mux21 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix157 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_5), .A0 (
          nx4491), .A1 (nx4493), .S0 (nx7973)) ;
    inv01 ix4490 (.Y (nx4491), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_6)) ;
    inv01 ix4492 (.Y (nx4493), .A (CacheWindow_3__0__4)) ;
    mux21 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix165 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_6), .A0 (
          nx4495), .A1 (nx4497), .S0 (nx7973)) ;
    inv01 ix4494 (.Y (nx4495), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_7)) ;
    inv01 ix4496 (.Y (nx4497), .A (CacheWindow_3__0__5)) ;
    mux21 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix173 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_7), .A0 (
          nx4499), .A1 (nx4501), .S0 (nx7975)) ;
    inv01 ix4498 (.Y (nx4499), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_8)) ;
    inv01 ix4500 (.Y (nx4501), .A (CacheWindow_3__0__6)) ;
    mux21 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix181 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_8), .A0 (
          nx4503), .A1 (nx4505), .S0 (nx7975)) ;
    inv01 ix4502 (.Y (nx4503), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_9)) ;
    inv01 ix4504 (.Y (nx4505), .A (CacheWindow_3__0__7)) ;
    nor02_2x CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix89 (.Y (
             CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_9), .A0 (
             nx7975), .A1 (nx4507)) ;
    inv01 ix4506 (.Y (nx4507), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_10)) ;
    nor02_2x CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix93 (.Y (
             CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_10), .A0 (
             nx7975), .A1 (nx4509)) ;
    inv01 ix4508 (.Y (nx4509), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_11)) ;
    nor02_2x CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix97 (.Y (
             CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_11), .A0 (
             nx7975), .A1 (nx4511)) ;
    inv01 ix4510 (.Y (nx4511), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_12)) ;
    nor02_2x CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix101 (.Y (
             CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_12), .A0 (
             nx7975), .A1 (nx4513)) ;
    inv01 ix4512 (.Y (nx4513), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_13)) ;
    nor02_2x CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix105 (.Y (
             CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_13), .A0 (
             nx7975), .A1 (nx4515)) ;
    inv01 ix4514 (.Y (nx4515), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_14)) ;
    nor02_2x CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix109 (.Y (
             CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_14), .A0 (
             nx7977), .A1 (nx4517)) ;
    inv01 ix4516 (.Y (nx4517), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_15)) ;
    nor02_2x CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix113 (.Y (
             CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_15), .A0 (
             nx7977), .A1 (nx4519)) ;
    inv01 ix4518 (.Y (nx4519), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_16)) ;
    nor02_2x CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix117 (.Y (
             CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_16), .A0 (
             nx7977), .A1 (nx4519)) ;
    mux21 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix189 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothOperand_0), .A0 (nx4521), .A1 (
          nx4523), .S0 (nx7965)) ;
    inv01 ix4520 (.Y (nx4521), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_0)) ;
    inv01 ix4522 (.Y (nx4523), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_0)) ;
    mux21 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix197 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothOperand_1), .A0 (nx4525), .A1 (
          nx4527), .S0 (nx7965)) ;
    inv01 ix4524 (.Y (nx4525), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_1)) ;
    inv01 ix4526 (.Y (nx4527), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_1)) ;
    mux21 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix205 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothOperand_2), .A0 (nx4529), .A1 (
          nx4531), .S0 (nx7965)) ;
    inv01 ix4528 (.Y (nx4529), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_2)) ;
    inv01 ix4530 (.Y (nx4531), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_2)) ;
    mux21 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix213 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothOperand_3), .A0 (nx4533), .A1 (
          nx4535), .S0 (nx7965)) ;
    inv01 ix4532 (.Y (nx4533), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_3)) ;
    inv01 ix4534 (.Y (nx4535), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_3)) ;
    mux21 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix221 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothOperand_4), .A0 (nx4537), .A1 (
          nx4539), .S0 (nx7965)) ;
    inv01 ix4536 (.Y (nx4537), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_4)) ;
    inv01 ix4538 (.Y (nx4539), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_4)) ;
    mux21 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix229 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothOperand_5), .A0 (nx4541), .A1 (
          nx4543), .S0 (nx7967)) ;
    inv01 ix4540 (.Y (nx4541), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_5)) ;
    inv01 ix4542 (.Y (nx4543), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_5)) ;
    mux21 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix237 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothOperand_6), .A0 (nx4545), .A1 (
          nx4547), .S0 (nx7967)) ;
    inv01 ix4544 (.Y (nx4545), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_6)) ;
    inv01 ix4546 (.Y (nx4547), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_6)) ;
    mux21 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix245 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothOperand_7), .A0 (nx4549), .A1 (
          nx4551), .S0 (nx7967)) ;
    inv01 ix4548 (.Y (nx4549), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_7)) ;
    inv01 ix4550 (.Y (nx4551), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_7)) ;
    mux21 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix253 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothOperand_8), .A0 (nx4553), .A1 (
          nx4555), .S0 (nx7967)) ;
    inv01 ix4552 (.Y (nx4553), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_8)) ;
    inv01 ix4554 (.Y (nx4555), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_8)) ;
    mux21 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix261 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothOperand_9), .A0 (nx4557), .A1 (
          nx4559), .S0 (nx7967)) ;
    inv01 ix4556 (.Y (nx4557), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_9)) ;
    inv01 ix4558 (.Y (nx4559), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_9)) ;
    mux21 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix269 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothOperand_10), .A0 (nx4561), .A1 (
          nx4563), .S0 (nx7967)) ;
    inv01 ix4560 (.Y (nx4561), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_10)) ;
    inv01 ix4562 (.Y (nx4563), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_10)) ;
    mux21 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix277 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothOperand_11), .A0 (nx4565), .A1 (
          nx4567), .S0 (nx7967)) ;
    inv01 ix4564 (.Y (nx4565), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_11)) ;
    inv01 ix4566 (.Y (nx4567), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_11)) ;
    mux21 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix285 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothOperand_12), .A0 (nx4569), .A1 (
          nx4571), .S0 (nx7969)) ;
    inv01 ix4568 (.Y (nx4569), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_12)) ;
    inv01 ix4570 (.Y (nx4571), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_12)) ;
    mux21 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix293 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothOperand_13), .A0 (nx4573), .A1 (
          nx4575), .S0 (nx7969)) ;
    inv01 ix4572 (.Y (nx4573), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_13)) ;
    inv01 ix4574 (.Y (nx4575), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_13)) ;
    mux21 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix301 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothOperand_14), .A0 (nx4577), .A1 (
          nx4579), .S0 (nx7969)) ;
    inv01 ix4576 (.Y (nx4577), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_14)) ;
    inv01 ix4578 (.Y (nx4579), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_14)) ;
    mux21 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix309 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothOperand_15), .A0 (nx4581), .A1 (
          nx4583), .S0 (nx7969)) ;
    inv01 ix4580 (.Y (nx4581), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_15)) ;
    inv01 ix4582 (.Y (nx4583), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_15)) ;
    mux21 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix317 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BoothOperand_16), .A0 (nx4585), .A1 (
          nx4587), .S0 (nx7969)) ;
    inv01 ix4584 (.Y (nx4585), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_16)) ;
    inv01 ix4586 (.Y (nx4587), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_16)) ;
    xnor2 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix321 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_AddPToBoothOperand), .A0 (nx7969), .A1 (
          nx4453)) ;
    oai32 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix393 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .A0 (
          nx8569), .A1 (RST), .A2 (nx7979), .B0 (nx4523), .B1 (nx4591)) ;
    oai32 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix403 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .A0 (
          nx8569), .A1 (RST), .A2 (nx7979), .B0 (nx4527), .B1 (nx4591)) ;
    oai32 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix413 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .A0 (
          nx8569), .A1 (RST), .A2 (nx7979), .B0 (nx4531), .B1 (nx4591)) ;
    oai32 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix423 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .A0 (
          nx8569), .A1 (RST), .A2 (nx7979), .B0 (nx4535), .B1 (nx4591)) ;
    oai32 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix433 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .A0 (
          nx8569), .A1 (RST), .A2 (nx7979), .B0 (nx4539), .B1 (nx4591)) ;
    oai32 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix443 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .A0 (
          nx8569), .A1 (RST), .A2 (nx7979), .B0 (nx4543), .B1 (nx4591)) ;
    oai32 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix453 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .A0 (
          nx8569), .A1 (RST), .A2 (nx7981), .B0 (nx4547), .B1 (nx4591)) ;
    oai32 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix463 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .A0 (
          nx8571), .A1 (RST), .A2 (nx7981), .B0 (nx4551), .B1 (nx4593)) ;
    oai32 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix473 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .A0 (
          nx8571), .A1 (RST), .A2 (nx7981), .B0 (nx4555), .B1 (nx4593)) ;
    oai32 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix483 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .A0 (
          nx4595), .A1 (RST), .A2 (nx7981), .B0 (nx4559), .B1 (nx4593)) ;
    inv01 ix4594 (.Y (nx4595), .A (CacheFilter_3__0__0)) ;
    oai32 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix493 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .A0 (
          nx4597), .A1 (RST), .A2 (nx7981), .B0 (nx4563), .B1 (nx4593)) ;
    inv01 ix4596 (.Y (nx4597), .A (CacheFilter_3__0__1)) ;
    oai32 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix503 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .A0 (
          nx4599), .A1 (RST), .A2 (nx7981), .B0 (nx4567), .B1 (nx4593)) ;
    inv01 ix4598 (.Y (nx4599), .A (CacheFilter_3__0__2)) ;
    oai32 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix513 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .A0 (
          nx4601), .A1 (RST), .A2 (nx7981), .B0 (nx4571), .B1 (nx4593)) ;
    inv01 ix4600 (.Y (nx4601), .A (CacheFilter_3__0__3)) ;
    oai32 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix523 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .A0 (
          nx4603), .A1 (RST), .A2 (nx7983), .B0 (nx4575), .B1 (nx4593)) ;
    inv01 ix4602 (.Y (nx4603), .A (CacheFilter_3__0__4)) ;
    oai32 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix533 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .A0 (
          nx4605), .A1 (RST), .A2 (nx7983), .B0 (nx4579), .B1 (nx4607)) ;
    inv01 ix4604 (.Y (nx4605), .A (CacheFilter_3__0__5)) ;
    inv01 ix4606 (.Y (nx4607), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566)) ;
    oai32 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix543 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .A0 (
          nx4609), .A1 (RST), .A2 (nx7983), .B0 (nx4583), .B1 (nx4607)) ;
    inv01 ix4608 (.Y (nx4609), .A (CacheFilter_3__0__6)) ;
    oai32 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix553 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .A0 (
          nx4611), .A1 (RST), .A2 (nx7983), .B0 (nx4587), .B1 (nx4607)) ;
    inv01 ix4610 (.Y (nx4611), .A (CacheFilter_3__0__7)) ;
    nand02_2x CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix633 (.Y (
              nx4591), .A0 (nx7363), .A1 (nx7983)) ;
    nand02_2x CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix635 (.Y (
              nx4593), .A0 (nx7363), .A1 (nx7983)) ;
    oai32 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix393 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .A0 (
          nx8571), .A1 (RST), .A2 (nx7985), .B0 (nx4521), .B1 (nx4613)) ;
    oai32 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix403 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .A0 (
          nx8571), .A1 (RST), .A2 (nx7985), .B0 (nx4525), .B1 (nx4613)) ;
    oai32 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix413 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .A0 (
          nx8571), .A1 (RST), .A2 (nx7985), .B0 (nx4529), .B1 (nx4613)) ;
    oai32 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix423 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .A0 (
          nx8571), .A1 (RST), .A2 (nx7985), .B0 (nx4533), .B1 (nx4613)) ;
    oai32 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix433 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .A0 (
          nx8571), .A1 (RST), .A2 (nx7985), .B0 (nx4537), .B1 (nx4613)) ;
    oai32 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix443 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .A0 (
          nx8573), .A1 (RST), .A2 (nx7985), .B0 (nx4541), .B1 (nx4613)) ;
    oai32 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix453 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .A0 (
          nx8573), .A1 (RST), .A2 (nx7987), .B0 (nx4545), .B1 (nx4613)) ;
    oai32 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix463 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .A0 (
          nx8573), .A1 (RST), .A2 (nx7987), .B0 (nx4549), .B1 (nx4615)) ;
    oai32 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix473 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .A0 (
          nx8573), .A1 (RST), .A2 (nx7987), .B0 (nx4553), .B1 (nx4615)) ;
    oai32 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix483 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .A0 (
          nx4595), .A1 (RST), .A2 (nx7987), .B0 (nx4557), .B1 (nx4615)) ;
    oai32 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix493 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .A0 (
          nx4617), .A1 (RST), .A2 (nx7987), .B0 (nx4561), .B1 (nx4615)) ;
    inv01 ix4616 (.Y (nx4617), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_10)) ;
    oai32 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix503 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .A0 (
          nx4619), .A1 (RST), .A2 (nx7987), .B0 (nx4565), .B1 (nx4615)) ;
    inv01 ix4618 (.Y (nx4619), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_11)) ;
    oai32 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix513 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .A0 (
          nx4621), .A1 (RST), .A2 (nx7987), .B0 (nx4569), .B1 (nx4615)) ;
    inv01 ix4620 (.Y (nx4621), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_12)) ;
    oai32 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix523 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .A0 (
          nx4623), .A1 (RST), .A2 (nx7989), .B0 (nx4573), .B1 (nx4615)) ;
    inv01 ix4622 (.Y (nx4623), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_13)) ;
    oai32 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix533 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .A0 (
          nx4625), .A1 (RST), .A2 (nx7989), .B0 (nx4577), .B1 (nx4627)) ;
    inv01 ix4624 (.Y (nx4625), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_14)) ;
    inv01 ix4626 (.Y (nx4627), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566)) ;
    oai32 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix543 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .A0 (
          nx4629), .A1 (RST), .A2 (nx7989), .B0 (nx4581), .B1 (nx4627)) ;
    inv01 ix4628 (.Y (nx4629), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_15)) ;
    oai32 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix553 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .A0 (
          nx4631), .A1 (RST), .A2 (nx7989), .B0 (nx4585), .B1 (nx4627)) ;
    inv01 ix4630 (.Y (nx4631), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_16)) ;
    nand02_2x CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix633 (.Y (
              nx4613), .A0 (nx7363), .A1 (nx7989)) ;
    nand02_2x CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix635 (.Y (
              nx4615), .A0 (nx7363), .A1 (nx7989)) ;
    oai32 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix393 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .A0 (
          nx4633), .A1 (RST), .A2 (nx7991), .B0 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_nx384), .B1 (nx4635)) ;
    inv01 ix4632 (.Y (nx4633), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_0)) ;
    oai32 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix403 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .A0 (
          nx4637), .A1 (RST), .A2 (nx7991), .B0 (nx4453), .B1 (nx4635)) ;
    inv01 ix4636 (.Y (nx4637), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_1)) ;
    oai32 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix413 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .A0 (
          nx4639), .A1 (RST), .A2 (nx7991), .B0 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx387), .B1 (nx4635)) ;
    inv01 ix4638 (.Y (nx4639), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_2)) ;
    oai32 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix423 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .A0 (
          nx4641), .A1 (RST), .A2 (nx7991), .B0 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx399), .B1 (nx4635)) ;
    inv01 ix4640 (.Y (nx4641), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_3)) ;
    oai32 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix433 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .A0 (
          nx4643), .A1 (RST), .A2 (nx7991), .B0 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx409), .B1 (nx4635)) ;
    inv01 ix4642 (.Y (nx4643), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_4)) ;
    oai32 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix443 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .A0 (
          nx4645), .A1 (RST), .A2 (nx7991), .B0 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx419), .B1 (nx4635)) ;
    inv01 ix4644 (.Y (nx4645), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_5)) ;
    oai32 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix453 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .A0 (
          nx4647), .A1 (RST), .A2 (nx7991), .B0 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx429), .B1 (nx4635)) ;
    inv01 ix4646 (.Y (nx4647), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_6)) ;
    oai32 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix463 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .A0 (
          nx4649), .A1 (RST), .A2 (nx7993), .B0 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx439), .B1 (nx4651)) ;
    inv01 ix4648 (.Y (nx4649), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_7)) ;
    oai32 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix473 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .A0 (
          nx4653), .A1 (RST), .A2 (nx7993), .B0 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx449), .B1 (nx4651)) ;
    inv01 ix4652 (.Y (nx4653), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_8)) ;
    oai32 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix483 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .A0 (
          nx4655), .A1 (RST), .A2 (nx7993), .B0 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx469), .B1 (nx4651)) ;
    inv01 ix4654 (.Y (nx4655), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_9)) ;
    oai32 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix493 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .A0 (
          nx4657), .A1 (RST), .A2 (nx7993), .B0 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx477), .B1 (nx4651)) ;
    inv01 ix4656 (.Y (nx4657), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_10)) ;
    oai32 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix503 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .A0 (
          nx4659), .A1 (RST), .A2 (nx7993), .B0 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx485), .B1 (nx4651)) ;
    inv01 ix4658 (.Y (nx4659), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_11)) ;
    oai32 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix513 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .A0 (
          nx4661), .A1 (RST), .A2 (nx7993), .B0 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx493), .B1 (nx4651)) ;
    inv01 ix4660 (.Y (nx4661), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_12)) ;
    oai32 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix523 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .A0 (
          nx4663), .A1 (RST), .A2 (nx7993), .B0 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx501), .B1 (nx4651)) ;
    inv01 ix4662 (.Y (nx4663), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_13)) ;
    oai32 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix533 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .A0 (
          nx4665), .A1 (RST), .A2 (nx7995), .B0 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx509), .B1 (nx4667)) ;
    inv01 ix4664 (.Y (nx4665), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_14)) ;
    inv01 ix4666 (.Y (nx4667), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566)) ;
    oai32 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix543 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .A0 (
          nx4669), .A1 (RST), .A2 (nx7995), .B0 (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_nx517), .B1 (nx4667)) ;
    inv01 ix4668 (.Y (nx4669), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_15)) ;
    oai32 CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix553 (.Y (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .A0 (
          nx4671), .A1 (RST), .A2 (nx7995), .B0 (nx4469), .B1 (nx4667)) ;
    inv01 ix4670 (.Y (nx4671), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_16)) ;
    nand02_2x CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix633 (.Y (
              nx4635), .A0 (nx7363), .A1 (nx7995)) ;
    nand02_2x CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix635 (.Y (
              nx4651), .A0 (nx7363), .A1 (nx7995)) ;
    mux21 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix404 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx403), .A0 (nx4673), .A1 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_2), .S0 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx395)) ;
    inv01 ix4672 (.Y (nx4673), .A (CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx391)) ;
    mux21 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix414 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx413), .A0 (nx4675), .A1 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_3), .S0 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx405)) ;
    inv01 ix4674 (.Y (nx4675), .A (CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx403)) ;
    mux21 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix424 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx423), .A0 (nx4677), .A1 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_4), .S0 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx415)) ;
    inv01 ix4676 (.Y (nx4677), .A (CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx413)) ;
    mux21 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix434 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx433), .A0 (nx4679), .A1 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_5), .S0 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx425)) ;
    inv01 ix4678 (.Y (nx4679), .A (CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx423)) ;
    mux21 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix444 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx443), .A0 (nx4681), .A1 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_6), .S0 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx435)) ;
    inv01 ix4680 (.Y (nx4681), .A (CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx433)) ;
    mux21 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix454 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx453), .A0 (nx4683), .A1 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_7), .S0 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx445)) ;
    inv01 ix4682 (.Y (nx4683), .A (CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx443)) ;
    mux21 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix462 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx461), .A0 (nx4685), .A1 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_8), .S0 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx455)) ;
    inv01 ix4684 (.Y (nx4685), .A (CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx453)) ;
    mux21 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix468 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx467), .A0 (nx4687), .A1 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_9), .S0 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx463)) ;
    inv01 ix4686 (.Y (nx4687), .A (CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx461)) ;
    mux21 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix476 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx475), .A0 (nx4689), .A1 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_10), .S0 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx471)) ;
    inv01 ix4688 (.Y (nx4689), .A (CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx467)) ;
    mux21 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix484 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx483), .A0 (nx4691), .A1 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_11), .S0 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx479)) ;
    inv01 ix4690 (.Y (nx4691), .A (CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx475)) ;
    mux21 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix492 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx491), .A0 (nx4693), .A1 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_12), .S0 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx487)) ;
    inv01 ix4692 (.Y (nx4693), .A (CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx483)) ;
    mux21 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix500 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx499), .A0 (nx4695), .A1 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_13), .S0 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx495)) ;
    inv01 ix4694 (.Y (nx4695), .A (CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx491)) ;
    mux21 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix508 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx507), .A0 (nx4697), .A1 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_14), .S0 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx503)) ;
    inv01 ix4696 (.Y (nx4697), .A (CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx499)) ;
    mux21 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix516 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx515), .A0 (nx4699), .A1 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_15), .S0 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx511)) ;
    inv01 ix4698 (.Y (nx4699), .A (CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx507)) ;
    mux21 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix161 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_1), .A0 (nx4701), .A1 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx379), .S0 (nx7999)) ;
    inv01 ix4700 (.Y (nx4701), .A (CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_1)) ;
    mux21 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix181 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_2), .A0 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx387), .A1 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx389), .S0 (nx7999)) ;
    mux21 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix201 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_3), .A0 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx399), .A1 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx401), .S0 (nx7999)) ;
    mux21 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix221 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_4), .A0 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx409), .A1 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx411), .S0 (nx7999)) ;
    mux21 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix241 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_5), .A0 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx419), .A1 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx421), .S0 (nx7999)) ;
    mux21 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix261 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_6), .A0 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx429), .A1 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx431), .S0 (nx7999)) ;
    mux21 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix281 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_7), .A0 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx439), .A1 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx441), .S0 (nx7999)) ;
    mux21 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix301 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_8), .A0 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx449), .A1 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx451), .S0 (nx8001)) ;
    mux21 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix321 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_9), .A0 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx469), .A1 (nx4703), .S0 (nx8001)) ;
    inv01 ix4702 (.Y (nx4703), .A (CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx316)) ;
    mux21 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix341 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_10), .A0 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx477), .A1 (nx4705), .S0 (nx8001)) ;
    inv01 ix4704 (.Y (nx4705), .A (CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx336)) ;
    mux21 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix361 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_11), .A0 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx485), .A1 (nx4707), .S0 (nx8001)) ;
    inv01 ix4706 (.Y (nx4707), .A (CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx356)) ;
    mux21 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix381 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_12), .A0 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx493), .A1 (nx4709), .S0 (nx8001)) ;
    inv01 ix4708 (.Y (nx4709), .A (CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx376)) ;
    mux21 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix401 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_13), .A0 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx501), .A1 (nx4711), .S0 (nx8001)) ;
    inv01 ix4710 (.Y (nx4711), .A (CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx396)) ;
    mux21 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix421 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_14), .A0 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx509), .A1 (nx4713), .S0 (nx8001)) ;
    inv01 ix4712 (.Y (nx4713), .A (CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx416)) ;
    mux21 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix441 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_15), .A0 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx517), .A1 (nx4715), .S0 (nx8003)) ;
    inv01 ix4714 (.Y (nx4715), .A (CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx436)) ;
    mux21 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_ix461 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_16), .A0 (nx4717), 
          .A1 (nx4719), .S0 (nx8003)) ;
    inv01 ix4716 (.Y (nx4717), .A (CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothP_16)
          ) ;
    inv01 ix4718 (.Y (nx4719), .A (CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx456)) ;
    nor02_2x CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix81 (.Y (
             CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_nx80), .A0 (Instr), .A1 (
             nx7313)) ;
    nor02_2x CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix319 (.Y (
             CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642), .A0 (
             CALCULATOR_Start_dup_1248), .A1 (
             CALCULATOR_CalculatingBooth_dup_1224)) ;
    nor02_2x CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix85 (.Y (
             CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_0), .A0 (
             nx8013), .A1 (nx4721)) ;
    inv01 ix4720 (.Y (nx4721), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_1)) ;
    mux21 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix125 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_1), .A0 (
          nx4723), .A1 (nx4725), .S0 (nx8013)) ;
    inv01 ix4722 (.Y (nx4723), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_2)) ;
    inv01 ix4724 (.Y (nx4725), .A (CacheWindow_3__1__0)) ;
    mux21 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix133 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_2), .A0 (
          nx4727), .A1 (nx4729), .S0 (nx8013)) ;
    inv01 ix4726 (.Y (nx4727), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_3)) ;
    inv01 ix4728 (.Y (nx4729), .A (CacheWindow_3__1__1)) ;
    mux21 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix141 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_3), .A0 (
          nx4731), .A1 (nx4733), .S0 (nx8013)) ;
    inv01 ix4730 (.Y (nx4731), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_4)) ;
    inv01 ix4732 (.Y (nx4733), .A (CacheWindow_3__1__2)) ;
    mux21 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix149 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_4), .A0 (
          nx4735), .A1 (nx4737), .S0 (nx8013)) ;
    inv01 ix4734 (.Y (nx4735), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_5)) ;
    inv01 ix4736 (.Y (nx4737), .A (CacheWindow_3__1__3)) ;
    mux21 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix157 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_5), .A0 (
          nx4739), .A1 (nx4741), .S0 (nx8013)) ;
    inv01 ix4738 (.Y (nx4739), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_6)) ;
    inv01 ix4740 (.Y (nx4741), .A (CacheWindow_3__1__4)) ;
    mux21 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix165 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_6), .A0 (
          nx4743), .A1 (nx4745), .S0 (nx8013)) ;
    inv01 ix4742 (.Y (nx4743), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_7)) ;
    inv01 ix4744 (.Y (nx4745), .A (CacheWindow_3__1__5)) ;
    mux21 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix173 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_7), .A0 (
          nx4747), .A1 (nx4749), .S0 (nx8015)) ;
    inv01 ix4746 (.Y (nx4747), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_8)) ;
    inv01 ix4748 (.Y (nx4749), .A (CacheWindow_3__1__6)) ;
    mux21 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix181 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_8), .A0 (
          nx4751), .A1 (nx4753), .S0 (nx8015)) ;
    inv01 ix4750 (.Y (nx4751), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_9)) ;
    inv01 ix4752 (.Y (nx4753), .A (CacheWindow_3__1__7)) ;
    nor02_2x CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix89 (.Y (
             CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_9), .A0 (
             nx8015), .A1 (nx4755)) ;
    inv01 ix4754 (.Y (nx4755), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_10)) ;
    nor02_2x CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix93 (.Y (
             CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_10), .A0 (
             nx8015), .A1 (nx4757)) ;
    inv01 ix4756 (.Y (nx4757), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_11)) ;
    nor02_2x CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix97 (.Y (
             CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_11), .A0 (
             nx8015), .A1 (nx4759)) ;
    inv01 ix4758 (.Y (nx4759), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_12)) ;
    nor02_2x CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix101 (.Y (
             CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_12), .A0 (
             nx8015), .A1 (nx4761)) ;
    inv01 ix4760 (.Y (nx4761), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_13)) ;
    nor02_2x CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix105 (.Y (
             CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_13), .A0 (
             nx8015), .A1 (nx4763)) ;
    inv01 ix4762 (.Y (nx4763), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_14)) ;
    nor02_2x CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix109 (.Y (
             CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_14), .A0 (
             nx8017), .A1 (nx4765)) ;
    inv01 ix4764 (.Y (nx4765), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_15)) ;
    nor02_2x CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix113 (.Y (
             CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_15), .A0 (
             nx8017), .A1 (nx4767)) ;
    inv01 ix4766 (.Y (nx4767), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_16)) ;
    nor02_2x CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix117 (.Y (
             CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_16), .A0 (
             nx8017), .A1 (nx4767)) ;
    mux21 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix189 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothOperand_0), .A0 (nx4769), .A1 (
          nx4771), .S0 (nx8005)) ;
    inv01 ix4768 (.Y (nx4769), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_0)) ;
    inv01 ix4770 (.Y (nx4771), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_0)) ;
    mux21 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix197 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothOperand_1), .A0 (nx4773), .A1 (
          nx4775), .S0 (nx8005)) ;
    inv01 ix4772 (.Y (nx4773), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_1)) ;
    inv01 ix4774 (.Y (nx4775), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_1)) ;
    mux21 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix205 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothOperand_2), .A0 (nx4777), .A1 (
          nx4779), .S0 (nx8005)) ;
    inv01 ix4776 (.Y (nx4777), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_2)) ;
    inv01 ix4778 (.Y (nx4779), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_2)) ;
    mux21 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix213 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothOperand_3), .A0 (nx4781), .A1 (
          nx4783), .S0 (nx8005)) ;
    inv01 ix4780 (.Y (nx4781), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_3)) ;
    inv01 ix4782 (.Y (nx4783), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_3)) ;
    mux21 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix221 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothOperand_4), .A0 (nx4785), .A1 (
          nx4787), .S0 (nx8005)) ;
    inv01 ix4784 (.Y (nx4785), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_4)) ;
    inv01 ix4786 (.Y (nx4787), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_4)) ;
    mux21 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix229 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothOperand_5), .A0 (nx4789), .A1 (
          nx4791), .S0 (nx8007)) ;
    inv01 ix4788 (.Y (nx4789), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_5)) ;
    inv01 ix4790 (.Y (nx4791), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_5)) ;
    mux21 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix237 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothOperand_6), .A0 (nx4793), .A1 (
          nx4795), .S0 (nx8007)) ;
    inv01 ix4792 (.Y (nx4793), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_6)) ;
    inv01 ix4794 (.Y (nx4795), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_6)) ;
    mux21 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix245 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothOperand_7), .A0 (nx4797), .A1 (
          nx4799), .S0 (nx8007)) ;
    inv01 ix4796 (.Y (nx4797), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_7)) ;
    inv01 ix4798 (.Y (nx4799), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_7)) ;
    mux21 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix253 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothOperand_8), .A0 (nx4801), .A1 (
          nx4803), .S0 (nx8007)) ;
    inv01 ix4800 (.Y (nx4801), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_8)) ;
    inv01 ix4802 (.Y (nx4803), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_8)) ;
    mux21 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix261 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothOperand_9), .A0 (nx4805), .A1 (
          nx4807), .S0 (nx8007)) ;
    inv01 ix4804 (.Y (nx4805), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_9)) ;
    inv01 ix4806 (.Y (nx4807), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_9)) ;
    mux21 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix269 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothOperand_10), .A0 (nx4809), .A1 (
          nx4811), .S0 (nx8007)) ;
    inv01 ix4808 (.Y (nx4809), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_10)) ;
    inv01 ix4810 (.Y (nx4811), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_10)) ;
    mux21 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix277 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothOperand_11), .A0 (nx4813), .A1 (
          nx4815), .S0 (nx8007)) ;
    inv01 ix4812 (.Y (nx4813), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_11)) ;
    inv01 ix4814 (.Y (nx4815), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_11)) ;
    mux21 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix285 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothOperand_12), .A0 (nx4817), .A1 (
          nx4819), .S0 (nx8009)) ;
    inv01 ix4816 (.Y (nx4817), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_12)) ;
    inv01 ix4818 (.Y (nx4819), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_12)) ;
    mux21 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix293 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothOperand_13), .A0 (nx4821), .A1 (
          nx4823), .S0 (nx8009)) ;
    inv01 ix4820 (.Y (nx4821), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_13)) ;
    inv01 ix4822 (.Y (nx4823), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_13)) ;
    mux21 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix301 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothOperand_14), .A0 (nx4825), .A1 (
          nx4827), .S0 (nx8009)) ;
    inv01 ix4824 (.Y (nx4825), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_14)) ;
    inv01 ix4826 (.Y (nx4827), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_14)) ;
    mux21 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix309 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothOperand_15), .A0 (nx4829), .A1 (
          nx4831), .S0 (nx8009)) ;
    inv01 ix4828 (.Y (nx4829), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_15)) ;
    inv01 ix4830 (.Y (nx4831), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_15)) ;
    mux21 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix317 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BoothOperand_16), .A0 (nx4833), .A1 (
          nx4835), .S0 (nx8009)) ;
    inv01 ix4832 (.Y (nx4833), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_16)) ;
    inv01 ix4834 (.Y (nx4835), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_16)) ;
    xnor2 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix321 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_AddPToBoothOperand), .A0 (nx8009), .A1 (
          nx4701)) ;
    oai32 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix393 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .A0 (
          nx8575), .A1 (RST), .A2 (nx8019), .B0 (nx4771), .B1 (nx4839)) ;
    oai32 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix403 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .A0 (
          nx8575), .A1 (RST), .A2 (nx8019), .B0 (nx4775), .B1 (nx4839)) ;
    oai32 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix413 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .A0 (
          nx8575), .A1 (RST), .A2 (nx8019), .B0 (nx4779), .B1 (nx4839)) ;
    oai32 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix423 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .A0 (
          nx8575), .A1 (RST), .A2 (nx8019), .B0 (nx4783), .B1 (nx4839)) ;
    oai32 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix433 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .A0 (
          nx8575), .A1 (RST), .A2 (nx8019), .B0 (nx4787), .B1 (nx4839)) ;
    oai32 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix443 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .A0 (
          nx8575), .A1 (RST), .A2 (nx8019), .B0 (nx4791), .B1 (nx4839)) ;
    oai32 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix453 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .A0 (
          nx8575), .A1 (RST), .A2 (nx8021), .B0 (nx4795), .B1 (nx4839)) ;
    oai32 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix463 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .A0 (
          nx8577), .A1 (RST), .A2 (nx8021), .B0 (nx4799), .B1 (nx4841)) ;
    oai32 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix473 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .A0 (
          nx8577), .A1 (RST), .A2 (nx8021), .B0 (nx4803), .B1 (nx4841)) ;
    oai32 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix483 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .A0 (
          nx4843), .A1 (RST), .A2 (nx8021), .B0 (nx4807), .B1 (nx4841)) ;
    inv01 ix4842 (.Y (nx4843), .A (CacheFilter_3__1__0)) ;
    oai32 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix493 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .A0 (
          nx4845), .A1 (RST), .A2 (nx8021), .B0 (nx4811), .B1 (nx4841)) ;
    inv01 ix4844 (.Y (nx4845), .A (CacheFilter_3__1__1)) ;
    oai32 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix503 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .A0 (
          nx4847), .A1 (RST), .A2 (nx8021), .B0 (nx4815), .B1 (nx4841)) ;
    inv01 ix4846 (.Y (nx4847), .A (CacheFilter_3__1__2)) ;
    oai32 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix513 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .A0 (
          nx4849), .A1 (RST), .A2 (nx8021), .B0 (nx4819), .B1 (nx4841)) ;
    inv01 ix4848 (.Y (nx4849), .A (CacheFilter_3__1__3)) ;
    oai32 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix523 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .A0 (
          nx4851), .A1 (RST), .A2 (nx8023), .B0 (nx4823), .B1 (nx4841)) ;
    inv01 ix4850 (.Y (nx4851), .A (CacheFilter_3__1__4)) ;
    oai32 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix533 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .A0 (
          nx4853), .A1 (RST), .A2 (nx8023), .B0 (nx4827), .B1 (nx4855)) ;
    inv01 ix4852 (.Y (nx4853), .A (CacheFilter_3__1__5)) ;
    inv01 ix4854 (.Y (nx4855), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566)) ;
    oai32 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix543 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .A0 (
          nx4857), .A1 (RST), .A2 (nx8023), .B0 (nx4831), .B1 (nx4855)) ;
    inv01 ix4856 (.Y (nx4857), .A (CacheFilter_3__1__6)) ;
    oai32 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix553 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .A0 (
          nx4859), .A1 (RST), .A2 (nx8023), .B0 (nx4835), .B1 (nx4855)) ;
    inv01 ix4858 (.Y (nx4859), .A (CacheFilter_3__1__7)) ;
    nand02_2x CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix633 (.Y (
              nx4839), .A0 (nx7363), .A1 (nx8023)) ;
    nand02_2x CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix635 (.Y (
              nx4841), .A0 (nx7365), .A1 (nx8023)) ;
    oai32 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix393 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .A0 (
          nx8577), .A1 (RST), .A2 (nx8025), .B0 (nx4769), .B1 (nx4861)) ;
    oai32 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix403 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .A0 (
          nx8577), .A1 (RST), .A2 (nx8025), .B0 (nx4773), .B1 (nx4861)) ;
    oai32 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix413 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .A0 (
          nx8577), .A1 (RST), .A2 (nx8025), .B0 (nx4777), .B1 (nx4861)) ;
    oai32 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix423 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .A0 (
          nx8577), .A1 (RST), .A2 (nx8025), .B0 (nx4781), .B1 (nx4861)) ;
    oai32 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix433 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .A0 (
          nx8577), .A1 (RST), .A2 (nx8025), .B0 (nx4785), .B1 (nx4861)) ;
    oai32 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix443 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .A0 (
          nx8579), .A1 (RST), .A2 (nx8025), .B0 (nx4789), .B1 (nx4861)) ;
    oai32 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix453 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .A0 (
          nx8579), .A1 (RST), .A2 (nx8027), .B0 (nx4793), .B1 (nx4861)) ;
    oai32 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix463 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .A0 (
          nx8579), .A1 (RST), .A2 (nx8027), .B0 (nx4797), .B1 (nx4863)) ;
    oai32 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix473 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .A0 (
          nx8579), .A1 (RST), .A2 (nx8027), .B0 (nx4801), .B1 (nx4863)) ;
    oai32 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix483 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .A0 (
          nx4843), .A1 (RST), .A2 (nx8027), .B0 (nx4805), .B1 (nx4863)) ;
    oai32 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix493 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .A0 (
          nx4865), .A1 (RST), .A2 (nx8027), .B0 (nx4809), .B1 (nx4863)) ;
    inv01 ix4864 (.Y (nx4865), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_10)) ;
    oai32 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix503 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .A0 (
          nx4867), .A1 (RST), .A2 (nx8027), .B0 (nx4813), .B1 (nx4863)) ;
    inv01 ix4866 (.Y (nx4867), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_11)) ;
    oai32 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix513 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .A0 (
          nx4869), .A1 (RST), .A2 (nx8027), .B0 (nx4817), .B1 (nx4863)) ;
    inv01 ix4868 (.Y (nx4869), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_12)) ;
    oai32 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix523 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .A0 (
          nx4871), .A1 (RST), .A2 (nx8029), .B0 (nx4821), .B1 (nx4863)) ;
    inv01 ix4870 (.Y (nx4871), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_13)) ;
    oai32 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix533 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .A0 (
          nx4873), .A1 (RST), .A2 (nx8029), .B0 (nx4825), .B1 (nx4875)) ;
    inv01 ix4872 (.Y (nx4873), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_14)) ;
    inv01 ix4874 (.Y (nx4875), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566)) ;
    oai32 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix543 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .A0 (
          nx4877), .A1 (RST), .A2 (nx8029), .B0 (nx4829), .B1 (nx4875)) ;
    inv01 ix4876 (.Y (nx4877), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_15)) ;
    oai32 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix553 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .A0 (
          nx4879), .A1 (RST), .A2 (nx8029), .B0 (nx4833), .B1 (nx4875)) ;
    inv01 ix4878 (.Y (nx4879), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_16)) ;
    nand02_2x CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix633 (.Y (
              nx4861), .A0 (nx7365), .A1 (nx8029)) ;
    nand02_2x CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix635 (.Y (
              nx4863), .A0 (nx7365), .A1 (nx8029)) ;
    oai32 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix393 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .A0 (
          nx4881), .A1 (RST), .A2 (nx8031), .B0 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_nx384), .B1 (nx4883)) ;
    inv01 ix4880 (.Y (nx4881), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_0)) ;
    oai32 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix403 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .A0 (
          nx4885), .A1 (RST), .A2 (nx8031), .B0 (nx4701), .B1 (nx4883)) ;
    inv01 ix4884 (.Y (nx4885), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_1)) ;
    oai32 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix413 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .A0 (
          nx4887), .A1 (RST), .A2 (nx8031), .B0 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx387), .B1 (nx4883)) ;
    inv01 ix4886 (.Y (nx4887), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_2)) ;
    oai32 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix423 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .A0 (
          nx4889), .A1 (RST), .A2 (nx8031), .B0 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx399), .B1 (nx4883)) ;
    inv01 ix4888 (.Y (nx4889), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_3)) ;
    oai32 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix433 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .A0 (
          nx4891), .A1 (RST), .A2 (nx8031), .B0 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx409), .B1 (nx4883)) ;
    inv01 ix4890 (.Y (nx4891), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_4)) ;
    oai32 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix443 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .A0 (
          nx4893), .A1 (RST), .A2 (nx8031), .B0 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx419), .B1 (nx4883)) ;
    inv01 ix4892 (.Y (nx4893), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_5)) ;
    oai32 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix453 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .A0 (
          nx4895), .A1 (RST), .A2 (nx8031), .B0 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx429), .B1 (nx4883)) ;
    inv01 ix4894 (.Y (nx4895), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_6)) ;
    oai32 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix463 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .A0 (
          nx4897), .A1 (RST), .A2 (nx8033), .B0 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx439), .B1 (nx4899)) ;
    inv01 ix4896 (.Y (nx4897), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_7)) ;
    oai32 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix473 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .A0 (
          nx4901), .A1 (RST), .A2 (nx8033), .B0 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx449), .B1 (nx4899)) ;
    inv01 ix4900 (.Y (nx4901), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_8)) ;
    oai32 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix483 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .A0 (
          nx4903), .A1 (RST), .A2 (nx8033), .B0 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx469), .B1 (nx4899)) ;
    inv01 ix4902 (.Y (nx4903), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_9)) ;
    oai32 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix493 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .A0 (
          nx4905), .A1 (RST), .A2 (nx8033), .B0 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx477), .B1 (nx4899)) ;
    inv01 ix4904 (.Y (nx4905), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_10)) ;
    oai32 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix503 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .A0 (
          nx4907), .A1 (RST), .A2 (nx8033), .B0 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx485), .B1 (nx4899)) ;
    inv01 ix4906 (.Y (nx4907), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_11)) ;
    oai32 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix513 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .A0 (
          nx4909), .A1 (RST), .A2 (nx8033), .B0 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx493), .B1 (nx4899)) ;
    inv01 ix4908 (.Y (nx4909), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_12)) ;
    oai32 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix523 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .A0 (
          nx4911), .A1 (RST), .A2 (nx8033), .B0 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx501), .B1 (nx4899)) ;
    inv01 ix4910 (.Y (nx4911), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_13)) ;
    oai32 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix533 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .A0 (
          nx4913), .A1 (RST), .A2 (nx8035), .B0 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx509), .B1 (nx4915)) ;
    inv01 ix4912 (.Y (nx4913), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_14)) ;
    inv01 ix4914 (.Y (nx4915), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566)) ;
    oai32 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix543 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .A0 (
          nx4917), .A1 (RST), .A2 (nx8035), .B0 (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_nx517), .B1 (nx4915)) ;
    inv01 ix4916 (.Y (nx4917), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_15)) ;
    oai32 CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix553 (.Y (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .A0 (
          nx4919), .A1 (RST), .A2 (nx8035), .B0 (nx4717), .B1 (nx4915)) ;
    inv01 ix4918 (.Y (nx4919), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_16)) ;
    nand02_2x CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix633 (.Y (
              nx4883), .A0 (nx7365), .A1 (nx8035)) ;
    nand02_2x CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix635 (.Y (
              nx4899), .A0 (nx7365), .A1 (nx8035)) ;
    mux21 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix404 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx403), .A0 (nx4921), .A1 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_2), .S0 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx395)) ;
    inv01 ix4920 (.Y (nx4921), .A (CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx391)) ;
    mux21 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix414 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx413), .A0 (nx4923), .A1 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_3), .S0 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx405)) ;
    inv01 ix4922 (.Y (nx4923), .A (CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx403)) ;
    mux21 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix424 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx423), .A0 (nx4925), .A1 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_4), .S0 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx415)) ;
    inv01 ix4924 (.Y (nx4925), .A (CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx413)) ;
    mux21 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix434 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx433), .A0 (nx4927), .A1 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_5), .S0 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx425)) ;
    inv01 ix4926 (.Y (nx4927), .A (CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx423)) ;
    mux21 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix444 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx443), .A0 (nx4929), .A1 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_6), .S0 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx435)) ;
    inv01 ix4928 (.Y (nx4929), .A (CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx433)) ;
    mux21 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix454 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx453), .A0 (nx4931), .A1 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_7), .S0 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx445)) ;
    inv01 ix4930 (.Y (nx4931), .A (CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx443)) ;
    mux21 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix462 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx461), .A0 (nx4933), .A1 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_8), .S0 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx455)) ;
    inv01 ix4932 (.Y (nx4933), .A (CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx453)) ;
    mux21 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix468 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx467), .A0 (nx4935), .A1 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_9), .S0 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx463)) ;
    inv01 ix4934 (.Y (nx4935), .A (CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx461)) ;
    mux21 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix476 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx475), .A0 (nx4937), .A1 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_10), .S0 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx471)) ;
    inv01 ix4936 (.Y (nx4937), .A (CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx467)) ;
    mux21 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix484 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx483), .A0 (nx4939), .A1 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_11), .S0 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx479)) ;
    inv01 ix4938 (.Y (nx4939), .A (CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx475)) ;
    mux21 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix492 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx491), .A0 (nx4941), .A1 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_12), .S0 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx487)) ;
    inv01 ix4940 (.Y (nx4941), .A (CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx483)) ;
    mux21 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix500 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx499), .A0 (nx4943), .A1 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_13), .S0 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx495)) ;
    inv01 ix4942 (.Y (nx4943), .A (CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx491)) ;
    mux21 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix508 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx507), .A0 (nx4945), .A1 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_14), .S0 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx503)) ;
    inv01 ix4944 (.Y (nx4945), .A (CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx499)) ;
    mux21 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix516 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx515), .A0 (nx4947), .A1 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_15), .S0 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx511)) ;
    inv01 ix4946 (.Y (nx4947), .A (CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx507)) ;
    mux21 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix161 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_1), .A0 (nx4949), .A1 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx379), .S0 (nx8039)) ;
    inv01 ix4948 (.Y (nx4949), .A (CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_1)) ;
    mux21 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix181 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_2), .A0 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx387), .A1 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx389), .S0 (nx8039)) ;
    mux21 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix201 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_3), .A0 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx399), .A1 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx401), .S0 (nx8039)) ;
    mux21 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix221 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_4), .A0 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx409), .A1 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx411), .S0 (nx8039)) ;
    mux21 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix241 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_5), .A0 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx419), .A1 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx421), .S0 (nx8039)) ;
    mux21 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix261 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_6), .A0 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx429), .A1 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx431), .S0 (nx8039)) ;
    mux21 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix281 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_7), .A0 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx439), .A1 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx441), .S0 (nx8039)) ;
    mux21 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix301 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_8), .A0 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx449), .A1 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx451), .S0 (nx8041)) ;
    mux21 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix321 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_9), .A0 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx469), .A1 (nx4951), .S0 (nx8041)) ;
    inv01 ix4950 (.Y (nx4951), .A (CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx316)) ;
    mux21 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix341 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_10), .A0 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx477), .A1 (nx4953), .S0 (nx8041)) ;
    inv01 ix4952 (.Y (nx4953), .A (CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx336)) ;
    mux21 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix361 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_11), .A0 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx485), .A1 (nx4955), .S0 (nx8041)) ;
    inv01 ix4954 (.Y (nx4955), .A (CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx356)) ;
    mux21 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix381 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_12), .A0 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx493), .A1 (nx4957), .S0 (nx8041)) ;
    inv01 ix4956 (.Y (nx4957), .A (CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx376)) ;
    mux21 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix401 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_13), .A0 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx501), .A1 (nx4959), .S0 (nx8041)) ;
    inv01 ix4958 (.Y (nx4959), .A (CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx396)) ;
    mux21 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix421 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_14), .A0 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx509), .A1 (nx4961), .S0 (nx8041)) ;
    inv01 ix4960 (.Y (nx4961), .A (CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx416)) ;
    mux21 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix441 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_15), .A0 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx517), .A1 (nx4963), .S0 (nx8043)) ;
    inv01 ix4962 (.Y (nx4963), .A (CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx436)) ;
    mux21 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_ix461 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_16), .A0 (nx4965), 
          .A1 (nx4967), .S0 (nx8043)) ;
    inv01 ix4964 (.Y (nx4965), .A (CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothP_16)
          ) ;
    inv01 ix4966 (.Y (nx4967), .A (CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx456)) ;
    nor02_2x CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix81 (.Y (
             CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_nx80), .A0 (Instr), .A1 (
             nx7313)) ;
    nor02_2x CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix319 (.Y (
             CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642), .A0 (
             CALCULATOR_Start_dup_1261), .A1 (
             CALCULATOR_CalculatingBooth_dup_1224)) ;
    nor02_2x CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix85 (.Y (
             CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_0), .A0 (
             nx8053), .A1 (nx4969)) ;
    inv01 ix4968 (.Y (nx4969), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_1)) ;
    mux21 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix125 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_1), .A0 (
          nx4971), .A1 (nx4973), .S0 (nx8053)) ;
    inv01 ix4970 (.Y (nx4971), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_2)) ;
    inv01 ix4972 (.Y (nx4973), .A (CacheWindow_3__2__0)) ;
    mux21 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix133 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_2), .A0 (
          nx4975), .A1 (nx4977), .S0 (nx8053)) ;
    inv01 ix4974 (.Y (nx4975), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_3)) ;
    inv01 ix4976 (.Y (nx4977), .A (CacheWindow_3__2__1)) ;
    mux21 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix141 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_3), .A0 (
          nx4979), .A1 (nx4981), .S0 (nx8053)) ;
    inv01 ix4978 (.Y (nx4979), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_4)) ;
    inv01 ix4980 (.Y (nx4981), .A (CacheWindow_3__2__2)) ;
    mux21 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix149 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_4), .A0 (
          nx4983), .A1 (nx4985), .S0 (nx8053)) ;
    inv01 ix4982 (.Y (nx4983), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_5)) ;
    inv01 ix4984 (.Y (nx4985), .A (CacheWindow_3__2__3)) ;
    mux21 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix157 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_5), .A0 (
          nx4987), .A1 (nx4989), .S0 (nx8053)) ;
    inv01 ix4986 (.Y (nx4987), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_6)) ;
    inv01 ix4988 (.Y (nx4989), .A (CacheWindow_3__2__4)) ;
    mux21 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix165 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_6), .A0 (
          nx4991), .A1 (nx4993), .S0 (nx8053)) ;
    inv01 ix4990 (.Y (nx4991), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_7)) ;
    inv01 ix4992 (.Y (nx4993), .A (CacheWindow_3__2__5)) ;
    mux21 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix173 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_7), .A0 (
          nx4995), .A1 (nx4997), .S0 (nx8055)) ;
    inv01 ix4994 (.Y (nx4995), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_8)) ;
    inv01 ix4996 (.Y (nx4997), .A (CacheWindow_3__2__6)) ;
    mux21 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix181 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_8), .A0 (
          nx4999), .A1 (nx5001), .S0 (nx8055)) ;
    inv01 ix4998 (.Y (nx4999), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_9)) ;
    inv01 ix5000 (.Y (nx5001), .A (CacheWindow_3__2__7)) ;
    nor02_2x CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix89 (.Y (
             CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_9), .A0 (
             nx8055), .A1 (nx5003)) ;
    inv01 ix5002 (.Y (nx5003), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_10)) ;
    nor02_2x CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix93 (.Y (
             CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_10), .A0 (
             nx8055), .A1 (nx5005)) ;
    inv01 ix5004 (.Y (nx5005), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_11)) ;
    nor02_2x CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix97 (.Y (
             CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_11), .A0 (
             nx8055), .A1 (nx5007)) ;
    inv01 ix5006 (.Y (nx5007), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_12)) ;
    nor02_2x CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix101 (.Y (
             CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_12), .A0 (
             nx8055), .A1 (nx5009)) ;
    inv01 ix5008 (.Y (nx5009), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_13)) ;
    nor02_2x CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix105 (.Y (
             CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_13), .A0 (
             nx8055), .A1 (nx5011)) ;
    inv01 ix5010 (.Y (nx5011), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_14)) ;
    nor02_2x CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix109 (.Y (
             CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_14), .A0 (
             nx8057), .A1 (nx5013)) ;
    inv01 ix5012 (.Y (nx5013), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_15)) ;
    nor02_2x CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix113 (.Y (
             CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_15), .A0 (
             nx8057), .A1 (nx5015)) ;
    inv01 ix5014 (.Y (nx5015), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_16)) ;
    nor02_2x CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix117 (.Y (
             CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_16), .A0 (
             nx8057), .A1 (nx5015)) ;
    mux21 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix189 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothOperand_0), .A0 (nx5017), .A1 (
          nx5019), .S0 (nx8045)) ;
    inv01 ix5016 (.Y (nx5017), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_0)) ;
    inv01 ix5018 (.Y (nx5019), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_0)) ;
    mux21 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix197 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothOperand_1), .A0 (nx5021), .A1 (
          nx5023), .S0 (nx8045)) ;
    inv01 ix5020 (.Y (nx5021), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_1)) ;
    inv01 ix5022 (.Y (nx5023), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_1)) ;
    mux21 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix205 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothOperand_2), .A0 (nx5025), .A1 (
          nx5027), .S0 (nx8045)) ;
    inv01 ix5024 (.Y (nx5025), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_2)) ;
    inv01 ix5026 (.Y (nx5027), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_2)) ;
    mux21 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix213 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothOperand_3), .A0 (nx5029), .A1 (
          nx5031), .S0 (nx8045)) ;
    inv01 ix5028 (.Y (nx5029), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_3)) ;
    inv01 ix5030 (.Y (nx5031), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_3)) ;
    mux21 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix221 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothOperand_4), .A0 (nx5033), .A1 (
          nx5035), .S0 (nx8045)) ;
    inv01 ix5032 (.Y (nx5033), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_4)) ;
    inv01 ix5034 (.Y (nx5035), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_4)) ;
    mux21 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix229 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothOperand_5), .A0 (nx5037), .A1 (
          nx5039), .S0 (nx8047)) ;
    inv01 ix5036 (.Y (nx5037), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_5)) ;
    inv01 ix5038 (.Y (nx5039), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_5)) ;
    mux21 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix237 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothOperand_6), .A0 (nx5041), .A1 (
          nx5043), .S0 (nx8047)) ;
    inv01 ix5040 (.Y (nx5041), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_6)) ;
    inv01 ix5042 (.Y (nx5043), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_6)) ;
    mux21 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix245 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothOperand_7), .A0 (nx5045), .A1 (
          nx5047), .S0 (nx8047)) ;
    inv01 ix5044 (.Y (nx5045), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_7)) ;
    inv01 ix5046 (.Y (nx5047), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_7)) ;
    mux21 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix253 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothOperand_8), .A0 (nx5049), .A1 (
          nx5051), .S0 (nx8047)) ;
    inv01 ix5048 (.Y (nx5049), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_8)) ;
    inv01 ix5050 (.Y (nx5051), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_8)) ;
    mux21 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix261 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothOperand_9), .A0 (nx5053), .A1 (
          nx5055), .S0 (nx8047)) ;
    inv01 ix5052 (.Y (nx5053), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_9)) ;
    inv01 ix5054 (.Y (nx5055), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_9)) ;
    mux21 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix269 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothOperand_10), .A0 (nx5057), .A1 (
          nx5059), .S0 (nx8047)) ;
    inv01 ix5056 (.Y (nx5057), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_10)) ;
    inv01 ix5058 (.Y (nx5059), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_10)) ;
    mux21 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix277 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothOperand_11), .A0 (nx5061), .A1 (
          nx5063), .S0 (nx8047)) ;
    inv01 ix5060 (.Y (nx5061), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_11)) ;
    inv01 ix5062 (.Y (nx5063), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_11)) ;
    mux21 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix285 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothOperand_12), .A0 (nx5065), .A1 (
          nx5067), .S0 (nx8049)) ;
    inv01 ix5064 (.Y (nx5065), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_12)) ;
    inv01 ix5066 (.Y (nx5067), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_12)) ;
    mux21 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix293 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothOperand_13), .A0 (nx5069), .A1 (
          nx5071), .S0 (nx8049)) ;
    inv01 ix5068 (.Y (nx5069), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_13)) ;
    inv01 ix5070 (.Y (nx5071), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_13)) ;
    mux21 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix301 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothOperand_14), .A0 (nx5073), .A1 (
          nx5075), .S0 (nx8049)) ;
    inv01 ix5072 (.Y (nx5073), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_14)) ;
    inv01 ix5074 (.Y (nx5075), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_14)) ;
    mux21 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix309 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothOperand_15), .A0 (nx5077), .A1 (
          nx5079), .S0 (nx8049)) ;
    inv01 ix5076 (.Y (nx5077), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_15)) ;
    inv01 ix5078 (.Y (nx5079), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_15)) ;
    mux21 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix317 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BoothOperand_16), .A0 (nx5081), .A1 (
          nx5083), .S0 (nx8049)) ;
    inv01 ix5080 (.Y (nx5081), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_16)) ;
    inv01 ix5082 (.Y (nx5083), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_16)) ;
    xnor2 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix321 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_AddPToBoothOperand), .A0 (nx8049), .A1 (
          nx4949)) ;
    oai32 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix393 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .A0 (
          nx8581), .A1 (RST), .A2 (nx8059), .B0 (nx5019), .B1 (nx5087)) ;
    oai32 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix403 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .A0 (
          nx8581), .A1 (RST), .A2 (nx8059), .B0 (nx5023), .B1 (nx5087)) ;
    oai32 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix413 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .A0 (
          nx8581), .A1 (RST), .A2 (nx8059), .B0 (nx5027), .B1 (nx5087)) ;
    oai32 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix423 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .A0 (
          nx8581), .A1 (RST), .A2 (nx8059), .B0 (nx5031), .B1 (nx5087)) ;
    oai32 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix433 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .A0 (
          nx8581), .A1 (RST), .A2 (nx8059), .B0 (nx5035), .B1 (nx5087)) ;
    oai32 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix443 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .A0 (
          nx8581), .A1 (RST), .A2 (nx8059), .B0 (nx5039), .B1 (nx5087)) ;
    oai32 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix453 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .A0 (
          nx8581), .A1 (RST), .A2 (nx8061), .B0 (nx5043), .B1 (nx5087)) ;
    oai32 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix463 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .A0 (
          nx8583), .A1 (RST), .A2 (nx8061), .B0 (nx5047), .B1 (nx5089)) ;
    oai32 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix473 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .A0 (
          nx8583), .A1 (RST), .A2 (nx8061), .B0 (nx5051), .B1 (nx5089)) ;
    oai32 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix483 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .A0 (
          nx5091), .A1 (RST), .A2 (nx8061), .B0 (nx5055), .B1 (nx5089)) ;
    inv01 ix5090 (.Y (nx5091), .A (CacheFilter_3__2__0)) ;
    oai32 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix493 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .A0 (
          nx5093), .A1 (RST), .A2 (nx8061), .B0 (nx5059), .B1 (nx5089)) ;
    inv01 ix5092 (.Y (nx5093), .A (CacheFilter_3__2__1)) ;
    oai32 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix503 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .A0 (
          nx5095), .A1 (RST), .A2 (nx8061), .B0 (nx5063), .B1 (nx5089)) ;
    inv01 ix5094 (.Y (nx5095), .A (CacheFilter_3__2__2)) ;
    oai32 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix513 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .A0 (
          nx5097), .A1 (RST), .A2 (nx8061), .B0 (nx5067), .B1 (nx5089)) ;
    inv01 ix5096 (.Y (nx5097), .A (CacheFilter_3__2__3)) ;
    oai32 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix523 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .A0 (
          nx5099), .A1 (RST), .A2 (nx8063), .B0 (nx5071), .B1 (nx5089)) ;
    inv01 ix5098 (.Y (nx5099), .A (CacheFilter_3__2__4)) ;
    oai32 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix533 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .A0 (
          nx5101), .A1 (RST), .A2 (nx8063), .B0 (nx5075), .B1 (nx5103)) ;
    inv01 ix5100 (.Y (nx5101), .A (CacheFilter_3__2__5)) ;
    inv01 ix5102 (.Y (nx5103), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566)) ;
    oai32 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix543 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .A0 (
          nx5105), .A1 (RST), .A2 (nx8063), .B0 (nx5079), .B1 (nx5103)) ;
    inv01 ix5104 (.Y (nx5105), .A (CacheFilter_3__2__6)) ;
    oai32 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix553 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .A0 (
          nx5107), .A1 (RST), .A2 (nx8063), .B0 (nx5083), .B1 (nx5103)) ;
    inv01 ix5106 (.Y (nx5107), .A (CacheFilter_3__2__7)) ;
    nand02_2x CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix633 (.Y (
              nx5087), .A0 (nx7365), .A1 (nx8063)) ;
    nand02_2x CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix635 (.Y (
              nx5089), .A0 (nx7365), .A1 (nx8063)) ;
    oai32 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix393 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .A0 (
          nx8583), .A1 (RST), .A2 (nx8065), .B0 (nx5017), .B1 (nx5109)) ;
    oai32 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix403 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .A0 (
          nx8583), .A1 (RST), .A2 (nx8065), .B0 (nx5021), .B1 (nx5109)) ;
    oai32 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix413 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .A0 (
          nx8583), .A1 (RST), .A2 (nx8065), .B0 (nx5025), .B1 (nx5109)) ;
    oai32 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix423 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .A0 (
          nx8583), .A1 (RST), .A2 (nx8065), .B0 (nx5029), .B1 (nx5109)) ;
    oai32 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix433 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .A0 (
          nx8583), .A1 (RST), .A2 (nx8065), .B0 (nx5033), .B1 (nx5109)) ;
    oai32 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix443 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .A0 (
          nx8585), .A1 (RST), .A2 (nx8065), .B0 (nx5037), .B1 (nx5109)) ;
    oai32 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix453 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .A0 (
          nx8585), .A1 (RST), .A2 (nx8067), .B0 (nx5041), .B1 (nx5109)) ;
    oai32 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix463 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .A0 (
          nx8585), .A1 (RST), .A2 (nx8067), .B0 (nx5045), .B1 (nx5111)) ;
    oai32 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix473 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .A0 (
          nx8585), .A1 (RST), .A2 (nx8067), .B0 (nx5049), .B1 (nx5111)) ;
    oai32 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix483 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .A0 (
          nx5091), .A1 (RST), .A2 (nx8067), .B0 (nx5053), .B1 (nx5111)) ;
    oai32 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix493 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .A0 (
          nx5113), .A1 (RST), .A2 (nx8067), .B0 (nx5057), .B1 (nx5111)) ;
    inv01 ix5112 (.Y (nx5113), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_10)) ;
    oai32 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix503 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .A0 (
          nx5115), .A1 (RST), .A2 (nx8067), .B0 (nx5061), .B1 (nx5111)) ;
    inv01 ix5114 (.Y (nx5115), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_11)) ;
    oai32 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix513 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .A0 (
          nx5117), .A1 (RST), .A2 (nx8067), .B0 (nx5065), .B1 (nx5111)) ;
    inv01 ix5116 (.Y (nx5117), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_12)) ;
    oai32 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix523 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .A0 (
          nx5119), .A1 (RST), .A2 (nx8069), .B0 (nx5069), .B1 (nx5111)) ;
    inv01 ix5118 (.Y (nx5119), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_13)) ;
    oai32 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix533 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .A0 (
          nx5121), .A1 (RST), .A2 (nx8069), .B0 (nx5073), .B1 (nx5123)) ;
    inv01 ix5120 (.Y (nx5121), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_14)) ;
    inv01 ix5122 (.Y (nx5123), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566)) ;
    oai32 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix543 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .A0 (
          nx5125), .A1 (RST), .A2 (nx8069), .B0 (nx5077), .B1 (nx5123)) ;
    inv01 ix5124 (.Y (nx5125), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_15)) ;
    oai32 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix553 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .A0 (
          nx5127), .A1 (RST), .A2 (nx8069), .B0 (nx5081), .B1 (nx5123)) ;
    inv01 ix5126 (.Y (nx5127), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_16)) ;
    nand02_2x CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix633 (.Y (
              nx5109), .A0 (nx7367), .A1 (nx8069)) ;
    nand02_2x CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix635 (.Y (
              nx5111), .A0 (nx7367), .A1 (nx8069)) ;
    oai32 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix393 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .A0 (
          nx5129), .A1 (RST), .A2 (nx8071), .B0 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_nx384), .B1 (nx5131)) ;
    inv01 ix5128 (.Y (nx5129), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_0)) ;
    oai32 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix403 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .A0 (
          nx5133), .A1 (RST), .A2 (nx8071), .B0 (nx4949), .B1 (nx5131)) ;
    inv01 ix5132 (.Y (nx5133), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_1)) ;
    oai32 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix413 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .A0 (
          nx5135), .A1 (RST), .A2 (nx8071), .B0 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx387), .B1 (nx5131)) ;
    inv01 ix5134 (.Y (nx5135), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_2)) ;
    oai32 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix423 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .A0 (
          nx5137), .A1 (RST), .A2 (nx8071), .B0 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx399), .B1 (nx5131)) ;
    inv01 ix5136 (.Y (nx5137), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_3)) ;
    oai32 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix433 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .A0 (
          nx5139), .A1 (RST), .A2 (nx8071), .B0 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx409), .B1 (nx5131)) ;
    inv01 ix5138 (.Y (nx5139), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_4)) ;
    oai32 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix443 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .A0 (
          nx5141), .A1 (RST), .A2 (nx8071), .B0 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx419), .B1 (nx5131)) ;
    inv01 ix5140 (.Y (nx5141), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_5)) ;
    oai32 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix453 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .A0 (
          nx5143), .A1 (RST), .A2 (nx8071), .B0 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx429), .B1 (nx5131)) ;
    inv01 ix5142 (.Y (nx5143), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_6)) ;
    oai32 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix463 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .A0 (
          nx5145), .A1 (RST), .A2 (nx8073), .B0 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx439), .B1 (nx5147)) ;
    inv01 ix5144 (.Y (nx5145), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_7)) ;
    oai32 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix473 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .A0 (
          nx5149), .A1 (RST), .A2 (nx8073), .B0 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx449), .B1 (nx5147)) ;
    inv01 ix5148 (.Y (nx5149), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_8)) ;
    oai32 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix483 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .A0 (
          nx5151), .A1 (RST), .A2 (nx8073), .B0 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx469), .B1 (nx5147)) ;
    inv01 ix5150 (.Y (nx5151), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_9)) ;
    oai32 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix493 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .A0 (
          nx5153), .A1 (RST), .A2 (nx8073), .B0 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx477), .B1 (nx5147)) ;
    inv01 ix5152 (.Y (nx5153), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_10)) ;
    oai32 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix503 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .A0 (
          nx5155), .A1 (RST), .A2 (nx8073), .B0 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx485), .B1 (nx5147)) ;
    inv01 ix5154 (.Y (nx5155), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_11)) ;
    oai32 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix513 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .A0 (
          nx5157), .A1 (RST), .A2 (nx8073), .B0 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx493), .B1 (nx5147)) ;
    inv01 ix5156 (.Y (nx5157), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_12)) ;
    oai32 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix523 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .A0 (
          nx5159), .A1 (RST), .A2 (nx8073), .B0 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx501), .B1 (nx5147)) ;
    inv01 ix5158 (.Y (nx5159), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_13)) ;
    oai32 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix533 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .A0 (
          nx5161), .A1 (RST), .A2 (nx8075), .B0 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx509), .B1 (nx5163)) ;
    inv01 ix5160 (.Y (nx5161), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_14)) ;
    inv01 ix5162 (.Y (nx5163), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566)) ;
    oai32 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix543 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .A0 (
          nx5165), .A1 (RST), .A2 (nx8075), .B0 (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_nx517), .B1 (nx5163)) ;
    inv01 ix5164 (.Y (nx5165), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_15)) ;
    oai32 CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix553 (.Y (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .A0 (
          nx5167), .A1 (RST), .A2 (nx8075), .B0 (nx4965), .B1 (nx5163)) ;
    inv01 ix5166 (.Y (nx5167), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_16)) ;
    nand02_2x CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix633 (.Y (
              nx5131), .A0 (nx7367), .A1 (nx8075)) ;
    nand02_2x CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix635 (.Y (
              nx5147), .A0 (nx7367), .A1 (nx8075)) ;
    mux21 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix404 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx403), .A0 (nx5169), .A1 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_2), .S0 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx395)) ;
    inv01 ix5168 (.Y (nx5169), .A (CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx391)) ;
    mux21 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix414 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx413), .A0 (nx5171), .A1 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_3), .S0 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx405)) ;
    inv01 ix5170 (.Y (nx5171), .A (CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx403)) ;
    mux21 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix424 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx423), .A0 (nx5173), .A1 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_4), .S0 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx415)) ;
    inv01 ix5172 (.Y (nx5173), .A (CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx413)) ;
    mux21 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix434 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx433), .A0 (nx5175), .A1 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_5), .S0 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx425)) ;
    inv01 ix5174 (.Y (nx5175), .A (CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx423)) ;
    mux21 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix444 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx443), .A0 (nx5177), .A1 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_6), .S0 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx435)) ;
    inv01 ix5176 (.Y (nx5177), .A (CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx433)) ;
    mux21 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix454 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx453), .A0 (nx5179), .A1 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_7), .S0 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx445)) ;
    inv01 ix5178 (.Y (nx5179), .A (CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx443)) ;
    mux21 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix462 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx461), .A0 (nx5181), .A1 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_8), .S0 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx455)) ;
    inv01 ix5180 (.Y (nx5181), .A (CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx453)) ;
    mux21 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix468 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx467), .A0 (nx5183), .A1 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_9), .S0 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx463)) ;
    inv01 ix5182 (.Y (nx5183), .A (CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx461)) ;
    mux21 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix476 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx475), .A0 (nx5185), .A1 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_10), .S0 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx471)) ;
    inv01 ix5184 (.Y (nx5185), .A (CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx467)) ;
    mux21 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix484 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx483), .A0 (nx5187), .A1 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_11), .S0 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx479)) ;
    inv01 ix5186 (.Y (nx5187), .A (CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx475)) ;
    mux21 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix492 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx491), .A0 (nx5189), .A1 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_12), .S0 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx487)) ;
    inv01 ix5188 (.Y (nx5189), .A (CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx483)) ;
    mux21 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix500 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx499), .A0 (nx5191), .A1 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_13), .S0 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx495)) ;
    inv01 ix5190 (.Y (nx5191), .A (CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx491)) ;
    mux21 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix508 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx507), .A0 (nx5193), .A1 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_14), .S0 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx503)) ;
    inv01 ix5192 (.Y (nx5193), .A (CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx499)) ;
    mux21 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix516 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx515), .A0 (nx5195), .A1 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_15), .S0 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx511)) ;
    inv01 ix5194 (.Y (nx5195), .A (CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx507)) ;
    mux21 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix161 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_1), .A0 (nx5197), .A1 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx379), .S0 (nx8079)) ;
    inv01 ix5196 (.Y (nx5197), .A (CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_1)) ;
    mux21 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix181 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_2), .A0 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx387), .A1 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx389), .S0 (nx8079)) ;
    mux21 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix201 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_3), .A0 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx399), .A1 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx401), .S0 (nx8079)) ;
    mux21 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix221 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_4), .A0 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx409), .A1 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx411), .S0 (nx8079)) ;
    mux21 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix241 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_5), .A0 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx419), .A1 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx421), .S0 (nx8079)) ;
    mux21 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix261 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_6), .A0 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx429), .A1 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx431), .S0 (nx8079)) ;
    mux21 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix281 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_7), .A0 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx439), .A1 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx441), .S0 (nx8079)) ;
    mux21 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix301 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_8), .A0 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx449), .A1 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx451), .S0 (nx8081)) ;
    mux21 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix321 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_9), .A0 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx469), .A1 (nx5199), .S0 (nx8081)) ;
    inv01 ix5198 (.Y (nx5199), .A (CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx316)) ;
    mux21 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix341 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_10), .A0 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx477), .A1 (nx5201), .S0 (nx8081)) ;
    inv01 ix5200 (.Y (nx5201), .A (CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx336)) ;
    mux21 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix361 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_11), .A0 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx485), .A1 (nx5203), .S0 (nx8081)) ;
    inv01 ix5202 (.Y (nx5203), .A (CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx356)) ;
    mux21 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix381 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_12), .A0 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx493), .A1 (nx5205), .S0 (nx8081)) ;
    inv01 ix5204 (.Y (nx5205), .A (CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx376)) ;
    mux21 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix401 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_13), .A0 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx501), .A1 (nx5207), .S0 (nx8081)) ;
    inv01 ix5206 (.Y (nx5207), .A (CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx396)) ;
    mux21 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix421 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_14), .A0 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx509), .A1 (nx5209), .S0 (nx8081)) ;
    inv01 ix5208 (.Y (nx5209), .A (CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx416)) ;
    mux21 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix441 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_15), .A0 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx517), .A1 (nx5211), .S0 (nx8083)) ;
    inv01 ix5210 (.Y (nx5211), .A (CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx436)) ;
    mux21 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_ix461 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_16), .A0 (nx5213), 
          .A1 (nx5215), .S0 (nx8083)) ;
    inv01 ix5212 (.Y (nx5213), .A (CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothP_16)
          ) ;
    inv01 ix5214 (.Y (nx5215), .A (CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx456)) ;
    nor02_2x CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix81 (.Y (
             CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx80), .A0 (Instr), .A1 (
             nx7313)) ;
    nor02_2x CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix319 (.Y (
             CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642), .A0 (
             CALCULATOR_Start_dup_1274), .A1 (
             CALCULATOR_CalculatingBooth_dup_1224)) ;
    nor02_2x CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix85 (.Y (
             CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_0), .A0 (
             nx8093), .A1 (nx5217)) ;
    inv01 ix5216 (.Y (nx5217), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_1)) ;
    mux21 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix125 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_1), .A0 (
          nx5219), .A1 (nx5221), .S0 (nx8093)) ;
    inv01 ix5218 (.Y (nx5219), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_2)) ;
    inv01 ix5220 (.Y (nx5221), .A (CacheWindow_3__3__0)) ;
    mux21 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix133 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_2), .A0 (
          nx5223), .A1 (nx5225), .S0 (nx8093)) ;
    inv01 ix5222 (.Y (nx5223), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_3)) ;
    inv01 ix5224 (.Y (nx5225), .A (CacheWindow_3__3__1)) ;
    mux21 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix141 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_3), .A0 (
          nx5227), .A1 (nx5229), .S0 (nx8093)) ;
    inv01 ix5226 (.Y (nx5227), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_4)) ;
    inv01 ix5228 (.Y (nx5229), .A (CacheWindow_3__3__2)) ;
    mux21 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix149 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_4), .A0 (
          nx5231), .A1 (nx5233), .S0 (nx8093)) ;
    inv01 ix5230 (.Y (nx5231), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_5)) ;
    inv01 ix5232 (.Y (nx5233), .A (CacheWindow_3__3__3)) ;
    mux21 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix157 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_5), .A0 (
          nx5235), .A1 (nx5237), .S0 (nx8093)) ;
    inv01 ix5234 (.Y (nx5235), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_6)) ;
    inv01 ix5236 (.Y (nx5237), .A (CacheWindow_3__3__4)) ;
    mux21 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix165 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_6), .A0 (
          nx5239), .A1 (nx5241), .S0 (nx8093)) ;
    inv01 ix5238 (.Y (nx5239), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_7)) ;
    inv01 ix5240 (.Y (nx5241), .A (CacheWindow_3__3__5)) ;
    mux21 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix173 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_7), .A0 (
          nx5243), .A1 (nx5245), .S0 (nx8095)) ;
    inv01 ix5242 (.Y (nx5243), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_8)) ;
    inv01 ix5244 (.Y (nx5245), .A (CacheWindow_3__3__6)) ;
    mux21 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix181 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_8), .A0 (
          nx5247), .A1 (nx5249), .S0 (nx8095)) ;
    inv01 ix5246 (.Y (nx5247), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_9)) ;
    inv01 ix5248 (.Y (nx5249), .A (CacheWindow_3__3__7)) ;
    nor02_2x CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix89 (.Y (
             CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_9), .A0 (
             nx8095), .A1 (nx5251)) ;
    inv01 ix5250 (.Y (nx5251), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_10)) ;
    nor02_2x CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix93 (.Y (
             CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_10), .A0 (
             nx8095), .A1 (nx5253)) ;
    inv01 ix5252 (.Y (nx5253), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_11)) ;
    nor02_2x CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix97 (.Y (
             CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_11), .A0 (
             nx8095), .A1 (nx5255)) ;
    inv01 ix5254 (.Y (nx5255), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_12)) ;
    nor02_2x CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix101 (.Y (
             CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_12), .A0 (
             nx8095), .A1 (nx5257)) ;
    inv01 ix5256 (.Y (nx5257), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_13)) ;
    nor02_2x CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix105 (.Y (
             CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_13), .A0 (
             nx8095), .A1 (nx5259)) ;
    inv01 ix5258 (.Y (nx5259), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_14)) ;
    nor02_2x CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix109 (.Y (
             CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_14), .A0 (
             nx8097), .A1 (nx5261)) ;
    inv01 ix5260 (.Y (nx5261), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_15)) ;
    nor02_2x CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix113 (.Y (
             CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_15), .A0 (
             nx8097), .A1 (nx5263)) ;
    inv01 ix5262 (.Y (nx5263), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_16)) ;
    nor02_2x CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix117 (.Y (
             CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_16), .A0 (
             nx8097), .A1 (nx5263)) ;
    mux21 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix189 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothOperand_0), .A0 (nx5265), .A1 (
          nx5267), .S0 (nx8085)) ;
    inv01 ix5264 (.Y (nx5265), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_0)) ;
    inv01 ix5266 (.Y (nx5267), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_0)) ;
    mux21 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix197 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothOperand_1), .A0 (nx5269), .A1 (
          nx5271), .S0 (nx8085)) ;
    inv01 ix5268 (.Y (nx5269), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_1)) ;
    inv01 ix5270 (.Y (nx5271), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_1)) ;
    mux21 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix205 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothOperand_2), .A0 (nx5273), .A1 (
          nx5275), .S0 (nx8085)) ;
    inv01 ix5272 (.Y (nx5273), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_2)) ;
    inv01 ix5274 (.Y (nx5275), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_2)) ;
    mux21 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix213 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothOperand_3), .A0 (nx5277), .A1 (
          nx5279), .S0 (nx8085)) ;
    inv01 ix5276 (.Y (nx5277), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_3)) ;
    inv01 ix5278 (.Y (nx5279), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_3)) ;
    mux21 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix221 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothOperand_4), .A0 (nx5281), .A1 (
          nx5283), .S0 (nx8085)) ;
    inv01 ix5280 (.Y (nx5281), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_4)) ;
    inv01 ix5282 (.Y (nx5283), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_4)) ;
    mux21 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix229 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothOperand_5), .A0 (nx5285), .A1 (
          nx5287), .S0 (nx8087)) ;
    inv01 ix5284 (.Y (nx5285), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_5)) ;
    inv01 ix5286 (.Y (nx5287), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_5)) ;
    mux21 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix237 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothOperand_6), .A0 (nx5289), .A1 (
          nx5291), .S0 (nx8087)) ;
    inv01 ix5288 (.Y (nx5289), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_6)) ;
    inv01 ix5290 (.Y (nx5291), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_6)) ;
    mux21 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix245 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothOperand_7), .A0 (nx5293), .A1 (
          nx5295), .S0 (nx8087)) ;
    inv01 ix5292 (.Y (nx5293), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_7)) ;
    inv01 ix5294 (.Y (nx5295), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_7)) ;
    mux21 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix253 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothOperand_8), .A0 (nx5297), .A1 (
          nx5299), .S0 (nx8087)) ;
    inv01 ix5296 (.Y (nx5297), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_8)) ;
    inv01 ix5298 (.Y (nx5299), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_8)) ;
    mux21 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix261 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothOperand_9), .A0 (nx5301), .A1 (
          nx5303), .S0 (nx8087)) ;
    inv01 ix5300 (.Y (nx5301), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_9)) ;
    inv01 ix5302 (.Y (nx5303), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_9)) ;
    mux21 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix269 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothOperand_10), .A0 (nx5305), .A1 (
          nx5307), .S0 (nx8087)) ;
    inv01 ix5304 (.Y (nx5305), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_10)) ;
    inv01 ix5306 (.Y (nx5307), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_10)) ;
    mux21 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix277 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothOperand_11), .A0 (nx5309), .A1 (
          nx5311), .S0 (nx8087)) ;
    inv01 ix5308 (.Y (nx5309), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_11)) ;
    inv01 ix5310 (.Y (nx5311), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_11)) ;
    mux21 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix285 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothOperand_12), .A0 (nx5313), .A1 (
          nx5315), .S0 (nx8089)) ;
    inv01 ix5312 (.Y (nx5313), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_12)) ;
    inv01 ix5314 (.Y (nx5315), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_12)) ;
    mux21 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix293 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothOperand_13), .A0 (nx5317), .A1 (
          nx5319), .S0 (nx8089)) ;
    inv01 ix5316 (.Y (nx5317), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_13)) ;
    inv01 ix5318 (.Y (nx5319), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_13)) ;
    mux21 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix301 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothOperand_14), .A0 (nx5321), .A1 (
          nx5323), .S0 (nx8089)) ;
    inv01 ix5320 (.Y (nx5321), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_14)) ;
    inv01 ix5322 (.Y (nx5323), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_14)) ;
    mux21 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix309 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothOperand_15), .A0 (nx5325), .A1 (
          nx5327), .S0 (nx8089)) ;
    inv01 ix5324 (.Y (nx5325), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_15)) ;
    inv01 ix5326 (.Y (nx5327), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_15)) ;
    mux21 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix317 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BoothOperand_16), .A0 (nx5329), .A1 (
          nx5331), .S0 (nx8089)) ;
    inv01 ix5328 (.Y (nx5329), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_16)) ;
    inv01 ix5330 (.Y (nx5331), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_16)) ;
    xnor2 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix321 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_AddPToBoothOperand), .A0 (nx8089), .A1 (
          nx5197)) ;
    oai32 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix393 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .A0 (
          nx8587), .A1 (RST), .A2 (nx8099), .B0 (nx5267), .B1 (nx5335)) ;
    oai32 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix403 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .A0 (
          nx8587), .A1 (RST), .A2 (nx8099), .B0 (nx5271), .B1 (nx5335)) ;
    oai32 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix413 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .A0 (
          nx8587), .A1 (RST), .A2 (nx8099), .B0 (nx5275), .B1 (nx5335)) ;
    oai32 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix423 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .A0 (
          nx8587), .A1 (RST), .A2 (nx8099), .B0 (nx5279), .B1 (nx5335)) ;
    oai32 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix433 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .A0 (
          nx8587), .A1 (RST), .A2 (nx8099), .B0 (nx5283), .B1 (nx5335)) ;
    oai32 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix443 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .A0 (
          nx8587), .A1 (RST), .A2 (nx8099), .B0 (nx5287), .B1 (nx5335)) ;
    oai32 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix453 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .A0 (
          nx8587), .A1 (RST), .A2 (nx8101), .B0 (nx5291), .B1 (nx5335)) ;
    oai32 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix463 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .A0 (
          nx8589), .A1 (RST), .A2 (nx8101), .B0 (nx5295), .B1 (nx5337)) ;
    oai32 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix473 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .A0 (
          nx8589), .A1 (RST), .A2 (nx8101), .B0 (nx5299), .B1 (nx5337)) ;
    oai32 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix483 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .A0 (
          nx5339), .A1 (RST), .A2 (nx8101), .B0 (nx5303), .B1 (nx5337)) ;
    inv01 ix5338 (.Y (nx5339), .A (CacheFilter_3__3__0)) ;
    oai32 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix493 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .A0 (
          nx5341), .A1 (RST), .A2 (nx8101), .B0 (nx5307), .B1 (nx5337)) ;
    inv01 ix5340 (.Y (nx5341), .A (CacheFilter_3__3__1)) ;
    oai32 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix503 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .A0 (
          nx5343), .A1 (RST), .A2 (nx8101), .B0 (nx5311), .B1 (nx5337)) ;
    inv01 ix5342 (.Y (nx5343), .A (CacheFilter_3__3__2)) ;
    oai32 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix513 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .A0 (
          nx5345), .A1 (RST), .A2 (nx8101), .B0 (nx5315), .B1 (nx5337)) ;
    inv01 ix5344 (.Y (nx5345), .A (CacheFilter_3__3__3)) ;
    oai32 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix523 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .A0 (
          nx5347), .A1 (RST), .A2 (nx8103), .B0 (nx5319), .B1 (nx5337)) ;
    inv01 ix5346 (.Y (nx5347), .A (CacheFilter_3__3__4)) ;
    oai32 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix533 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .A0 (
          nx5349), .A1 (RST), .A2 (nx8103), .B0 (nx5323), .B1 (nx5351)) ;
    inv01 ix5348 (.Y (nx5349), .A (CacheFilter_3__3__5)) ;
    inv01 ix5350 (.Y (nx5351), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566)) ;
    oai32 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix543 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .A0 (
          nx5353), .A1 (RST), .A2 (nx8103), .B0 (nx5327), .B1 (nx5351)) ;
    inv01 ix5352 (.Y (nx5353), .A (CacheFilter_3__3__6)) ;
    oai32 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix553 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .A0 (
          nx5355), .A1 (RST), .A2 (nx8103), .B0 (nx5331), .B1 (nx5351)) ;
    inv01 ix5354 (.Y (nx5355), .A (CacheFilter_3__3__7)) ;
    nand02_2x CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix633 (.Y (
              nx5335), .A0 (nx7367), .A1 (nx8103)) ;
    nand02_2x CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix635 (.Y (
              nx5337), .A0 (nx7367), .A1 (nx8103)) ;
    oai32 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix393 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .A0 (
          nx8589), .A1 (RST), .A2 (nx8105), .B0 (nx5265), .B1 (nx5357)) ;
    oai32 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix403 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .A0 (
          nx8589), .A1 (RST), .A2 (nx8105), .B0 (nx5269), .B1 (nx5357)) ;
    oai32 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix413 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .A0 (
          nx8589), .A1 (RST), .A2 (nx8105), .B0 (nx5273), .B1 (nx5357)) ;
    oai32 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix423 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .A0 (
          nx8589), .A1 (RST), .A2 (nx8105), .B0 (nx5277), .B1 (nx5357)) ;
    oai32 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix433 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .A0 (
          nx8589), .A1 (RST), .A2 (nx8105), .B0 (nx5281), .B1 (nx5357)) ;
    oai32 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix443 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .A0 (
          nx8591), .A1 (RST), .A2 (nx8105), .B0 (nx5285), .B1 (nx5357)) ;
    oai32 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix453 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .A0 (
          nx8591), .A1 (RST), .A2 (nx8107), .B0 (nx5289), .B1 (nx5357)) ;
    oai32 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix463 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .A0 (
          nx8591), .A1 (RST), .A2 (nx8107), .B0 (nx5293), .B1 (nx5359)) ;
    oai32 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix473 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .A0 (
          nx8591), .A1 (RST), .A2 (nx8107), .B0 (nx5297), .B1 (nx5359)) ;
    oai32 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix483 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .A0 (
          nx5339), .A1 (RST), .A2 (nx8107), .B0 (nx5301), .B1 (nx5359)) ;
    oai32 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix493 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .A0 (
          nx5361), .A1 (RST), .A2 (nx8107), .B0 (nx5305), .B1 (nx5359)) ;
    inv01 ix5360 (.Y (nx5361), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_10)) ;
    oai32 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix503 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .A0 (
          nx5363), .A1 (RST), .A2 (nx8107), .B0 (nx5309), .B1 (nx5359)) ;
    inv01 ix5362 (.Y (nx5363), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_11)) ;
    oai32 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix513 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .A0 (
          nx5365), .A1 (RST), .A2 (nx8107), .B0 (nx5313), .B1 (nx5359)) ;
    inv01 ix5364 (.Y (nx5365), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_12)) ;
    oai32 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix523 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .A0 (
          nx5367), .A1 (RST), .A2 (nx8109), .B0 (nx5317), .B1 (nx5359)) ;
    inv01 ix5366 (.Y (nx5367), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_13)) ;
    oai32 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix533 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .A0 (
          nx5369), .A1 (RST), .A2 (nx8109), .B0 (nx5321), .B1 (nx5371)) ;
    inv01 ix5368 (.Y (nx5369), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_14)) ;
    inv01 ix5370 (.Y (nx5371), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566)) ;
    oai32 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix543 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .A0 (
          nx5373), .A1 (RST), .A2 (nx8109), .B0 (nx5325), .B1 (nx5371)) ;
    inv01 ix5372 (.Y (nx5373), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_15)) ;
    oai32 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix553 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .A0 (
          nx5375), .A1 (RST), .A2 (nx8109), .B0 (nx5329), .B1 (nx5371)) ;
    inv01 ix5374 (.Y (nx5375), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_16)) ;
    nand02_2x CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix633 (.Y (
              nx5357), .A0 (nx7367), .A1 (nx8109)) ;
    nand02_2x CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix635 (.Y (
              nx5359), .A0 (nx7369), .A1 (nx8109)) ;
    oai32 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix393 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .A0 (
          nx5377), .A1 (RST), .A2 (nx8111), .B0 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx384), .B1 (nx5379)) ;
    inv01 ix5376 (.Y (nx5377), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_0)) ;
    oai32 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix403 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .A0 (
          nx5381), .A1 (RST), .A2 (nx8111), .B0 (nx5197), .B1 (nx5379)) ;
    inv01 ix5380 (.Y (nx5381), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_1)) ;
    oai32 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix413 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .A0 (
          nx5383), .A1 (RST), .A2 (nx8111), .B0 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx387), .B1 (nx5379)) ;
    inv01 ix5382 (.Y (nx5383), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_2)) ;
    oai32 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix423 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .A0 (
          nx5385), .A1 (RST), .A2 (nx8111), .B0 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx399), .B1 (nx5379)) ;
    inv01 ix5384 (.Y (nx5385), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_3)) ;
    oai32 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix433 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .A0 (
          nx5387), .A1 (RST), .A2 (nx8111), .B0 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx409), .B1 (nx5379)) ;
    inv01 ix5386 (.Y (nx5387), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_4)) ;
    oai32 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix443 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .A0 (
          nx5389), .A1 (RST), .A2 (nx8111), .B0 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx419), .B1 (nx5379)) ;
    inv01 ix5388 (.Y (nx5389), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_5)) ;
    oai32 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix453 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .A0 (
          nx5391), .A1 (RST), .A2 (nx8111), .B0 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx429), .B1 (nx5379)) ;
    inv01 ix5390 (.Y (nx5391), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_6)) ;
    oai32 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix463 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .A0 (
          nx5393), .A1 (RST), .A2 (nx8113), .B0 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx439), .B1 (nx5395)) ;
    inv01 ix5392 (.Y (nx5393), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_7)) ;
    oai32 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix473 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .A0 (
          nx5397), .A1 (RST), .A2 (nx8113), .B0 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx449), .B1 (nx5395)) ;
    inv01 ix5396 (.Y (nx5397), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_8)) ;
    oai32 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix483 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .A0 (
          nx5399), .A1 (RST), .A2 (nx8113), .B0 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx469), .B1 (nx5395)) ;
    inv01 ix5398 (.Y (nx5399), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_9)) ;
    oai32 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix493 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .A0 (
          nx5401), .A1 (RST), .A2 (nx8113), .B0 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx477), .B1 (nx5395)) ;
    inv01 ix5400 (.Y (nx5401), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_10)) ;
    oai32 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix503 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .A0 (
          nx5403), .A1 (RST), .A2 (nx8113), .B0 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx485), .B1 (nx5395)) ;
    inv01 ix5402 (.Y (nx5403), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_11)) ;
    oai32 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix513 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .A0 (
          nx5405), .A1 (RST), .A2 (nx8113), .B0 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx493), .B1 (nx5395)) ;
    inv01 ix5404 (.Y (nx5405), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_12)) ;
    oai32 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix523 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .A0 (
          nx5407), .A1 (RST), .A2 (nx8113), .B0 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx501), .B1 (nx5395)) ;
    inv01 ix5406 (.Y (nx5407), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_13)) ;
    oai32 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix533 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .A0 (
          nx5409), .A1 (RST), .A2 (nx8115), .B0 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx509), .B1 (nx5411)) ;
    inv01 ix5408 (.Y (nx5409), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_14)) ;
    inv01 ix5410 (.Y (nx5411), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566)) ;
    oai32 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix543 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .A0 (
          nx5413), .A1 (RST), .A2 (nx8115), .B0 (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_nx517), .B1 (nx5411)) ;
    inv01 ix5412 (.Y (nx5413), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_15)) ;
    oai32 CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix553 (.Y (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .A0 (
          nx5415), .A1 (RST), .A2 (nx8115), .B0 (nx5213), .B1 (nx5411)) ;
    inv01 ix5414 (.Y (nx5415), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_16)) ;
    nand02_2x CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix633 (.Y (
              nx5379), .A0 (nx7369), .A1 (nx8115)) ;
    nand02_2x CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix635 (.Y (
              nx5395), .A0 (nx7369), .A1 (nx8115)) ;
    mux21 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix404 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx403), .A0 (nx5417), .A1 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_2), .S0 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx395)) ;
    inv01 ix5416 (.Y (nx5417), .A (CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx391)) ;
    mux21 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix414 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx413), .A0 (nx5419), .A1 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_3), .S0 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx405)) ;
    inv01 ix5418 (.Y (nx5419), .A (CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx403)) ;
    mux21 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix424 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx423), .A0 (nx5421), .A1 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_4), .S0 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx415)) ;
    inv01 ix5420 (.Y (nx5421), .A (CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx413)) ;
    mux21 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix434 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx433), .A0 (nx5423), .A1 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_5), .S0 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx425)) ;
    inv01 ix5422 (.Y (nx5423), .A (CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx423)) ;
    mux21 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix444 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx443), .A0 (nx5425), .A1 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_6), .S0 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx435)) ;
    inv01 ix5424 (.Y (nx5425), .A (CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx433)) ;
    mux21 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix454 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx453), .A0 (nx5427), .A1 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_7), .S0 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx445)) ;
    inv01 ix5426 (.Y (nx5427), .A (CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx443)) ;
    mux21 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix462 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx461), .A0 (nx5429), .A1 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_8), .S0 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx455)) ;
    inv01 ix5428 (.Y (nx5429), .A (CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx453)) ;
    mux21 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix468 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx467), .A0 (nx5431), .A1 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_9), .S0 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx463)) ;
    inv01 ix5430 (.Y (nx5431), .A (CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx461)) ;
    mux21 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix476 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx475), .A0 (nx5433), .A1 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_10), .S0 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx471)) ;
    inv01 ix5432 (.Y (nx5433), .A (CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx467)) ;
    mux21 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix484 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx483), .A0 (nx5435), .A1 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_11), .S0 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx479)) ;
    inv01 ix5434 (.Y (nx5435), .A (CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx475)) ;
    mux21 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix492 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx491), .A0 (nx5437), .A1 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_12), .S0 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx487)) ;
    inv01 ix5436 (.Y (nx5437), .A (CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx483)) ;
    mux21 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix500 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx499), .A0 (nx5439), .A1 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_13), .S0 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx495)) ;
    inv01 ix5438 (.Y (nx5439), .A (CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx491)) ;
    mux21 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix508 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx507), .A0 (nx5441), .A1 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_14), .S0 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx503)) ;
    inv01 ix5440 (.Y (nx5441), .A (CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx499)) ;
    mux21 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix516 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx515), .A0 (nx5443), .A1 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_15), .S0 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx511)) ;
    inv01 ix5442 (.Y (nx5443), .A (CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx507)) ;
    mux21 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix161 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_1), .A0 (nx5445), .A1 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx379), .S0 (nx8119)) ;
    inv01 ix5444 (.Y (nx5445), .A (CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_1)) ;
    mux21 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix181 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_2), .A0 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx387), .A1 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx389), .S0 (nx8119)) ;
    mux21 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix201 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_3), .A0 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx399), .A1 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx401), .S0 (nx8119)) ;
    mux21 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix221 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_4), .A0 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx409), .A1 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx411), .S0 (nx8119)) ;
    mux21 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix241 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_5), .A0 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx419), .A1 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx421), .S0 (nx8119)) ;
    mux21 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix261 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_6), .A0 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx429), .A1 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx431), .S0 (nx8119)) ;
    mux21 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix281 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_7), .A0 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx439), .A1 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx441), .S0 (nx8119)) ;
    mux21 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix301 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_8), .A0 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx449), .A1 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx451), .S0 (nx8121)) ;
    mux21 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix321 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_9), .A0 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx469), .A1 (nx5447), .S0 (nx8121)) ;
    inv01 ix5446 (.Y (nx5447), .A (CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx316)) ;
    mux21 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix341 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_10), .A0 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx477), .A1 (nx5449), .S0 (nx8121)) ;
    inv01 ix5448 (.Y (nx5449), .A (CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx336)) ;
    mux21 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix361 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_11), .A0 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx485), .A1 (nx5451), .S0 (nx8121)) ;
    inv01 ix5450 (.Y (nx5451), .A (CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx356)) ;
    mux21 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix381 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_12), .A0 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx493), .A1 (nx5453), .S0 (nx8121)) ;
    inv01 ix5452 (.Y (nx5453), .A (CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx376)) ;
    mux21 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix401 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_13), .A0 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx501), .A1 (nx5455), .S0 (nx8121)) ;
    inv01 ix5454 (.Y (nx5455), .A (CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx396)) ;
    mux21 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix421 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_14), .A0 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx509), .A1 (nx5457), .S0 (nx8121)) ;
    inv01 ix5456 (.Y (nx5457), .A (CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx416)) ;
    mux21 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix441 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_15), .A0 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx517), .A1 (nx5459), .S0 (nx8123)) ;
    inv01 ix5458 (.Y (nx5459), .A (CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx436)) ;
    mux21 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_ix461 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_16), .A0 (nx5461), 
          .A1 (nx5463), .S0 (nx8123)) ;
    inv01 ix5460 (.Y (nx5461), .A (CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothP_16)
          ) ;
    inv01 ix5462 (.Y (nx5463), .A (CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx456)) ;
    nor02_2x CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix81 (.Y (
             CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_nx80), .A0 (Instr), .A1 (
             nx7313)) ;
    nor02_2x CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix319 (.Y (
             CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642), .A0 (
             CALCULATOR_Start_dup_1287), .A1 (
             CALCULATOR_CalculatingBooth_dup_1224)) ;
    nor02_2x CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix85 (.Y (
             CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_0), .A0 (
             nx8133), .A1 (nx5465)) ;
    inv01 ix5464 (.Y (nx5465), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_1)) ;
    mux21 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix125 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_1), .A0 (
          nx5467), .A1 (nx5469), .S0 (nx8133)) ;
    inv01 ix5466 (.Y (nx5467), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_2)) ;
    inv01 ix5468 (.Y (nx5469), .A (CacheWindow_3__4__0)) ;
    mux21 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix133 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_2), .A0 (
          nx5471), .A1 (nx5473), .S0 (nx8133)) ;
    inv01 ix5470 (.Y (nx5471), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_3)) ;
    inv01 ix5472 (.Y (nx5473), .A (CacheWindow_3__4__1)) ;
    mux21 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix141 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_3), .A0 (
          nx5475), .A1 (nx5477), .S0 (nx8133)) ;
    inv01 ix5474 (.Y (nx5475), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_4)) ;
    inv01 ix5476 (.Y (nx5477), .A (CacheWindow_3__4__2)) ;
    mux21 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix149 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_4), .A0 (
          nx5479), .A1 (nx5481), .S0 (nx8133)) ;
    inv01 ix5478 (.Y (nx5479), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_5)) ;
    inv01 ix5480 (.Y (nx5481), .A (CacheWindow_3__4__3)) ;
    mux21 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix157 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_5), .A0 (
          nx5483), .A1 (nx5485), .S0 (nx8133)) ;
    inv01 ix5482 (.Y (nx5483), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_6)) ;
    inv01 ix5484 (.Y (nx5485), .A (CacheWindow_3__4__4)) ;
    mux21 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix165 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_6), .A0 (
          nx5487), .A1 (nx5489), .S0 (nx8133)) ;
    inv01 ix5486 (.Y (nx5487), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_7)) ;
    inv01 ix5488 (.Y (nx5489), .A (CacheWindow_3__4__5)) ;
    mux21 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix173 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_7), .A0 (
          nx5491), .A1 (nx5493), .S0 (nx8135)) ;
    inv01 ix5490 (.Y (nx5491), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_8)) ;
    inv01 ix5492 (.Y (nx5493), .A (CacheWindow_3__4__6)) ;
    mux21 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix181 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_8), .A0 (
          nx5495), .A1 (nx5497), .S0 (nx8135)) ;
    inv01 ix5494 (.Y (nx5495), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_9)) ;
    inv01 ix5496 (.Y (nx5497), .A (CacheWindow_3__4__7)) ;
    nor02_2x CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix89 (.Y (
             CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_9), .A0 (
             nx8135), .A1 (nx5499)) ;
    inv01 ix5498 (.Y (nx5499), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_10)) ;
    nor02_2x CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix93 (.Y (
             CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_10), .A0 (
             nx8135), .A1 (nx5501)) ;
    inv01 ix5500 (.Y (nx5501), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_11)) ;
    nor02_2x CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix97 (.Y (
             CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_11), .A0 (
             nx8135), .A1 (nx5503)) ;
    inv01 ix5502 (.Y (nx5503), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_12)) ;
    nor02_2x CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix101 (.Y (
             CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_12), .A0 (
             nx8135), .A1 (nx5505)) ;
    inv01 ix5504 (.Y (nx5505), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_13)) ;
    nor02_2x CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix105 (.Y (
             CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_13), .A0 (
             nx8135), .A1 (nx5507)) ;
    inv01 ix5506 (.Y (nx5507), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_14)) ;
    nor02_2x CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix109 (.Y (
             CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_14), .A0 (
             nx8137), .A1 (nx5509)) ;
    inv01 ix5508 (.Y (nx5509), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_15)) ;
    nor02_2x CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix113 (.Y (
             CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_15), .A0 (
             nx8137), .A1 (nx5511)) ;
    inv01 ix5510 (.Y (nx5511), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_16)) ;
    nor02_2x CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix117 (.Y (
             CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_16), .A0 (
             nx8137), .A1 (nx5511)) ;
    mux21 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix189 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothOperand_0), .A0 (nx5513), .A1 (
          nx5515), .S0 (nx8125)) ;
    inv01 ix5512 (.Y (nx5513), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_0)) ;
    inv01 ix5514 (.Y (nx5515), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_0)) ;
    mux21 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix197 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothOperand_1), .A0 (nx5517), .A1 (
          nx5519), .S0 (nx8125)) ;
    inv01 ix5516 (.Y (nx5517), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_1)) ;
    inv01 ix5518 (.Y (nx5519), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_1)) ;
    mux21 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix205 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothOperand_2), .A0 (nx5521), .A1 (
          nx5523), .S0 (nx8125)) ;
    inv01 ix5520 (.Y (nx5521), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_2)) ;
    inv01 ix5522 (.Y (nx5523), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_2)) ;
    mux21 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix213 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothOperand_3), .A0 (nx5525), .A1 (
          nx5527), .S0 (nx8125)) ;
    inv01 ix5524 (.Y (nx5525), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_3)) ;
    inv01 ix5526 (.Y (nx5527), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_3)) ;
    mux21 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix221 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothOperand_4), .A0 (nx5529), .A1 (
          nx5531), .S0 (nx8125)) ;
    inv01 ix5528 (.Y (nx5529), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_4)) ;
    inv01 ix5530 (.Y (nx5531), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_4)) ;
    mux21 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix229 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothOperand_5), .A0 (nx5533), .A1 (
          nx5535), .S0 (nx8127)) ;
    inv01 ix5532 (.Y (nx5533), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_5)) ;
    inv01 ix5534 (.Y (nx5535), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_5)) ;
    mux21 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix237 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothOperand_6), .A0 (nx5537), .A1 (
          nx5539), .S0 (nx8127)) ;
    inv01 ix5536 (.Y (nx5537), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_6)) ;
    inv01 ix5538 (.Y (nx5539), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_6)) ;
    mux21 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix245 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothOperand_7), .A0 (nx5541), .A1 (
          nx5543), .S0 (nx8127)) ;
    inv01 ix5540 (.Y (nx5541), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_7)) ;
    inv01 ix5542 (.Y (nx5543), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_7)) ;
    mux21 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix253 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothOperand_8), .A0 (nx5545), .A1 (
          nx5547), .S0 (nx8127)) ;
    inv01 ix5544 (.Y (nx5545), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_8)) ;
    inv01 ix5546 (.Y (nx5547), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_8)) ;
    mux21 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix261 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothOperand_9), .A0 (nx5549), .A1 (
          nx5551), .S0 (nx8127)) ;
    inv01 ix5548 (.Y (nx5549), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_9)) ;
    inv01 ix5550 (.Y (nx5551), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_9)) ;
    mux21 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix269 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothOperand_10), .A0 (nx5553), .A1 (
          nx5555), .S0 (nx8127)) ;
    inv01 ix5552 (.Y (nx5553), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_10)) ;
    inv01 ix5554 (.Y (nx5555), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_10)) ;
    mux21 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix277 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothOperand_11), .A0 (nx5557), .A1 (
          nx5559), .S0 (nx8127)) ;
    inv01 ix5556 (.Y (nx5557), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_11)) ;
    inv01 ix5558 (.Y (nx5559), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_11)) ;
    mux21 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix285 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothOperand_12), .A0 (nx5561), .A1 (
          nx5563), .S0 (nx8129)) ;
    inv01 ix5560 (.Y (nx5561), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_12)) ;
    inv01 ix5562 (.Y (nx5563), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_12)) ;
    mux21 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix293 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothOperand_13), .A0 (nx5565), .A1 (
          nx5567), .S0 (nx8129)) ;
    inv01 ix5564 (.Y (nx5565), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_13)) ;
    inv01 ix5566 (.Y (nx5567), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_13)) ;
    mux21 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix301 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothOperand_14), .A0 (nx5569), .A1 (
          nx5571), .S0 (nx8129)) ;
    inv01 ix5568 (.Y (nx5569), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_14)) ;
    inv01 ix5570 (.Y (nx5571), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_14)) ;
    mux21 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix309 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothOperand_15), .A0 (nx5573), .A1 (
          nx5575), .S0 (nx8129)) ;
    inv01 ix5572 (.Y (nx5573), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_15)) ;
    inv01 ix5574 (.Y (nx5575), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_15)) ;
    mux21 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix317 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BoothOperand_16), .A0 (nx5577), .A1 (
          nx5579), .S0 (nx8129)) ;
    inv01 ix5576 (.Y (nx5577), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_16)) ;
    inv01 ix5578 (.Y (nx5579), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_16)) ;
    xnor2 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix321 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_AddPToBoothOperand), .A0 (nx8129), .A1 (
          nx5445)) ;
    oai32 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix393 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .A0 (
          nx8593), .A1 (RST), .A2 (nx8139), .B0 (nx5515), .B1 (nx5583)) ;
    oai32 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix403 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .A0 (
          nx8593), .A1 (RST), .A2 (nx8139), .B0 (nx5519), .B1 (nx5583)) ;
    oai32 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix413 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .A0 (
          nx8593), .A1 (RST), .A2 (nx8139), .B0 (nx5523), .B1 (nx5583)) ;
    oai32 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix423 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .A0 (
          nx8593), .A1 (RST), .A2 (nx8139), .B0 (nx5527), .B1 (nx5583)) ;
    oai32 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix433 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .A0 (
          nx8593), .A1 (RST), .A2 (nx8139), .B0 (nx5531), .B1 (nx5583)) ;
    oai32 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix443 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .A0 (
          nx8593), .A1 (RST), .A2 (nx8139), .B0 (nx5535), .B1 (nx5583)) ;
    oai32 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix453 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .A0 (
          nx8593), .A1 (RST), .A2 (nx8141), .B0 (nx5539), .B1 (nx5583)) ;
    oai32 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix463 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .A0 (
          nx8595), .A1 (RST), .A2 (nx8141), .B0 (nx5543), .B1 (nx5585)) ;
    oai32 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix473 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .A0 (
          nx8595), .A1 (RST), .A2 (nx8141), .B0 (nx5547), .B1 (nx5585)) ;
    oai32 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix483 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .A0 (
          nx5587), .A1 (RST), .A2 (nx8141), .B0 (nx5551), .B1 (nx5585)) ;
    inv01 ix5586 (.Y (nx5587), .A (CacheFilter_3__4__0)) ;
    oai32 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix493 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .A0 (
          nx5589), .A1 (RST), .A2 (nx8141), .B0 (nx5555), .B1 (nx5585)) ;
    inv01 ix5588 (.Y (nx5589), .A (CacheFilter_3__4__1)) ;
    oai32 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix503 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .A0 (
          nx5591), .A1 (RST), .A2 (nx8141), .B0 (nx5559), .B1 (nx5585)) ;
    inv01 ix5590 (.Y (nx5591), .A (CacheFilter_3__4__2)) ;
    oai32 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix513 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .A0 (
          nx5593), .A1 (RST), .A2 (nx8141), .B0 (nx5563), .B1 (nx5585)) ;
    inv01 ix5592 (.Y (nx5593), .A (CacheFilter_3__4__3)) ;
    oai32 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix523 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .A0 (
          nx5595), .A1 (RST), .A2 (nx8143), .B0 (nx5567), .B1 (nx5585)) ;
    inv01 ix5594 (.Y (nx5595), .A (CacheFilter_3__4__4)) ;
    oai32 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix533 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .A0 (
          nx5597), .A1 (RST), .A2 (nx8143), .B0 (nx5571), .B1 (nx5599)) ;
    inv01 ix5596 (.Y (nx5597), .A (CacheFilter_3__4__5)) ;
    inv01 ix5598 (.Y (nx5599), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566)) ;
    oai32 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix543 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .A0 (
          nx5601), .A1 (RST), .A2 (nx8143), .B0 (nx5575), .B1 (nx5599)) ;
    inv01 ix5600 (.Y (nx5601), .A (CacheFilter_3__4__6)) ;
    oai32 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix553 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .A0 (
          nx5603), .A1 (RST), .A2 (nx8143), .B0 (nx5579), .B1 (nx5599)) ;
    inv01 ix5602 (.Y (nx5603), .A (CacheFilter_3__4__7)) ;
    nand02_2x CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix633 (.Y (
              nx5583), .A0 (nx7369), .A1 (nx8143)) ;
    nand02_2x CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix635 (.Y (
              nx5585), .A0 (nx7369), .A1 (nx8143)) ;
    oai32 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix393 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .A0 (
          nx8595), .A1 (RST), .A2 (nx8145), .B0 (nx5513), .B1 (nx5605)) ;
    oai32 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix403 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .A0 (
          nx8595), .A1 (RST), .A2 (nx8145), .B0 (nx5517), .B1 (nx5605)) ;
    oai32 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix413 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .A0 (
          nx8595), .A1 (RST), .A2 (nx8145), .B0 (nx5521), .B1 (nx5605)) ;
    oai32 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix423 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .A0 (
          nx8595), .A1 (RST), .A2 (nx8145), .B0 (nx5525), .B1 (nx5605)) ;
    oai32 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix433 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .A0 (
          nx8595), .A1 (RST), .A2 (nx8145), .B0 (nx5529), .B1 (nx5605)) ;
    oai32 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix443 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .A0 (
          nx8597), .A1 (RST), .A2 (nx8145), .B0 (nx5533), .B1 (nx5605)) ;
    oai32 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix453 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .A0 (
          nx8597), .A1 (RST), .A2 (nx8147), .B0 (nx5537), .B1 (nx5605)) ;
    oai32 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix463 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .A0 (
          nx8597), .A1 (RST), .A2 (nx8147), .B0 (nx5541), .B1 (nx5607)) ;
    oai32 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix473 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .A0 (
          nx8597), .A1 (RST), .A2 (nx8147), .B0 (nx5545), .B1 (nx5607)) ;
    oai32 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix483 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .A0 (
          nx5587), .A1 (RST), .A2 (nx8147), .B0 (nx5549), .B1 (nx5607)) ;
    oai32 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix493 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .A0 (
          nx5609), .A1 (RST), .A2 (nx8147), .B0 (nx5553), .B1 (nx5607)) ;
    inv01 ix5608 (.Y (nx5609), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_10)) ;
    oai32 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix503 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .A0 (
          nx5611), .A1 (RST), .A2 (nx8147), .B0 (nx5557), .B1 (nx5607)) ;
    inv01 ix5610 (.Y (nx5611), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_11)) ;
    oai32 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix513 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .A0 (
          nx5613), .A1 (RST), .A2 (nx8147), .B0 (nx5561), .B1 (nx5607)) ;
    inv01 ix5612 (.Y (nx5613), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_12)) ;
    oai32 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix523 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .A0 (
          nx5615), .A1 (RST), .A2 (nx8149), .B0 (nx5565), .B1 (nx5607)) ;
    inv01 ix5614 (.Y (nx5615), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_13)) ;
    oai32 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix533 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .A0 (
          nx5617), .A1 (RST), .A2 (nx8149), .B0 (nx5569), .B1 (nx5619)) ;
    inv01 ix5616 (.Y (nx5617), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_14)) ;
    inv01 ix5618 (.Y (nx5619), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566)) ;
    oai32 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix543 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .A0 (
          nx5621), .A1 (RST), .A2 (nx8149), .B0 (nx5573), .B1 (nx5619)) ;
    inv01 ix5620 (.Y (nx5621), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_15)) ;
    oai32 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix553 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .A0 (
          nx5623), .A1 (RST), .A2 (nx8149), .B0 (nx5577), .B1 (nx5619)) ;
    inv01 ix5622 (.Y (nx5623), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_16)) ;
    nand02_2x CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix633 (.Y (
              nx5605), .A0 (nx7369), .A1 (nx8149)) ;
    nand02_2x CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix635 (.Y (
              nx5607), .A0 (nx7369), .A1 (nx8149)) ;
    oai32 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix393 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .A0 (
          nx5625), .A1 (RST), .A2 (nx8151), .B0 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_nx384), .B1 (nx5627)) ;
    inv01 ix5624 (.Y (nx5625), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_0)) ;
    oai32 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix403 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .A0 (
          nx5629), .A1 (RST), .A2 (nx8151), .B0 (nx5445), .B1 (nx5627)) ;
    inv01 ix5628 (.Y (nx5629), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_1)) ;
    oai32 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix413 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .A0 (
          nx5631), .A1 (RST), .A2 (nx8151), .B0 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx387), .B1 (nx5627)) ;
    inv01 ix5630 (.Y (nx5631), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_2)) ;
    oai32 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix423 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .A0 (
          nx5633), .A1 (RST), .A2 (nx8151), .B0 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx399), .B1 (nx5627)) ;
    inv01 ix5632 (.Y (nx5633), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_3)) ;
    oai32 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix433 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .A0 (
          nx5635), .A1 (RST), .A2 (nx8151), .B0 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx409), .B1 (nx5627)) ;
    inv01 ix5634 (.Y (nx5635), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_4)) ;
    oai32 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix443 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .A0 (
          nx5637), .A1 (RST), .A2 (nx8151), .B0 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx419), .B1 (nx5627)) ;
    inv01 ix5636 (.Y (nx5637), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_5)) ;
    oai32 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix453 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .A0 (
          nx5639), .A1 (RST), .A2 (nx8151), .B0 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx429), .B1 (nx5627)) ;
    inv01 ix5638 (.Y (nx5639), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_6)) ;
    oai32 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix463 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .A0 (
          nx5641), .A1 (RST), .A2 (nx8153), .B0 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx439), .B1 (nx5643)) ;
    inv01 ix5640 (.Y (nx5641), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_7)) ;
    oai32 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix473 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .A0 (
          nx5645), .A1 (RST), .A2 (nx8153), .B0 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx449), .B1 (nx5643)) ;
    inv01 ix5644 (.Y (nx5645), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_8)) ;
    oai32 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix483 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .A0 (
          nx5647), .A1 (RST), .A2 (nx8153), .B0 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx469), .B1 (nx5643)) ;
    inv01 ix5646 (.Y (nx5647), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_9)) ;
    oai32 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix493 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .A0 (
          nx5649), .A1 (RST), .A2 (nx8153), .B0 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx477), .B1 (nx5643)) ;
    inv01 ix5648 (.Y (nx5649), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_10)) ;
    oai32 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix503 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .A0 (
          nx5651), .A1 (RST), .A2 (nx8153), .B0 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx485), .B1 (nx5643)) ;
    inv01 ix5650 (.Y (nx5651), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_11)) ;
    oai32 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix513 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .A0 (
          nx5653), .A1 (RST), .A2 (nx8153), .B0 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx493), .B1 (nx5643)) ;
    inv01 ix5652 (.Y (nx5653), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_12)) ;
    oai32 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix523 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .A0 (
          nx5655), .A1 (RST), .A2 (nx8153), .B0 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx501), .B1 (nx5643)) ;
    inv01 ix5654 (.Y (nx5655), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_13)) ;
    oai32 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix533 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .A0 (
          nx5657), .A1 (RST), .A2 (nx8155), .B0 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx509), .B1 (nx5659)) ;
    inv01 ix5656 (.Y (nx5657), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_14)) ;
    inv01 ix5658 (.Y (nx5659), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566)) ;
    oai32 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix543 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .A0 (
          nx5661), .A1 (RST), .A2 (nx8155), .B0 (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_nx517), .B1 (nx5659)) ;
    inv01 ix5660 (.Y (nx5661), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_15)) ;
    oai32 CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix553 (.Y (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .A0 (
          nx5663), .A1 (RST), .A2 (nx8155), .B0 (nx5461), .B1 (nx5659)) ;
    inv01 ix5662 (.Y (nx5663), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_16)) ;
    nand02_2x CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix633 (.Y (
              nx5627), .A0 (nx7371), .A1 (nx8155)) ;
    nand02_2x CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix635 (.Y (
              nx5643), .A0 (nx7371), .A1 (nx8155)) ;
    mux21 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix404 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx403), .A0 (nx5665), .A1 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_2), .S0 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx395)) ;
    inv01 ix5664 (.Y (nx5665), .A (CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx391)) ;
    mux21 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix414 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx413), .A0 (nx5667), .A1 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_3), .S0 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx405)) ;
    inv01 ix5666 (.Y (nx5667), .A (CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx403)) ;
    mux21 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix424 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx423), .A0 (nx5669), .A1 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_4), .S0 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx415)) ;
    inv01 ix5668 (.Y (nx5669), .A (CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx413)) ;
    mux21 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix434 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx433), .A0 (nx5671), .A1 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_5), .S0 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx425)) ;
    inv01 ix5670 (.Y (nx5671), .A (CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx423)) ;
    mux21 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix444 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx443), .A0 (nx5673), .A1 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_6), .S0 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx435)) ;
    inv01 ix5672 (.Y (nx5673), .A (CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx433)) ;
    mux21 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix454 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx453), .A0 (nx5675), .A1 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_7), .S0 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx445)) ;
    inv01 ix5674 (.Y (nx5675), .A (CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx443)) ;
    mux21 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix462 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx461), .A0 (nx5677), .A1 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_8), .S0 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx455)) ;
    inv01 ix5676 (.Y (nx5677), .A (CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx453)) ;
    mux21 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix468 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx467), .A0 (nx5679), .A1 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_9), .S0 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx463)) ;
    inv01 ix5678 (.Y (nx5679), .A (CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx461)) ;
    mux21 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix476 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx475), .A0 (nx5681), .A1 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_10), .S0 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx471)) ;
    inv01 ix5680 (.Y (nx5681), .A (CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx467)) ;
    mux21 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix484 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx483), .A0 (nx5683), .A1 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_11), .S0 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx479)) ;
    inv01 ix5682 (.Y (nx5683), .A (CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx475)) ;
    mux21 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix492 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx491), .A0 (nx5685), .A1 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_12), .S0 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx487)) ;
    inv01 ix5684 (.Y (nx5685), .A (CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx483)) ;
    mux21 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix500 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx499), .A0 (nx5687), .A1 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_13), .S0 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx495)) ;
    inv01 ix5686 (.Y (nx5687), .A (CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx491)) ;
    mux21 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix508 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx507), .A0 (nx5689), .A1 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_14), .S0 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx503)) ;
    inv01 ix5688 (.Y (nx5689), .A (CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx499)) ;
    mux21 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix516 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx515), .A0 (nx5691), .A1 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_15), .S0 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx511)) ;
    inv01 ix5690 (.Y (nx5691), .A (CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx507)) ;
    mux21 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix161 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_1), .A0 (nx5693), .A1 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx379), .S0 (nx8159)) ;
    inv01 ix5692 (.Y (nx5693), .A (CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_1)) ;
    mux21 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix181 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_2), .A0 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx387), .A1 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx389), .S0 (nx8159)) ;
    mux21 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix201 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_3), .A0 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx399), .A1 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx401), .S0 (nx8159)) ;
    mux21 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix221 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_4), .A0 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx409), .A1 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx411), .S0 (nx8159)) ;
    mux21 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix241 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_5), .A0 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx419), .A1 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx421), .S0 (nx8159)) ;
    mux21 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix261 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_6), .A0 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx429), .A1 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx431), .S0 (nx8159)) ;
    mux21 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix281 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_7), .A0 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx439), .A1 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx441), .S0 (nx8159)) ;
    mux21 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix301 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_8), .A0 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx449), .A1 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx451), .S0 (nx8161)) ;
    mux21 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix321 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_9), .A0 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx469), .A1 (nx5695), .S0 (nx8161)) ;
    inv01 ix5694 (.Y (nx5695), .A (CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx316)) ;
    mux21 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix341 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_10), .A0 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx477), .A1 (nx5697), .S0 (nx8161)) ;
    inv01 ix5696 (.Y (nx5697), .A (CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx336)) ;
    mux21 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix361 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_11), .A0 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx485), .A1 (nx5699), .S0 (nx8161)) ;
    inv01 ix5698 (.Y (nx5699), .A (CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx356)) ;
    mux21 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix381 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_12), .A0 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx493), .A1 (nx5701), .S0 (nx8161)) ;
    inv01 ix5700 (.Y (nx5701), .A (CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx376)) ;
    mux21 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix401 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_13), .A0 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx501), .A1 (nx5703), .S0 (nx8161)) ;
    inv01 ix5702 (.Y (nx5703), .A (CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx396)) ;
    mux21 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix421 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_14), .A0 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx509), .A1 (nx5705), .S0 (nx8161)) ;
    inv01 ix5704 (.Y (nx5705), .A (CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx416)) ;
    mux21 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix441 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_15), .A0 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx517), .A1 (nx5707), .S0 (nx8163)) ;
    inv01 ix5706 (.Y (nx5707), .A (CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx436)) ;
    mux21 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_ix461 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_16), .A0 (nx5709), 
          .A1 (nx5711), .S0 (nx8163)) ;
    inv01 ix5708 (.Y (nx5709), .A (CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothP_16)
          ) ;
    inv01 ix5710 (.Y (nx5711), .A (CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx456)) ;
    nor02_2x CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix81 (.Y (
             CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_nx80), .A0 (Instr), .A1 (
             nx7313)) ;
    nor02_2x CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix319 (.Y (
             CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642), .A0 (
             CALCULATOR_Start_dup_1300), .A1 (
             CALCULATOR_CalculatingBooth_dup_1224)) ;
    nor02_2x CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix85 (.Y (
             CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_0), .A0 (
             nx8173), .A1 (nx5713)) ;
    inv01 ix5712 (.Y (nx5713), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_1)) ;
    mux21 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix125 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_1), .A0 (
          nx5715), .A1 (nx5717), .S0 (nx8173)) ;
    inv01 ix5714 (.Y (nx5715), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_2)) ;
    inv01 ix5716 (.Y (nx5717), .A (CacheWindow_4__0__0)) ;
    mux21 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix133 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_2), .A0 (
          nx5719), .A1 (nx5721), .S0 (nx8173)) ;
    inv01 ix5718 (.Y (nx5719), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_3)) ;
    inv01 ix5720 (.Y (nx5721), .A (CacheWindow_4__0__1)) ;
    mux21 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix141 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_3), .A0 (
          nx5723), .A1 (nx5725), .S0 (nx8173)) ;
    inv01 ix5722 (.Y (nx5723), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_4)) ;
    inv01 ix5724 (.Y (nx5725), .A (CacheWindow_4__0__2)) ;
    mux21 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix149 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_4), .A0 (
          nx5727), .A1 (nx5729), .S0 (nx8173)) ;
    inv01 ix5726 (.Y (nx5727), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_5)) ;
    inv01 ix5728 (.Y (nx5729), .A (CacheWindow_4__0__3)) ;
    mux21 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix157 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_5), .A0 (
          nx5731), .A1 (nx5733), .S0 (nx8173)) ;
    inv01 ix5730 (.Y (nx5731), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_6)) ;
    inv01 ix5732 (.Y (nx5733), .A (CacheWindow_4__0__4)) ;
    mux21 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix165 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_6), .A0 (
          nx5735), .A1 (nx5737), .S0 (nx8173)) ;
    inv01 ix5734 (.Y (nx5735), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_7)) ;
    inv01 ix5736 (.Y (nx5737), .A (CacheWindow_4__0__5)) ;
    mux21 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix173 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_7), .A0 (
          nx5739), .A1 (nx5741), .S0 (nx8175)) ;
    inv01 ix5738 (.Y (nx5739), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_8)) ;
    inv01 ix5740 (.Y (nx5741), .A (CacheWindow_4__0__6)) ;
    mux21 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix181 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_8), .A0 (
          nx5743), .A1 (nx5745), .S0 (nx8175)) ;
    inv01 ix5742 (.Y (nx5743), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_9)) ;
    inv01 ix5744 (.Y (nx5745), .A (CacheWindow_4__0__7)) ;
    nor02_2x CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix89 (.Y (
             CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_9), .A0 (
             nx8175), .A1 (nx5747)) ;
    inv01 ix5746 (.Y (nx5747), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_10)) ;
    nor02_2x CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix93 (.Y (
             CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_10), .A0 (
             nx8175), .A1 (nx5749)) ;
    inv01 ix5748 (.Y (nx5749), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_11)) ;
    nor02_2x CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix97 (.Y (
             CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_11), .A0 (
             nx8175), .A1 (nx5751)) ;
    inv01 ix5750 (.Y (nx5751), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_12)) ;
    nor02_2x CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix101 (.Y (
             CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_12), .A0 (
             nx8175), .A1 (nx5753)) ;
    inv01 ix5752 (.Y (nx5753), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_13)) ;
    nor02_2x CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix105 (.Y (
             CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_13), .A0 (
             nx8175), .A1 (nx5755)) ;
    inv01 ix5754 (.Y (nx5755), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_14)) ;
    nor02_2x CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix109 (.Y (
             CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_14), .A0 (
             nx8177), .A1 (nx5757)) ;
    inv01 ix5756 (.Y (nx5757), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_15)) ;
    nor02_2x CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix113 (.Y (
             CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_15), .A0 (
             nx8177), .A1 (nx5759)) ;
    inv01 ix5758 (.Y (nx5759), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_16)) ;
    nor02_2x CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix117 (.Y (
             CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_16), .A0 (
             nx8177), .A1 (nx5759)) ;
    mux21 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix189 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothOperand_0), .A0 (nx5761), .A1 (
          nx5763), .S0 (nx8165)) ;
    inv01 ix5760 (.Y (nx5761), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_0)) ;
    inv01 ix5762 (.Y (nx5763), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_0)) ;
    mux21 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix197 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothOperand_1), .A0 (nx5765), .A1 (
          nx5767), .S0 (nx8165)) ;
    inv01 ix5764 (.Y (nx5765), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_1)) ;
    inv01 ix5766 (.Y (nx5767), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_1)) ;
    mux21 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix205 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothOperand_2), .A0 (nx5769), .A1 (
          nx5771), .S0 (nx8165)) ;
    inv01 ix5768 (.Y (nx5769), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_2)) ;
    inv01 ix5770 (.Y (nx5771), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_2)) ;
    mux21 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix213 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothOperand_3), .A0 (nx5773), .A1 (
          nx5775), .S0 (nx8165)) ;
    inv01 ix5772 (.Y (nx5773), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_3)) ;
    inv01 ix5774 (.Y (nx5775), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_3)) ;
    mux21 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix221 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothOperand_4), .A0 (nx5777), .A1 (
          nx5779), .S0 (nx8165)) ;
    inv01 ix5776 (.Y (nx5777), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_4)) ;
    inv01 ix5778 (.Y (nx5779), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_4)) ;
    mux21 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix229 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothOperand_5), .A0 (nx5781), .A1 (
          nx5783), .S0 (nx8167)) ;
    inv01 ix5780 (.Y (nx5781), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_5)) ;
    inv01 ix5782 (.Y (nx5783), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_5)) ;
    mux21 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix237 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothOperand_6), .A0 (nx5785), .A1 (
          nx5787), .S0 (nx8167)) ;
    inv01 ix5784 (.Y (nx5785), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_6)) ;
    inv01 ix5786 (.Y (nx5787), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_6)) ;
    mux21 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix245 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothOperand_7), .A0 (nx5789), .A1 (
          nx5791), .S0 (nx8167)) ;
    inv01 ix5788 (.Y (nx5789), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_7)) ;
    inv01 ix5790 (.Y (nx5791), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_7)) ;
    mux21 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix253 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothOperand_8), .A0 (nx5793), .A1 (
          nx5795), .S0 (nx8167)) ;
    inv01 ix5792 (.Y (nx5793), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_8)) ;
    inv01 ix5794 (.Y (nx5795), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_8)) ;
    mux21 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix261 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothOperand_9), .A0 (nx5797), .A1 (
          nx5799), .S0 (nx8167)) ;
    inv01 ix5796 (.Y (nx5797), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_9)) ;
    inv01 ix5798 (.Y (nx5799), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_9)) ;
    mux21 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix269 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothOperand_10), .A0 (nx5801), .A1 (
          nx5803), .S0 (nx8167)) ;
    inv01 ix5800 (.Y (nx5801), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_10)) ;
    inv01 ix5802 (.Y (nx5803), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_10)) ;
    mux21 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix277 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothOperand_11), .A0 (nx5805), .A1 (
          nx5807), .S0 (nx8167)) ;
    inv01 ix5804 (.Y (nx5805), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_11)) ;
    inv01 ix5806 (.Y (nx5807), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_11)) ;
    mux21 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix285 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothOperand_12), .A0 (nx5809), .A1 (
          nx5811), .S0 (nx8169)) ;
    inv01 ix5808 (.Y (nx5809), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_12)) ;
    inv01 ix5810 (.Y (nx5811), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_12)) ;
    mux21 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix293 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothOperand_13), .A0 (nx5813), .A1 (
          nx5815), .S0 (nx8169)) ;
    inv01 ix5812 (.Y (nx5813), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_13)) ;
    inv01 ix5814 (.Y (nx5815), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_13)) ;
    mux21 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix301 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothOperand_14), .A0 (nx5817), .A1 (
          nx5819), .S0 (nx8169)) ;
    inv01 ix5816 (.Y (nx5817), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_14)) ;
    inv01 ix5818 (.Y (nx5819), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_14)) ;
    mux21 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix309 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothOperand_15), .A0 (nx5821), .A1 (
          nx5823), .S0 (nx8169)) ;
    inv01 ix5820 (.Y (nx5821), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_15)) ;
    inv01 ix5822 (.Y (nx5823), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_15)) ;
    mux21 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix317 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BoothOperand_16), .A0 (nx5825), .A1 (
          nx5827), .S0 (nx8169)) ;
    inv01 ix5824 (.Y (nx5825), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_16)) ;
    inv01 ix5826 (.Y (nx5827), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_16)) ;
    xnor2 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix321 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_AddPToBoothOperand), .A0 (nx8169), .A1 (
          nx5693)) ;
    oai32 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix393 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .A0 (
          nx8599), .A1 (RST), .A2 (nx8179), .B0 (nx5763), .B1 (nx5831)) ;
    oai32 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix403 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .A0 (
          nx8599), .A1 (RST), .A2 (nx8179), .B0 (nx5767), .B1 (nx5831)) ;
    oai32 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix413 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .A0 (
          nx8599), .A1 (RST), .A2 (nx8179), .B0 (nx5771), .B1 (nx5831)) ;
    oai32 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix423 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .A0 (
          nx8599), .A1 (RST), .A2 (nx8179), .B0 (nx5775), .B1 (nx5831)) ;
    oai32 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix433 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .A0 (
          nx8599), .A1 (RST), .A2 (nx8179), .B0 (nx5779), .B1 (nx5831)) ;
    oai32 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix443 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .A0 (
          nx8599), .A1 (RST), .A2 (nx8179), .B0 (nx5783), .B1 (nx5831)) ;
    oai32 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix453 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .A0 (
          nx8599), .A1 (RST), .A2 (nx8181), .B0 (nx5787), .B1 (nx5831)) ;
    oai32 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix463 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .A0 (
          nx8601), .A1 (RST), .A2 (nx8181), .B0 (nx5791), .B1 (nx5833)) ;
    oai32 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix473 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .A0 (
          nx8601), .A1 (RST), .A2 (nx8181), .B0 (nx5795), .B1 (nx5833)) ;
    oai32 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix483 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .A0 (
          nx5835), .A1 (RST), .A2 (nx8181), .B0 (nx5799), .B1 (nx5833)) ;
    inv01 ix5834 (.Y (nx5835), .A (CacheFilter_4__0__0)) ;
    oai32 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix493 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .A0 (
          nx5837), .A1 (RST), .A2 (nx8181), .B0 (nx5803), .B1 (nx5833)) ;
    inv01 ix5836 (.Y (nx5837), .A (CacheFilter_4__0__1)) ;
    oai32 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix503 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .A0 (
          nx5839), .A1 (RST), .A2 (nx8181), .B0 (nx5807), .B1 (nx5833)) ;
    inv01 ix5838 (.Y (nx5839), .A (CacheFilter_4__0__2)) ;
    oai32 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix513 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .A0 (
          nx5841), .A1 (RST), .A2 (nx8181), .B0 (nx5811), .B1 (nx5833)) ;
    inv01 ix5840 (.Y (nx5841), .A (CacheFilter_4__0__3)) ;
    oai32 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix523 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .A0 (
          nx5843), .A1 (RST), .A2 (nx8183), .B0 (nx5815), .B1 (nx5833)) ;
    inv01 ix5842 (.Y (nx5843), .A (CacheFilter_4__0__4)) ;
    oai32 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix533 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .A0 (
          nx5845), .A1 (RST), .A2 (nx8183), .B0 (nx5819), .B1 (nx5847)) ;
    inv01 ix5844 (.Y (nx5845), .A (CacheFilter_4__0__5)) ;
    inv01 ix5846 (.Y (nx5847), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566)) ;
    oai32 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix543 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .A0 (
          nx5849), .A1 (RST), .A2 (nx8183), .B0 (nx5823), .B1 (nx5847)) ;
    inv01 ix5848 (.Y (nx5849), .A (CacheFilter_4__0__6)) ;
    oai32 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix553 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .A0 (
          nx5851), .A1 (RST), .A2 (nx8183), .B0 (nx5827), .B1 (nx5847)) ;
    inv01 ix5850 (.Y (nx5851), .A (CacheFilter_4__0__7)) ;
    nand02_2x CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix633 (.Y (
              nx5831), .A0 (nx7371), .A1 (nx8183)) ;
    nand02_2x CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix635 (.Y (
              nx5833), .A0 (nx7371), .A1 (nx8183)) ;
    oai32 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix393 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .A0 (
          nx8601), .A1 (RST), .A2 (nx8185), .B0 (nx5761), .B1 (nx5853)) ;
    oai32 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix403 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .A0 (
          nx8601), .A1 (RST), .A2 (nx8185), .B0 (nx5765), .B1 (nx5853)) ;
    oai32 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix413 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .A0 (
          nx8601), .A1 (RST), .A2 (nx8185), .B0 (nx5769), .B1 (nx5853)) ;
    oai32 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix423 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .A0 (
          nx8601), .A1 (RST), .A2 (nx8185), .B0 (nx5773), .B1 (nx5853)) ;
    oai32 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix433 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .A0 (
          nx8601), .A1 (RST), .A2 (nx8185), .B0 (nx5777), .B1 (nx5853)) ;
    oai32 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix443 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .A0 (
          nx8603), .A1 (RST), .A2 (nx8185), .B0 (nx5781), .B1 (nx5853)) ;
    oai32 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix453 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .A0 (
          nx8603), .A1 (RST), .A2 (nx8187), .B0 (nx5785), .B1 (nx5853)) ;
    oai32 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix463 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .A0 (
          nx8603), .A1 (RST), .A2 (nx8187), .B0 (nx5789), .B1 (nx5855)) ;
    oai32 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix473 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .A0 (
          nx8603), .A1 (RST), .A2 (nx8187), .B0 (nx5793), .B1 (nx5855)) ;
    oai32 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix483 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .A0 (
          nx5835), .A1 (RST), .A2 (nx8187), .B0 (nx5797), .B1 (nx5855)) ;
    oai32 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix493 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .A0 (
          nx5857), .A1 (RST), .A2 (nx8187), .B0 (nx5801), .B1 (nx5855)) ;
    inv01 ix5856 (.Y (nx5857), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_10)) ;
    oai32 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix503 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .A0 (
          nx5859), .A1 (RST), .A2 (nx8187), .B0 (nx5805), .B1 (nx5855)) ;
    inv01 ix5858 (.Y (nx5859), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_11)) ;
    oai32 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix513 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .A0 (
          nx5861), .A1 (RST), .A2 (nx8187), .B0 (nx5809), .B1 (nx5855)) ;
    inv01 ix5860 (.Y (nx5861), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_12)) ;
    oai32 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix523 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .A0 (
          nx5863), .A1 (RST), .A2 (nx8189), .B0 (nx5813), .B1 (nx5855)) ;
    inv01 ix5862 (.Y (nx5863), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_13)) ;
    oai32 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix533 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .A0 (
          nx5865), .A1 (RST), .A2 (nx8189), .B0 (nx5817), .B1 (nx5867)) ;
    inv01 ix5864 (.Y (nx5865), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_14)) ;
    inv01 ix5866 (.Y (nx5867), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566)) ;
    oai32 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix543 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .A0 (
          nx5869), .A1 (RST), .A2 (nx8189), .B0 (nx5821), .B1 (nx5867)) ;
    inv01 ix5868 (.Y (nx5869), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_15)) ;
    oai32 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix553 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .A0 (
          nx5871), .A1 (RST), .A2 (nx8189), .B0 (nx5825), .B1 (nx5867)) ;
    inv01 ix5870 (.Y (nx5871), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_16)) ;
    nand02_2x CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix633 (.Y (
              nx5853), .A0 (nx7371), .A1 (nx8189)) ;
    nand02_2x CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix635 (.Y (
              nx5855), .A0 (nx7371), .A1 (nx8189)) ;
    oai32 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix393 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .A0 (
          nx5873), .A1 (RST), .A2 (nx8191), .B0 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_nx384), .B1 (nx5875)) ;
    inv01 ix5872 (.Y (nx5873), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_0)) ;
    oai32 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix403 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .A0 (
          nx5877), .A1 (RST), .A2 (nx8191), .B0 (nx5693), .B1 (nx5875)) ;
    inv01 ix5876 (.Y (nx5877), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_1)) ;
    oai32 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix413 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .A0 (
          nx5879), .A1 (RST), .A2 (nx8191), .B0 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx387), .B1 (nx5875)) ;
    inv01 ix5878 (.Y (nx5879), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_2)) ;
    oai32 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix423 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .A0 (
          nx5881), .A1 (RST), .A2 (nx8191), .B0 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx399), .B1 (nx5875)) ;
    inv01 ix5880 (.Y (nx5881), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_3)) ;
    oai32 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix433 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .A0 (
          nx5883), .A1 (RST), .A2 (nx8191), .B0 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx409), .B1 (nx5875)) ;
    inv01 ix5882 (.Y (nx5883), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_4)) ;
    oai32 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix443 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .A0 (
          nx5885), .A1 (RST), .A2 (nx8191), .B0 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx419), .B1 (nx5875)) ;
    inv01 ix5884 (.Y (nx5885), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_5)) ;
    oai32 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix453 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .A0 (
          nx5887), .A1 (RST), .A2 (nx8191), .B0 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx429), .B1 (nx5875)) ;
    inv01 ix5886 (.Y (nx5887), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_6)) ;
    oai32 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix463 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .A0 (
          nx5889), .A1 (RST), .A2 (nx8193), .B0 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx439), .B1 (nx5891)) ;
    inv01 ix5888 (.Y (nx5889), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_7)) ;
    oai32 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix473 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .A0 (
          nx5893), .A1 (RST), .A2 (nx8193), .B0 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx449), .B1 (nx5891)) ;
    inv01 ix5892 (.Y (nx5893), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_8)) ;
    oai32 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix483 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .A0 (
          nx5895), .A1 (RST), .A2 (nx8193), .B0 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx469), .B1 (nx5891)) ;
    inv01 ix5894 (.Y (nx5895), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_9)) ;
    oai32 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix493 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .A0 (
          nx5897), .A1 (RST), .A2 (nx8193), .B0 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx477), .B1 (nx5891)) ;
    inv01 ix5896 (.Y (nx5897), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_10)) ;
    oai32 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix503 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .A0 (
          nx5899), .A1 (RST), .A2 (nx8193), .B0 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx485), .B1 (nx5891)) ;
    inv01 ix5898 (.Y (nx5899), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_11)) ;
    oai32 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix513 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .A0 (
          nx5901), .A1 (RST), .A2 (nx8193), .B0 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx493), .B1 (nx5891)) ;
    inv01 ix5900 (.Y (nx5901), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_12)) ;
    oai32 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix523 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .A0 (
          nx5903), .A1 (RST), .A2 (nx8193), .B0 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx501), .B1 (nx5891)) ;
    inv01 ix5902 (.Y (nx5903), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_13)) ;
    oai32 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix533 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .A0 (
          nx5905), .A1 (RST), .A2 (nx8195), .B0 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx509), .B1 (nx5907)) ;
    inv01 ix5904 (.Y (nx5905), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_14)) ;
    inv01 ix5906 (.Y (nx5907), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566)) ;
    oai32 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix543 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .A0 (
          nx5909), .A1 (RST), .A2 (nx8195), .B0 (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_nx517), .B1 (nx5907)) ;
    inv01 ix5908 (.Y (nx5909), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_15)) ;
    oai32 CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix553 (.Y (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .A0 (
          nx5911), .A1 (RST), .A2 (nx8195), .B0 (nx5709), .B1 (nx5907)) ;
    inv01 ix5910 (.Y (nx5911), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_16)) ;
    nand02_2x CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix633 (.Y (
              nx5875), .A0 (nx7371), .A1 (nx8195)) ;
    nand02_2x CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix635 (.Y (
              nx5891), .A0 (nx7373), .A1 (nx8195)) ;
    mux21 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix404 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx403), .A0 (nx5913), .A1 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_2), .S0 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx395)) ;
    inv01 ix5912 (.Y (nx5913), .A (CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx391)) ;
    mux21 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix414 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx413), .A0 (nx5915), .A1 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_3), .S0 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx405)) ;
    inv01 ix5914 (.Y (nx5915), .A (CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx403)) ;
    mux21 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix424 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx423), .A0 (nx5917), .A1 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_4), .S0 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx415)) ;
    inv01 ix5916 (.Y (nx5917), .A (CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx413)) ;
    mux21 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix434 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx433), .A0 (nx5919), .A1 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_5), .S0 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx425)) ;
    inv01 ix5918 (.Y (nx5919), .A (CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx423)) ;
    mux21 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix444 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx443), .A0 (nx5921), .A1 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_6), .S0 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx435)) ;
    inv01 ix5920 (.Y (nx5921), .A (CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx433)) ;
    mux21 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix454 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx453), .A0 (nx5923), .A1 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_7), .S0 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx445)) ;
    inv01 ix5922 (.Y (nx5923), .A (CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx443)) ;
    mux21 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix462 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx461), .A0 (nx5925), .A1 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_8), .S0 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx455)) ;
    inv01 ix5924 (.Y (nx5925), .A (CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx453)) ;
    mux21 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix468 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx467), .A0 (nx5927), .A1 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_9), .S0 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx463)) ;
    inv01 ix5926 (.Y (nx5927), .A (CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx461)) ;
    mux21 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix476 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx475), .A0 (nx5929), .A1 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_10), .S0 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx471)) ;
    inv01 ix5928 (.Y (nx5929), .A (CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx467)) ;
    mux21 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix484 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx483), .A0 (nx5931), .A1 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_11), .S0 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx479)) ;
    inv01 ix5930 (.Y (nx5931), .A (CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx475)) ;
    mux21 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix492 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx491), .A0 (nx5933), .A1 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_12), .S0 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx487)) ;
    inv01 ix5932 (.Y (nx5933), .A (CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx483)) ;
    mux21 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix500 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx499), .A0 (nx5935), .A1 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_13), .S0 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx495)) ;
    inv01 ix5934 (.Y (nx5935), .A (CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx491)) ;
    mux21 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix508 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx507), .A0 (nx5937), .A1 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_14), .S0 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx503)) ;
    inv01 ix5936 (.Y (nx5937), .A (CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx499)) ;
    mux21 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix516 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx515), .A0 (nx5939), .A1 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_15), .S0 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx511)) ;
    inv01 ix5938 (.Y (nx5939), .A (CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx507)) ;
    mux21 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix161 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_1), .A0 (nx5941), .A1 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx379), .S0 (nx8199)) ;
    inv01 ix5940 (.Y (nx5941), .A (CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_1)) ;
    mux21 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix181 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_2), .A0 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx387), .A1 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx389), .S0 (nx8199)) ;
    mux21 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix201 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_3), .A0 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx399), .A1 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx401), .S0 (nx8199)) ;
    mux21 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix221 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_4), .A0 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx409), .A1 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx411), .S0 (nx8199)) ;
    mux21 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix241 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_5), .A0 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx419), .A1 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx421), .S0 (nx8199)) ;
    mux21 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix261 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_6), .A0 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx429), .A1 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx431), .S0 (nx8199)) ;
    mux21 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix281 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_7), .A0 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx439), .A1 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx441), .S0 (nx8199)) ;
    mux21 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix301 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_8), .A0 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx449), .A1 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx451), .S0 (nx8201)) ;
    mux21 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix321 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_9), .A0 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx469), .A1 (nx5943), .S0 (nx8201)) ;
    inv01 ix5942 (.Y (nx5943), .A (CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx316)) ;
    mux21 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix341 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_10), .A0 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx477), .A1 (nx5945), .S0 (nx8201)) ;
    inv01 ix5944 (.Y (nx5945), .A (CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx336)) ;
    mux21 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix361 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_11), .A0 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx485), .A1 (nx5947), .S0 (nx8201)) ;
    inv01 ix5946 (.Y (nx5947), .A (CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx356)) ;
    mux21 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix381 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_12), .A0 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx493), .A1 (nx5949), .S0 (nx8201)) ;
    inv01 ix5948 (.Y (nx5949), .A (CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx376)) ;
    mux21 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix401 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_13), .A0 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx501), .A1 (nx5951), .S0 (nx8201)) ;
    inv01 ix5950 (.Y (nx5951), .A (CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx396)) ;
    mux21 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix421 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_14), .A0 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx509), .A1 (nx5953), .S0 (nx8201)) ;
    inv01 ix5952 (.Y (nx5953), .A (CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx416)) ;
    mux21 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix441 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_15), .A0 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx517), .A1 (nx5955), .S0 (nx8203)) ;
    inv01 ix5954 (.Y (nx5955), .A (CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx436)) ;
    mux21 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_ix461 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_16), .A0 (nx5957), 
          .A1 (nx5959), .S0 (nx8203)) ;
    inv01 ix5956 (.Y (nx5957), .A (CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothP_16)
          ) ;
    inv01 ix5958 (.Y (nx5959), .A (CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx456)) ;
    nor02_2x CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix81 (.Y (
             CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_nx80), .A0 (Instr), .A1 (
             nx7299)) ;
    nor02_2x CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix319 (.Y (
             CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642), .A0 (
             CALCULATOR_Start_dup_1313), .A1 (
             CALCULATOR_CalculatingBooth_dup_1315)) ;
    nor02_2x CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix85 (.Y (
             CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_0), .A0 (
             nx8213), .A1 (nx5961)) ;
    inv01 ix5960 (.Y (nx5961), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_1)) ;
    mux21 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix125 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_1), .A0 (
          nx5963), .A1 (nx5965), .S0 (nx8213)) ;
    inv01 ix5962 (.Y (nx5963), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_2)) ;
    inv01 ix5964 (.Y (nx5965), .A (CacheWindow_4__1__0)) ;
    mux21 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix133 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_2), .A0 (
          nx5967), .A1 (nx5969), .S0 (nx8213)) ;
    inv01 ix5966 (.Y (nx5967), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_3)) ;
    inv01 ix5968 (.Y (nx5969), .A (CacheWindow_4__1__1)) ;
    mux21 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix141 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_3), .A0 (
          nx5971), .A1 (nx5973), .S0 (nx8213)) ;
    inv01 ix5970 (.Y (nx5971), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_4)) ;
    inv01 ix5972 (.Y (nx5973), .A (CacheWindow_4__1__2)) ;
    mux21 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix149 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_4), .A0 (
          nx5975), .A1 (nx5977), .S0 (nx8213)) ;
    inv01 ix5974 (.Y (nx5975), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_5)) ;
    inv01 ix5976 (.Y (nx5977), .A (CacheWindow_4__1__3)) ;
    mux21 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix157 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_5), .A0 (
          nx5979), .A1 (nx5981), .S0 (nx8213)) ;
    inv01 ix5978 (.Y (nx5979), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_6)) ;
    inv01 ix5980 (.Y (nx5981), .A (CacheWindow_4__1__4)) ;
    mux21 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix165 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_6), .A0 (
          nx5983), .A1 (nx5985), .S0 (nx8213)) ;
    inv01 ix5982 (.Y (nx5983), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_7)) ;
    inv01 ix5984 (.Y (nx5985), .A (CacheWindow_4__1__5)) ;
    mux21 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix173 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_7), .A0 (
          nx5987), .A1 (nx5989), .S0 (nx8215)) ;
    inv01 ix5986 (.Y (nx5987), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_8)) ;
    inv01 ix5988 (.Y (nx5989), .A (CacheWindow_4__1__6)) ;
    mux21 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix181 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_8), .A0 (
          nx5991), .A1 (nx5993), .S0 (nx8215)) ;
    inv01 ix5990 (.Y (nx5991), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_9)) ;
    inv01 ix5992 (.Y (nx5993), .A (CacheWindow_4__1__7)) ;
    nor02_2x CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix89 (.Y (
             CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_9), .A0 (
             nx8215), .A1 (nx5995)) ;
    inv01 ix5994 (.Y (nx5995), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_10)) ;
    nor02_2x CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix93 (.Y (
             CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_10), .A0 (
             nx8215), .A1 (nx5997)) ;
    inv01 ix5996 (.Y (nx5997), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_11)) ;
    nor02_2x CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix97 (.Y (
             CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_11), .A0 (
             nx8215), .A1 (nx5999)) ;
    inv01 ix5998 (.Y (nx5999), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_12)) ;
    nor02_2x CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix101 (.Y (
             CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_12), .A0 (
             nx8215), .A1 (nx6001)) ;
    inv01 ix6000 (.Y (nx6001), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_13)) ;
    nor02_2x CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix105 (.Y (
             CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_13), .A0 (
             nx8215), .A1 (nx6003)) ;
    inv01 ix6002 (.Y (nx6003), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_14)) ;
    nor02_2x CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix109 (.Y (
             CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_14), .A0 (
             nx8217), .A1 (nx6005)) ;
    inv01 ix6004 (.Y (nx6005), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_15)) ;
    nor02_2x CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix113 (.Y (
             CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_15), .A0 (
             nx8217), .A1 (nx6007)) ;
    inv01 ix6006 (.Y (nx6007), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_16)) ;
    nor02_2x CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix117 (.Y (
             CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_16), .A0 (
             nx8217), .A1 (nx6007)) ;
    mux21 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix189 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothOperand_0), .A0 (nx6009), .A1 (
          nx6011), .S0 (nx8205)) ;
    inv01 ix6008 (.Y (nx6009), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_0)) ;
    inv01 ix6010 (.Y (nx6011), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_0)) ;
    mux21 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix197 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothOperand_1), .A0 (nx6013), .A1 (
          nx6015), .S0 (nx8205)) ;
    inv01 ix6012 (.Y (nx6013), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_1)) ;
    inv01 ix6014 (.Y (nx6015), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_1)) ;
    mux21 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix205 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothOperand_2), .A0 (nx6017), .A1 (
          nx6019), .S0 (nx8205)) ;
    inv01 ix6016 (.Y (nx6017), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_2)) ;
    inv01 ix6018 (.Y (nx6019), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_2)) ;
    mux21 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix213 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothOperand_3), .A0 (nx6021), .A1 (
          nx6023), .S0 (nx8205)) ;
    inv01 ix6020 (.Y (nx6021), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_3)) ;
    inv01 ix6022 (.Y (nx6023), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_3)) ;
    mux21 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix221 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothOperand_4), .A0 (nx6025), .A1 (
          nx6027), .S0 (nx8205)) ;
    inv01 ix6024 (.Y (nx6025), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_4)) ;
    inv01 ix6026 (.Y (nx6027), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_4)) ;
    mux21 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix229 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothOperand_5), .A0 (nx6029), .A1 (
          nx6031), .S0 (nx8207)) ;
    inv01 ix6028 (.Y (nx6029), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_5)) ;
    inv01 ix6030 (.Y (nx6031), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_5)) ;
    mux21 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix237 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothOperand_6), .A0 (nx6033), .A1 (
          nx6035), .S0 (nx8207)) ;
    inv01 ix6032 (.Y (nx6033), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_6)) ;
    inv01 ix6034 (.Y (nx6035), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_6)) ;
    mux21 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix245 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothOperand_7), .A0 (nx6037), .A1 (
          nx6039), .S0 (nx8207)) ;
    inv01 ix6036 (.Y (nx6037), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_7)) ;
    inv01 ix6038 (.Y (nx6039), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_7)) ;
    mux21 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix253 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothOperand_8), .A0 (nx6041), .A1 (
          nx6043), .S0 (nx8207)) ;
    inv01 ix6040 (.Y (nx6041), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_8)) ;
    inv01 ix6042 (.Y (nx6043), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_8)) ;
    mux21 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix261 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothOperand_9), .A0 (nx6045), .A1 (
          nx6047), .S0 (nx8207)) ;
    inv01 ix6044 (.Y (nx6045), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_9)) ;
    inv01 ix6046 (.Y (nx6047), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_9)) ;
    mux21 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix269 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothOperand_10), .A0 (nx6049), .A1 (
          nx6051), .S0 (nx8207)) ;
    inv01 ix6048 (.Y (nx6049), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_10)) ;
    inv01 ix6050 (.Y (nx6051), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_10)) ;
    mux21 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix277 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothOperand_11), .A0 (nx6053), .A1 (
          nx6055), .S0 (nx8207)) ;
    inv01 ix6052 (.Y (nx6053), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_11)) ;
    inv01 ix6054 (.Y (nx6055), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_11)) ;
    mux21 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix285 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothOperand_12), .A0 (nx6057), .A1 (
          nx6059), .S0 (nx8209)) ;
    inv01 ix6056 (.Y (nx6057), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_12)) ;
    inv01 ix6058 (.Y (nx6059), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_12)) ;
    mux21 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix293 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothOperand_13), .A0 (nx6061), .A1 (
          nx6063), .S0 (nx8209)) ;
    inv01 ix6060 (.Y (nx6061), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_13)) ;
    inv01 ix6062 (.Y (nx6063), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_13)) ;
    mux21 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix301 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothOperand_14), .A0 (nx6065), .A1 (
          nx6067), .S0 (nx8209)) ;
    inv01 ix6064 (.Y (nx6065), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_14)) ;
    inv01 ix6066 (.Y (nx6067), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_14)) ;
    mux21 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix309 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothOperand_15), .A0 (nx6069), .A1 (
          nx6071), .S0 (nx8209)) ;
    inv01 ix6068 (.Y (nx6069), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_15)) ;
    inv01 ix6070 (.Y (nx6071), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_15)) ;
    mux21 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix317 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BoothOperand_16), .A0 (nx6073), .A1 (
          nx6075), .S0 (nx8209)) ;
    inv01 ix6072 (.Y (nx6073), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_16)) ;
    inv01 ix6074 (.Y (nx6075), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_16)) ;
    xnor2 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix321 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_AddPToBoothOperand), .A0 (nx8209), .A1 (
          nx5941)) ;
    oai32 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix393 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .A0 (
          nx8605), .A1 (RST), .A2 (nx8219), .B0 (nx6011), .B1 (nx6079)) ;
    oai32 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix403 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .A0 (
          nx8605), .A1 (RST), .A2 (nx8219), .B0 (nx6015), .B1 (nx6079)) ;
    oai32 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix413 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .A0 (
          nx8605), .A1 (RST), .A2 (nx8219), .B0 (nx6019), .B1 (nx6079)) ;
    oai32 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix423 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .A0 (
          nx8605), .A1 (RST), .A2 (nx8219), .B0 (nx6023), .B1 (nx6079)) ;
    oai32 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix433 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .A0 (
          nx8605), .A1 (RST), .A2 (nx8219), .B0 (nx6027), .B1 (nx6079)) ;
    oai32 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix443 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .A0 (
          nx8605), .A1 (RST), .A2 (nx8219), .B0 (nx6031), .B1 (nx6079)) ;
    oai32 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix453 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .A0 (
          nx8605), .A1 (RST), .A2 (nx8221), .B0 (nx6035), .B1 (nx6079)) ;
    oai32 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix463 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .A0 (
          nx8607), .A1 (RST), .A2 (nx8221), .B0 (nx6039), .B1 (nx6081)) ;
    oai32 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix473 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .A0 (
          nx8607), .A1 (RST), .A2 (nx8221), .B0 (nx6043), .B1 (nx6081)) ;
    oai32 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix483 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .A0 (
          nx6083), .A1 (RST), .A2 (nx8221), .B0 (nx6047), .B1 (nx6081)) ;
    inv01 ix6082 (.Y (nx6083), .A (CacheFilter_4__1__0)) ;
    oai32 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix493 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .A0 (
          nx6085), .A1 (RST), .A2 (nx8221), .B0 (nx6051), .B1 (nx6081)) ;
    inv01 ix6084 (.Y (nx6085), .A (CacheFilter_4__1__1)) ;
    oai32 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix503 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .A0 (
          nx6087), .A1 (RST), .A2 (nx8221), .B0 (nx6055), .B1 (nx6081)) ;
    inv01 ix6086 (.Y (nx6087), .A (CacheFilter_4__1__2)) ;
    oai32 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix513 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .A0 (
          nx6089), .A1 (RST), .A2 (nx8221), .B0 (nx6059), .B1 (nx6081)) ;
    inv01 ix6088 (.Y (nx6089), .A (CacheFilter_4__1__3)) ;
    oai32 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix523 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .A0 (
          nx6091), .A1 (RST), .A2 (nx8223), .B0 (nx6063), .B1 (nx6081)) ;
    inv01 ix6090 (.Y (nx6091), .A (CacheFilter_4__1__4)) ;
    oai32 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix533 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .A0 (
          nx6093), .A1 (RST), .A2 (nx8223), .B0 (nx6067), .B1 (nx6095)) ;
    inv01 ix6092 (.Y (nx6093), .A (CacheFilter_4__1__5)) ;
    inv01 ix6094 (.Y (nx6095), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566)) ;
    oai32 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix543 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .A0 (
          nx6097), .A1 (RST), .A2 (nx8223), .B0 (nx6071), .B1 (nx6095)) ;
    inv01 ix6096 (.Y (nx6097), .A (CacheFilter_4__1__6)) ;
    oai32 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix553 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .A0 (
          nx6099), .A1 (RST), .A2 (nx8223), .B0 (nx6075), .B1 (nx6095)) ;
    inv01 ix6098 (.Y (nx6099), .A (CacheFilter_4__1__7)) ;
    nand02_2x CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix633 (.Y (
              nx6079), .A0 (nx7373), .A1 (nx8223)) ;
    nand02_2x CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix635 (.Y (
              nx6081), .A0 (nx7373), .A1 (nx8223)) ;
    oai32 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix393 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .A0 (
          nx8607), .A1 (RST), .A2 (nx8225), .B0 (nx6009), .B1 (nx6101)) ;
    oai32 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix403 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .A0 (
          nx8607), .A1 (RST), .A2 (nx8225), .B0 (nx6013), .B1 (nx6101)) ;
    oai32 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix413 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .A0 (
          nx8607), .A1 (RST), .A2 (nx8225), .B0 (nx6017), .B1 (nx6101)) ;
    oai32 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix423 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .A0 (
          nx8607), .A1 (RST), .A2 (nx8225), .B0 (nx6021), .B1 (nx6101)) ;
    oai32 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix433 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .A0 (
          nx8607), .A1 (RST), .A2 (nx8225), .B0 (nx6025), .B1 (nx6101)) ;
    oai32 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix443 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .A0 (
          nx8609), .A1 (RST), .A2 (nx8225), .B0 (nx6029), .B1 (nx6101)) ;
    oai32 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix453 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .A0 (
          nx8609), .A1 (RST), .A2 (nx8227), .B0 (nx6033), .B1 (nx6101)) ;
    oai32 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix463 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .A0 (
          nx8609), .A1 (RST), .A2 (nx8227), .B0 (nx6037), .B1 (nx6103)) ;
    oai32 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix473 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .A0 (
          nx8609), .A1 (RST), .A2 (nx8227), .B0 (nx6041), .B1 (nx6103)) ;
    oai32 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix483 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .A0 (
          nx6083), .A1 (RST), .A2 (nx8227), .B0 (nx6045), .B1 (nx6103)) ;
    oai32 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix493 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .A0 (
          nx6105), .A1 (RST), .A2 (nx8227), .B0 (nx6049), .B1 (nx6103)) ;
    inv01 ix6104 (.Y (nx6105), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_10)) ;
    oai32 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix503 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .A0 (
          nx6107), .A1 (RST), .A2 (nx8227), .B0 (nx6053), .B1 (nx6103)) ;
    inv01 ix6106 (.Y (nx6107), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_11)) ;
    oai32 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix513 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .A0 (
          nx6109), .A1 (RST), .A2 (nx8227), .B0 (nx6057), .B1 (nx6103)) ;
    inv01 ix6108 (.Y (nx6109), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_12)) ;
    oai32 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix523 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .A0 (
          nx6111), .A1 (RST), .A2 (nx8229), .B0 (nx6061), .B1 (nx6103)) ;
    inv01 ix6110 (.Y (nx6111), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_13)) ;
    oai32 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix533 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .A0 (
          nx6113), .A1 (RST), .A2 (nx8229), .B0 (nx6065), .B1 (nx6115)) ;
    inv01 ix6112 (.Y (nx6113), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_14)) ;
    inv01 ix6114 (.Y (nx6115), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566)) ;
    oai32 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix543 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .A0 (
          nx6117), .A1 (RST), .A2 (nx8229), .B0 (nx6069), .B1 (nx6115)) ;
    inv01 ix6116 (.Y (nx6117), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_15)) ;
    oai32 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix553 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .A0 (
          nx6119), .A1 (RST), .A2 (nx8229), .B0 (nx6073), .B1 (nx6115)) ;
    inv01 ix6118 (.Y (nx6119), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_16)) ;
    nand02_2x CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix633 (.Y (
              nx6101), .A0 (nx7373), .A1 (nx8229)) ;
    nand02_2x CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix635 (.Y (
              nx6103), .A0 (nx7373), .A1 (nx8229)) ;
    oai32 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix393 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .A0 (
          nx6121), .A1 (RST), .A2 (nx8231), .B0 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_nx384), .B1 (nx6123)) ;
    inv01 ix6120 (.Y (nx6121), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_0)) ;
    oai32 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix403 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .A0 (
          nx6125), .A1 (RST), .A2 (nx8231), .B0 (nx5941), .B1 (nx6123)) ;
    inv01 ix6124 (.Y (nx6125), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_1)) ;
    oai32 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix413 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .A0 (
          nx6127), .A1 (RST), .A2 (nx8231), .B0 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx387), .B1 (nx6123)) ;
    inv01 ix6126 (.Y (nx6127), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_2)) ;
    oai32 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix423 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .A0 (
          nx6129), .A1 (RST), .A2 (nx8231), .B0 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx399), .B1 (nx6123)) ;
    inv01 ix6128 (.Y (nx6129), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_3)) ;
    oai32 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix433 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .A0 (
          nx6131), .A1 (RST), .A2 (nx8231), .B0 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx409), .B1 (nx6123)) ;
    inv01 ix6130 (.Y (nx6131), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_4)) ;
    oai32 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix443 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .A0 (
          nx6133), .A1 (RST), .A2 (nx8231), .B0 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx419), .B1 (nx6123)) ;
    inv01 ix6132 (.Y (nx6133), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_5)) ;
    oai32 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix453 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .A0 (
          nx6135), .A1 (RST), .A2 (nx8231), .B0 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx429), .B1 (nx6123)) ;
    inv01 ix6134 (.Y (nx6135), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_6)) ;
    oai32 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix463 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .A0 (
          nx6137), .A1 (RST), .A2 (nx8233), .B0 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx439), .B1 (nx6139)) ;
    inv01 ix6136 (.Y (nx6137), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_7)) ;
    oai32 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix473 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .A0 (
          nx6141), .A1 (RST), .A2 (nx8233), .B0 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx449), .B1 (nx6139)) ;
    inv01 ix6140 (.Y (nx6141), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_8)) ;
    oai32 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix483 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .A0 (
          nx6143), .A1 (RST), .A2 (nx8233), .B0 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx469), .B1 (nx6139)) ;
    inv01 ix6142 (.Y (nx6143), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_9)) ;
    oai32 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix493 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .A0 (
          nx6145), .A1 (RST), .A2 (nx8233), .B0 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx477), .B1 (nx6139)) ;
    inv01 ix6144 (.Y (nx6145), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_10)) ;
    oai32 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix503 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .A0 (
          nx6147), .A1 (RST), .A2 (nx8233), .B0 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx485), .B1 (nx6139)) ;
    inv01 ix6146 (.Y (nx6147), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_11)) ;
    oai32 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix513 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .A0 (
          nx6149), .A1 (RST), .A2 (nx8233), .B0 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx493), .B1 (nx6139)) ;
    inv01 ix6148 (.Y (nx6149), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_12)) ;
    oai32 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix523 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .A0 (
          nx6151), .A1 (RST), .A2 (nx8233), .B0 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx501), .B1 (nx6139)) ;
    inv01 ix6150 (.Y (nx6151), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_13)) ;
    oai32 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix533 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .A0 (
          nx6153), .A1 (RST), .A2 (nx8235), .B0 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx509), .B1 (nx6155)) ;
    inv01 ix6152 (.Y (nx6153), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_14)) ;
    inv01 ix6154 (.Y (nx6155), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566)) ;
    oai32 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix543 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .A0 (
          nx6157), .A1 (RST), .A2 (nx8235), .B0 (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_nx517), .B1 (nx6155)) ;
    inv01 ix6156 (.Y (nx6157), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_15)) ;
    oai32 CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix553 (.Y (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .A0 (
          nx6159), .A1 (RST), .A2 (nx8235), .B0 (nx5957), .B1 (nx6155)) ;
    inv01 ix6158 (.Y (nx6159), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_16)) ;
    nand02_2x CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix633 (.Y (
              nx6123), .A0 (nx7373), .A1 (nx8235)) ;
    nand02_2x CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix635 (.Y (
              nx6139), .A0 (nx7373), .A1 (nx8235)) ;
    mux21 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix404 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx403), .A0 (nx6161), .A1 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_2), .S0 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx395)) ;
    inv01 ix6160 (.Y (nx6161), .A (CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx391)) ;
    mux21 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix414 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx413), .A0 (nx6163), .A1 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_3), .S0 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx405)) ;
    inv01 ix6162 (.Y (nx6163), .A (CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx403)) ;
    mux21 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix424 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx423), .A0 (nx6165), .A1 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_4), .S0 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx415)) ;
    inv01 ix6164 (.Y (nx6165), .A (CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx413)) ;
    mux21 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix434 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx433), .A0 (nx6167), .A1 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_5), .S0 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx425)) ;
    inv01 ix6166 (.Y (nx6167), .A (CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx423)) ;
    mux21 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix444 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx443), .A0 (nx6169), .A1 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_6), .S0 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx435)) ;
    inv01 ix6168 (.Y (nx6169), .A (CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx433)) ;
    mux21 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix454 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx453), .A0 (nx6171), .A1 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_7), .S0 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx445)) ;
    inv01 ix6170 (.Y (nx6171), .A (CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx443)) ;
    mux21 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix462 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx461), .A0 (nx6173), .A1 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_8), .S0 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx455)) ;
    inv01 ix6172 (.Y (nx6173), .A (CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx453)) ;
    mux21 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix468 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx467), .A0 (nx6175), .A1 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_9), .S0 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx463)) ;
    inv01 ix6174 (.Y (nx6175), .A (CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx461)) ;
    mux21 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix476 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx475), .A0 (nx6177), .A1 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_10), .S0 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx471)) ;
    inv01 ix6176 (.Y (nx6177), .A (CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx467)) ;
    mux21 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix484 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx483), .A0 (nx6179), .A1 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_11), .S0 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx479)) ;
    inv01 ix6178 (.Y (nx6179), .A (CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx475)) ;
    mux21 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix492 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx491), .A0 (nx6181), .A1 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_12), .S0 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx487)) ;
    inv01 ix6180 (.Y (nx6181), .A (CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx483)) ;
    mux21 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix500 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx499), .A0 (nx6183), .A1 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_13), .S0 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx495)) ;
    inv01 ix6182 (.Y (nx6183), .A (CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx491)) ;
    mux21 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix508 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx507), .A0 (nx6185), .A1 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_14), .S0 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx503)) ;
    inv01 ix6184 (.Y (nx6185), .A (CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx499)) ;
    mux21 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix516 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx515), .A0 (nx6187), .A1 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_15), .S0 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx511)) ;
    inv01 ix6186 (.Y (nx6187), .A (CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx507)) ;
    mux21 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix161 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_1), .A0 (nx6189), .A1 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx379), .S0 (nx8239)) ;
    inv01 ix6188 (.Y (nx6189), .A (CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_1)) ;
    mux21 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix181 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_2), .A0 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx387), .A1 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx389), .S0 (nx8239)) ;
    mux21 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix201 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_3), .A0 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx399), .A1 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx401), .S0 (nx8239)) ;
    mux21 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix221 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_4), .A0 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx409), .A1 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx411), .S0 (nx8239)) ;
    mux21 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix241 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_5), .A0 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx419), .A1 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx421), .S0 (nx8239)) ;
    mux21 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix261 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_6), .A0 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx429), .A1 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx431), .S0 (nx8239)) ;
    mux21 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix281 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_7), .A0 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx439), .A1 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx441), .S0 (nx8239)) ;
    mux21 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix301 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_8), .A0 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx449), .A1 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx451), .S0 (nx8241)) ;
    mux21 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix321 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_9), .A0 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx469), .A1 (nx6191), .S0 (nx8241)) ;
    inv01 ix6190 (.Y (nx6191), .A (CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx316)) ;
    mux21 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix341 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_10), .A0 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx477), .A1 (nx6193), .S0 (nx8241)) ;
    inv01 ix6192 (.Y (nx6193), .A (CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx336)) ;
    mux21 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix361 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_11), .A0 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx485), .A1 (nx6195), .S0 (nx8241)) ;
    inv01 ix6194 (.Y (nx6195), .A (CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx356)) ;
    mux21 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix381 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_12), .A0 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx493), .A1 (nx6197), .S0 (nx8241)) ;
    inv01 ix6196 (.Y (nx6197), .A (CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx376)) ;
    mux21 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix401 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_13), .A0 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx501), .A1 (nx6199), .S0 (nx8241)) ;
    inv01 ix6198 (.Y (nx6199), .A (CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx396)) ;
    mux21 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix421 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_14), .A0 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx509), .A1 (nx6201), .S0 (nx8241)) ;
    inv01 ix6200 (.Y (nx6201), .A (CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx416)) ;
    mux21 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix441 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_15), .A0 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx517), .A1 (nx6203), .S0 (nx8243)) ;
    inv01 ix6202 (.Y (nx6203), .A (CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx436)) ;
    mux21 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_ix461 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_16), .A0 (nx6205), 
          .A1 (nx6207), .S0 (nx8243)) ;
    inv01 ix6204 (.Y (nx6205), .A (CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothP_16)
          ) ;
    inv01 ix6206 (.Y (nx6207), .A (CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx456)) ;
    nor02_2x CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix81 (.Y (
             CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_nx80), .A0 (Instr), .A1 (
             nx7299)) ;
    nor02_2x CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix319 (.Y (
             CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642), .A0 (
             CALCULATOR_Start_dup_1326), .A1 (
             CALCULATOR_CalculatingBooth_dup_1315)) ;
    nor02_2x CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix85 (.Y (
             CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_0), .A0 (
             nx8253), .A1 (nx6209)) ;
    inv01 ix6208 (.Y (nx6209), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_1)) ;
    mux21 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix125 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_1), .A0 (
          nx6211), .A1 (nx6213), .S0 (nx8253)) ;
    inv01 ix6210 (.Y (nx6211), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_2)) ;
    inv01 ix6212 (.Y (nx6213), .A (CacheWindow_4__2__0)) ;
    mux21 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix133 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_2), .A0 (
          nx6215), .A1 (nx6217), .S0 (nx8253)) ;
    inv01 ix6214 (.Y (nx6215), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_3)) ;
    inv01 ix6216 (.Y (nx6217), .A (CacheWindow_4__2__1)) ;
    mux21 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix141 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_3), .A0 (
          nx6219), .A1 (nx6221), .S0 (nx8253)) ;
    inv01 ix6218 (.Y (nx6219), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_4)) ;
    inv01 ix6220 (.Y (nx6221), .A (CacheWindow_4__2__2)) ;
    mux21 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix149 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_4), .A0 (
          nx6223), .A1 (nx6225), .S0 (nx8253)) ;
    inv01 ix6222 (.Y (nx6223), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_5)) ;
    inv01 ix6224 (.Y (nx6225), .A (CacheWindow_4__2__3)) ;
    mux21 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix157 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_5), .A0 (
          nx6227), .A1 (nx6229), .S0 (nx8253)) ;
    inv01 ix6226 (.Y (nx6227), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_6)) ;
    inv01 ix6228 (.Y (nx6229), .A (CacheWindow_4__2__4)) ;
    mux21 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix165 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_6), .A0 (
          nx6231), .A1 (nx6233), .S0 (nx8253)) ;
    inv01 ix6230 (.Y (nx6231), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_7)) ;
    inv01 ix6232 (.Y (nx6233), .A (CacheWindow_4__2__5)) ;
    mux21 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix173 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_7), .A0 (
          nx6235), .A1 (nx6237), .S0 (nx8255)) ;
    inv01 ix6234 (.Y (nx6235), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_8)) ;
    inv01 ix6236 (.Y (nx6237), .A (CacheWindow_4__2__6)) ;
    mux21 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix181 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_8), .A0 (
          nx6239), .A1 (nx6241), .S0 (nx8255)) ;
    inv01 ix6238 (.Y (nx6239), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_9)) ;
    inv01 ix6240 (.Y (nx6241), .A (CacheWindow_4__2__7)) ;
    nor02_2x CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix89 (.Y (
             CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_9), .A0 (
             nx8255), .A1 (nx6243)) ;
    inv01 ix6242 (.Y (nx6243), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_10)) ;
    nor02_2x CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix93 (.Y (
             CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_10), .A0 (
             nx8255), .A1 (nx6245)) ;
    inv01 ix6244 (.Y (nx6245), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_11)) ;
    nor02_2x CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix97 (.Y (
             CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_11), .A0 (
             nx8255), .A1 (nx6247)) ;
    inv01 ix6246 (.Y (nx6247), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_12)) ;
    nor02_2x CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix101 (.Y (
             CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_12), .A0 (
             nx8255), .A1 (nx6249)) ;
    inv01 ix6248 (.Y (nx6249), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_13)) ;
    nor02_2x CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix105 (.Y (
             CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_13), .A0 (
             nx8255), .A1 (nx6251)) ;
    inv01 ix6250 (.Y (nx6251), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_14)) ;
    nor02_2x CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix109 (.Y (
             CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_14), .A0 (
             nx8257), .A1 (nx6253)) ;
    inv01 ix6252 (.Y (nx6253), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_15)) ;
    nor02_2x CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix113 (.Y (
             CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_15), .A0 (
             nx8257), .A1 (nx6255)) ;
    inv01 ix6254 (.Y (nx6255), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_16)) ;
    nor02_2x CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix117 (.Y (
             CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_16), .A0 (
             nx8257), .A1 (nx6255)) ;
    mux21 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix189 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothOperand_0), .A0 (nx6257), .A1 (
          nx6259), .S0 (nx8245)) ;
    inv01 ix6256 (.Y (nx6257), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_0)) ;
    inv01 ix6258 (.Y (nx6259), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_0)) ;
    mux21 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix197 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothOperand_1), .A0 (nx6261), .A1 (
          nx6263), .S0 (nx8245)) ;
    inv01 ix6260 (.Y (nx6261), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_1)) ;
    inv01 ix6262 (.Y (nx6263), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_1)) ;
    mux21 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix205 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothOperand_2), .A0 (nx6265), .A1 (
          nx6267), .S0 (nx8245)) ;
    inv01 ix6264 (.Y (nx6265), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_2)) ;
    inv01 ix6266 (.Y (nx6267), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_2)) ;
    mux21 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix213 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothOperand_3), .A0 (nx6269), .A1 (
          nx6271), .S0 (nx8245)) ;
    inv01 ix6268 (.Y (nx6269), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_3)) ;
    inv01 ix6270 (.Y (nx6271), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_3)) ;
    mux21 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix221 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothOperand_4), .A0 (nx6273), .A1 (
          nx6275), .S0 (nx8245)) ;
    inv01 ix6272 (.Y (nx6273), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_4)) ;
    inv01 ix6274 (.Y (nx6275), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_4)) ;
    mux21 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix229 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothOperand_5), .A0 (nx6277), .A1 (
          nx6279), .S0 (nx8247)) ;
    inv01 ix6276 (.Y (nx6277), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_5)) ;
    inv01 ix6278 (.Y (nx6279), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_5)) ;
    mux21 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix237 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothOperand_6), .A0 (nx6281), .A1 (
          nx6283), .S0 (nx8247)) ;
    inv01 ix6280 (.Y (nx6281), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_6)) ;
    inv01 ix6282 (.Y (nx6283), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_6)) ;
    mux21 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix245 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothOperand_7), .A0 (nx6285), .A1 (
          nx6287), .S0 (nx8247)) ;
    inv01 ix6284 (.Y (nx6285), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_7)) ;
    inv01 ix6286 (.Y (nx6287), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_7)) ;
    mux21 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix253 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothOperand_8), .A0 (nx6289), .A1 (
          nx6291), .S0 (nx8247)) ;
    inv01 ix6288 (.Y (nx6289), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_8)) ;
    inv01 ix6290 (.Y (nx6291), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_8)) ;
    mux21 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix261 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothOperand_9), .A0 (nx6293), .A1 (
          nx6295), .S0 (nx8247)) ;
    inv01 ix6292 (.Y (nx6293), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_9)) ;
    inv01 ix6294 (.Y (nx6295), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_9)) ;
    mux21 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix269 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothOperand_10), .A0 (nx6297), .A1 (
          nx6299), .S0 (nx8247)) ;
    inv01 ix6296 (.Y (nx6297), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_10)) ;
    inv01 ix6298 (.Y (nx6299), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_10)) ;
    mux21 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix277 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothOperand_11), .A0 (nx6301), .A1 (
          nx6303), .S0 (nx8247)) ;
    inv01 ix6300 (.Y (nx6301), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_11)) ;
    inv01 ix6302 (.Y (nx6303), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_11)) ;
    mux21 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix285 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothOperand_12), .A0 (nx6305), .A1 (
          nx6307), .S0 (nx8249)) ;
    inv01 ix6304 (.Y (nx6305), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_12)) ;
    inv01 ix6306 (.Y (nx6307), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_12)) ;
    mux21 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix293 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothOperand_13), .A0 (nx6309), .A1 (
          nx6311), .S0 (nx8249)) ;
    inv01 ix6308 (.Y (nx6309), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_13)) ;
    inv01 ix6310 (.Y (nx6311), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_13)) ;
    mux21 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix301 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothOperand_14), .A0 (nx6313), .A1 (
          nx6315), .S0 (nx8249)) ;
    inv01 ix6312 (.Y (nx6313), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_14)) ;
    inv01 ix6314 (.Y (nx6315), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_14)) ;
    mux21 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix309 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothOperand_15), .A0 (nx6317), .A1 (
          nx6319), .S0 (nx8249)) ;
    inv01 ix6316 (.Y (nx6317), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_15)) ;
    inv01 ix6318 (.Y (nx6319), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_15)) ;
    mux21 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix317 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BoothOperand_16), .A0 (nx6321), .A1 (
          nx6323), .S0 (nx8249)) ;
    inv01 ix6320 (.Y (nx6321), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_16)) ;
    inv01 ix6322 (.Y (nx6323), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_16)) ;
    xnor2 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix321 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_AddPToBoothOperand), .A0 (nx8249), .A1 (
          nx6189)) ;
    oai32 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix393 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .A0 (
          nx8611), .A1 (RST), .A2 (nx8259), .B0 (nx6259), .B1 (nx6327)) ;
    oai32 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix403 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .A0 (
          nx8611), .A1 (RST), .A2 (nx8259), .B0 (nx6263), .B1 (nx6327)) ;
    oai32 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix413 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .A0 (
          nx8611), .A1 (RST), .A2 (nx8259), .B0 (nx6267), .B1 (nx6327)) ;
    oai32 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix423 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .A0 (
          nx8611), .A1 (RST), .A2 (nx8259), .B0 (nx6271), .B1 (nx6327)) ;
    oai32 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix433 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .A0 (
          nx8611), .A1 (RST), .A2 (nx8259), .B0 (nx6275), .B1 (nx6327)) ;
    oai32 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix443 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .A0 (
          nx8611), .A1 (RST), .A2 (nx8259), .B0 (nx6279), .B1 (nx6327)) ;
    oai32 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix453 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .A0 (
          nx8611), .A1 (RST), .A2 (nx8261), .B0 (nx6283), .B1 (nx6327)) ;
    oai32 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix463 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .A0 (
          nx8613), .A1 (RST), .A2 (nx8261), .B0 (nx6287), .B1 (nx6329)) ;
    oai32 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix473 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .A0 (
          nx8613), .A1 (RST), .A2 (nx8261), .B0 (nx6291), .B1 (nx6329)) ;
    oai32 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix483 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .A0 (
          nx6331), .A1 (RST), .A2 (nx8261), .B0 (nx6295), .B1 (nx6329)) ;
    inv01 ix6330 (.Y (nx6331), .A (CacheFilter_4__2__0)) ;
    oai32 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix493 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .A0 (
          nx6333), .A1 (RST), .A2 (nx8261), .B0 (nx6299), .B1 (nx6329)) ;
    inv01 ix6332 (.Y (nx6333), .A (CacheFilter_4__2__1)) ;
    oai32 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix503 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .A0 (
          nx6335), .A1 (RST), .A2 (nx8261), .B0 (nx6303), .B1 (nx6329)) ;
    inv01 ix6334 (.Y (nx6335), .A (CacheFilter_4__2__2)) ;
    oai32 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix513 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .A0 (
          nx6337), .A1 (RST), .A2 (nx8261), .B0 (nx6307), .B1 (nx6329)) ;
    inv01 ix6336 (.Y (nx6337), .A (CacheFilter_4__2__3)) ;
    oai32 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix523 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .A0 (
          nx6339), .A1 (RST), .A2 (nx8263), .B0 (nx6311), .B1 (nx6329)) ;
    inv01 ix6338 (.Y (nx6339), .A (CacheFilter_4__2__4)) ;
    oai32 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix533 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .A0 (
          nx6341), .A1 (RST), .A2 (nx8263), .B0 (nx6315), .B1 (nx6343)) ;
    inv01 ix6340 (.Y (nx6341), .A (CacheFilter_4__2__5)) ;
    inv01 ix6342 (.Y (nx6343), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566)) ;
    oai32 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix543 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .A0 (
          nx6345), .A1 (RST), .A2 (nx8263), .B0 (nx6319), .B1 (nx6343)) ;
    inv01 ix6344 (.Y (nx6345), .A (CacheFilter_4__2__6)) ;
    oai32 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix553 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .A0 (
          nx6347), .A1 (RST), .A2 (nx8263), .B0 (nx6323), .B1 (nx6343)) ;
    inv01 ix6346 (.Y (nx6347), .A (CacheFilter_4__2__7)) ;
    nand02_2x CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix633 (.Y (
              nx6327), .A0 (nx7375), .A1 (nx8263)) ;
    nand02_2x CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix635 (.Y (
              nx6329), .A0 (nx7375), .A1 (nx8263)) ;
    oai32 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix393 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .A0 (
          nx8613), .A1 (RST), .A2 (nx8265), .B0 (nx6257), .B1 (nx6349)) ;
    oai32 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix403 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .A0 (
          nx8613), .A1 (RST), .A2 (nx8265), .B0 (nx6261), .B1 (nx6349)) ;
    oai32 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix413 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .A0 (
          nx8613), .A1 (RST), .A2 (nx8265), .B0 (nx6265), .B1 (nx6349)) ;
    oai32 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix423 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .A0 (
          nx8613), .A1 (RST), .A2 (nx8265), .B0 (nx6269), .B1 (nx6349)) ;
    oai32 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix433 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .A0 (
          nx8613), .A1 (RST), .A2 (nx8265), .B0 (nx6273), .B1 (nx6349)) ;
    oai32 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix443 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .A0 (
          nx8615), .A1 (RST), .A2 (nx8265), .B0 (nx6277), .B1 (nx6349)) ;
    oai32 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix453 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .A0 (
          nx8615), .A1 (RST), .A2 (nx8267), .B0 (nx6281), .B1 (nx6349)) ;
    oai32 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix463 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .A0 (
          nx8615), .A1 (RST), .A2 (nx8267), .B0 (nx6285), .B1 (nx6351)) ;
    oai32 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix473 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .A0 (
          nx8615), .A1 (RST), .A2 (nx8267), .B0 (nx6289), .B1 (nx6351)) ;
    oai32 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix483 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .A0 (
          nx6331), .A1 (RST), .A2 (nx8267), .B0 (nx6293), .B1 (nx6351)) ;
    oai32 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix493 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .A0 (
          nx6353), .A1 (RST), .A2 (nx8267), .B0 (nx6297), .B1 (nx6351)) ;
    inv01 ix6352 (.Y (nx6353), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDin_10)) ;
    oai32 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix503 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .A0 (
          nx6355), .A1 (RST), .A2 (nx8267), .B0 (nx6301), .B1 (nx6351)) ;
    inv01 ix6354 (.Y (nx6355), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDin_11)) ;
    oai32 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix513 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .A0 (
          nx6357), .A1 (RST), .A2 (nx8267), .B0 (nx6305), .B1 (nx6351)) ;
    inv01 ix6356 (.Y (nx6357), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDin_12)) ;
    oai32 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix523 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .A0 (
          nx6359), .A1 (RST), .A2 (nx8269), .B0 (nx6309), .B1 (nx6351)) ;
    inv01 ix6358 (.Y (nx6359), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDin_13)) ;
    oai32 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix533 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .A0 (
          nx6361), .A1 (RST), .A2 (nx8269), .B0 (nx6313), .B1 (nx6363)) ;
    inv01 ix6360 (.Y (nx6361), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDin_14)) ;
    inv01 ix6362 (.Y (nx6363), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566)) ;
    oai32 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix543 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .A0 (
          nx6365), .A1 (RST), .A2 (nx8269), .B0 (nx6317), .B1 (nx6363)) ;
    inv01 ix6364 (.Y (nx6365), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDin_15)) ;
    oai32 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix553 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .A0 (
          nx6367), .A1 (RST), .A2 (nx8269), .B0 (nx6321), .B1 (nx6363)) ;
    inv01 ix6366 (.Y (nx6367), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDin_16)) ;
    nand02_2x CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix633 (.Y (
              nx6349), .A0 (nx7375), .A1 (nx8269)) ;
    nand02_2x CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix635 (.Y (
              nx6351), .A0 (nx7375), .A1 (nx8269)) ;
    oai32 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix393 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .A0 (
          nx6369), .A1 (RST), .A2 (nx8271), .B0 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_nx384), .B1 (nx6371)) ;
    inv01 ix6368 (.Y (nx6369), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_0)) ;
    oai32 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix403 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .A0 (
          nx6373), .A1 (RST), .A2 (nx8271), .B0 (nx6189), .B1 (nx6371)) ;
    inv01 ix6372 (.Y (nx6373), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_1)) ;
    oai32 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix413 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .A0 (
          nx6375), .A1 (RST), .A2 (nx8271), .B0 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx387), .B1 (nx6371)) ;
    inv01 ix6374 (.Y (nx6375), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_2)) ;
    oai32 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix423 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .A0 (
          nx6377), .A1 (RST), .A2 (nx8271), .B0 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx399), .B1 (nx6371)) ;
    inv01 ix6376 (.Y (nx6377), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_3)) ;
    oai32 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix433 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .A0 (
          nx6379), .A1 (RST), .A2 (nx8271), .B0 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx409), .B1 (nx6371)) ;
    inv01 ix6378 (.Y (nx6379), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_4)) ;
    oai32 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix443 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .A0 (
          nx6381), .A1 (RST), .A2 (nx8271), .B0 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx419), .B1 (nx6371)) ;
    inv01 ix6380 (.Y (nx6381), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_5)) ;
    oai32 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix453 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .A0 (
          nx6383), .A1 (RST), .A2 (nx8271), .B0 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx429), .B1 (nx6371)) ;
    inv01 ix6382 (.Y (nx6383), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_6)) ;
    oai32 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix463 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .A0 (
          nx6385), .A1 (RST), .A2 (nx8273), .B0 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx439), .B1 (nx6387)) ;
    inv01 ix6384 (.Y (nx6385), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_7)) ;
    oai32 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix473 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .A0 (
          nx6389), .A1 (RST), .A2 (nx8273), .B0 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx449), .B1 (nx6387)) ;
    inv01 ix6388 (.Y (nx6389), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_8)) ;
    oai32 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix483 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .A0 (
          nx6391), .A1 (RST), .A2 (nx8273), .B0 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx469), .B1 (nx6387)) ;
    inv01 ix6390 (.Y (nx6391), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_9)) ;
    oai32 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix493 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .A0 (
          nx6393), .A1 (RST), .A2 (nx8273), .B0 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx477), .B1 (nx6387)) ;
    inv01 ix6392 (.Y (nx6393), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_10)) ;
    oai32 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix503 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .A0 (
          nx6395), .A1 (RST), .A2 (nx8273), .B0 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx485), .B1 (nx6387)) ;
    inv01 ix6394 (.Y (nx6395), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_11)) ;
    oai32 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix513 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .A0 (
          nx6397), .A1 (RST), .A2 (nx8273), .B0 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx493), .B1 (nx6387)) ;
    inv01 ix6396 (.Y (nx6397), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_12)) ;
    oai32 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix523 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .A0 (
          nx6399), .A1 (RST), .A2 (nx8273), .B0 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx501), .B1 (nx6387)) ;
    inv01 ix6398 (.Y (nx6399), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_13)) ;
    oai32 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix533 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .A0 (
          nx6401), .A1 (RST), .A2 (nx8275), .B0 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx509), .B1 (nx6403)) ;
    inv01 ix6400 (.Y (nx6401), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_14)) ;
    inv01 ix6402 (.Y (nx6403), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566)) ;
    oai32 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix543 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .A0 (
          nx6405), .A1 (RST), .A2 (nx8275), .B0 (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_nx517), .B1 (nx6403)) ;
    inv01 ix6404 (.Y (nx6405), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_15)) ;
    oai32 CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix553 (.Y (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .A0 (
          nx6407), .A1 (RST), .A2 (nx8275), .B0 (nx6205), .B1 (nx6403)) ;
    inv01 ix6406 (.Y (nx6407), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_16)) ;
    nand02_2x CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix633 (.Y (
              nx6371), .A0 (nx7375), .A1 (nx8275)) ;
    nand02_2x CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix635 (.Y (
              nx6387), .A0 (nx7375), .A1 (nx8275)) ;
    mux21 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix404 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx403), .A0 (nx6409), .A1 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_2), .S0 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx395)) ;
    inv01 ix6408 (.Y (nx6409), .A (CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx391)) ;
    mux21 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix414 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx413), .A0 (nx6411), .A1 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_3), .S0 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx405)) ;
    inv01 ix6410 (.Y (nx6411), .A (CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx403)) ;
    mux21 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix424 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx423), .A0 (nx6413), .A1 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_4), .S0 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx415)) ;
    inv01 ix6412 (.Y (nx6413), .A (CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx413)) ;
    mux21 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix434 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx433), .A0 (nx6415), .A1 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_5), .S0 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx425)) ;
    inv01 ix6414 (.Y (nx6415), .A (CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx423)) ;
    mux21 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix444 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx443), .A0 (nx6417), .A1 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_6), .S0 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx435)) ;
    inv01 ix6416 (.Y (nx6417), .A (CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx433)) ;
    mux21 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix454 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx453), .A0 (nx6419), .A1 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_7), .S0 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx445)) ;
    inv01 ix6418 (.Y (nx6419), .A (CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx443)) ;
    mux21 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix462 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx461), .A0 (nx6421), .A1 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_8), .S0 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx455)) ;
    inv01 ix6420 (.Y (nx6421), .A (CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx453)) ;
    mux21 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix468 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx467), .A0 (nx6423), .A1 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_9), .S0 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx463)) ;
    inv01 ix6422 (.Y (nx6423), .A (CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx461)) ;
    mux21 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix476 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx475), .A0 (nx6425), .A1 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_10), .S0 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx471)) ;
    inv01 ix6424 (.Y (nx6425), .A (CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx467)) ;
    mux21 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix484 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx483), .A0 (nx6427), .A1 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_11), .S0 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx479)) ;
    inv01 ix6426 (.Y (nx6427), .A (CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx475)) ;
    mux21 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix492 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx491), .A0 (nx6429), .A1 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_12), .S0 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx487)) ;
    inv01 ix6428 (.Y (nx6429), .A (CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx483)) ;
    mux21 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix500 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx499), .A0 (nx6431), .A1 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_13), .S0 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx495)) ;
    inv01 ix6430 (.Y (nx6431), .A (CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx491)) ;
    mux21 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix508 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx507), .A0 (nx6433), .A1 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_14), .S0 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx503)) ;
    inv01 ix6432 (.Y (nx6433), .A (CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx499)) ;
    mux21 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix516 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx515), .A0 (nx6435), .A1 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_15), .S0 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx511)) ;
    inv01 ix6434 (.Y (nx6435), .A (CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx507)) ;
    mux21 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix161 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_1), .A0 (nx6437), .A1 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx379), .S0 (nx8279)) ;
    inv01 ix6436 (.Y (nx6437), .A (CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_1)) ;
    mux21 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix181 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_2), .A0 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx387), .A1 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx389), .S0 (nx8279)) ;
    mux21 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix201 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_3), .A0 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx399), .A1 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx401), .S0 (nx8279)) ;
    mux21 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix221 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_4), .A0 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx409), .A1 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx411), .S0 (nx8279)) ;
    mux21 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix241 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_5), .A0 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx419), .A1 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx421), .S0 (nx8279)) ;
    mux21 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix261 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_6), .A0 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx429), .A1 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx431), .S0 (nx8279)) ;
    mux21 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix281 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_7), .A0 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx439), .A1 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx441), .S0 (nx8279)) ;
    mux21 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix301 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_8), .A0 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx449), .A1 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx451), .S0 (nx8281)) ;
    mux21 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix321 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_9), .A0 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx469), .A1 (nx6439), .S0 (nx8281)) ;
    inv01 ix6438 (.Y (nx6439), .A (CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx316)) ;
    mux21 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix341 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_10), .A0 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx477), .A1 (nx6441), .S0 (nx8281)) ;
    inv01 ix6440 (.Y (nx6441), .A (CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx336)) ;
    mux21 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix361 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_11), .A0 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx485), .A1 (nx6443), .S0 (nx8281)) ;
    inv01 ix6442 (.Y (nx6443), .A (CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx356)) ;
    mux21 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix381 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_12), .A0 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx493), .A1 (nx6445), .S0 (nx8281)) ;
    inv01 ix6444 (.Y (nx6445), .A (CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx376)) ;
    mux21 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix401 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_13), .A0 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx501), .A1 (nx6447), .S0 (nx8281)) ;
    inv01 ix6446 (.Y (nx6447), .A (CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx396)) ;
    mux21 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix421 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_14), .A0 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx509), .A1 (nx6449), .S0 (nx8281)) ;
    inv01 ix6448 (.Y (nx6449), .A (CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx416)) ;
    mux21 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix441 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_15), .A0 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx517), .A1 (nx6451), .S0 (nx8283)) ;
    inv01 ix6450 (.Y (nx6451), .A (CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx436)) ;
    mux21 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_ix461 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_16), .A0 (nx6453), 
          .A1 (nx6455), .S0 (nx8283)) ;
    inv01 ix6452 (.Y (nx6453), .A (CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothP_16)
          ) ;
    inv01 ix6454 (.Y (nx6455), .A (CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx456)) ;
    nor02_2x CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix81 (.Y (
             CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_nx80), .A0 (Instr), .A1 (
             nx7299)) ;
    nor02_2x CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix319 (.Y (
             CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642), .A0 (
             CALCULATOR_Start_dup_1339), .A1 (
             CALCULATOR_CalculatingBooth_dup_1315)) ;
    nor02_2x CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix85 (.Y (
             CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_0), .A0 (
             nx8293), .A1 (nx6457)) ;
    inv01 ix6456 (.Y (nx6457), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_1)) ;
    mux21 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix125 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_1), .A0 (
          nx6459), .A1 (nx6461), .S0 (nx8293)) ;
    inv01 ix6458 (.Y (nx6459), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_2)) ;
    inv01 ix6460 (.Y (nx6461), .A (CacheWindow_4__3__0)) ;
    mux21 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix133 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_2), .A0 (
          nx6463), .A1 (nx6465), .S0 (nx8293)) ;
    inv01 ix6462 (.Y (nx6463), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_3)) ;
    inv01 ix6464 (.Y (nx6465), .A (CacheWindow_4__3__1)) ;
    mux21 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix141 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_3), .A0 (
          nx6467), .A1 (nx6469), .S0 (nx8293)) ;
    inv01 ix6466 (.Y (nx6467), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_4)) ;
    inv01 ix6468 (.Y (nx6469), .A (CacheWindow_4__3__2)) ;
    mux21 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix149 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_4), .A0 (
          nx6471), .A1 (nx6473), .S0 (nx8293)) ;
    inv01 ix6470 (.Y (nx6471), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_5)) ;
    inv01 ix6472 (.Y (nx6473), .A (CacheWindow_4__3__3)) ;
    mux21 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix157 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_5), .A0 (
          nx6475), .A1 (nx6477), .S0 (nx8293)) ;
    inv01 ix6474 (.Y (nx6475), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_6)) ;
    inv01 ix6476 (.Y (nx6477), .A (CacheWindow_4__3__4)) ;
    mux21 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix165 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_6), .A0 (
          nx6479), .A1 (nx6481), .S0 (nx8293)) ;
    inv01 ix6478 (.Y (nx6479), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_7)) ;
    inv01 ix6480 (.Y (nx6481), .A (CacheWindow_4__3__5)) ;
    mux21 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix173 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_7), .A0 (
          nx6483), .A1 (nx6485), .S0 (nx8295)) ;
    inv01 ix6482 (.Y (nx6483), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_8)) ;
    inv01 ix6484 (.Y (nx6485), .A (CacheWindow_4__3__6)) ;
    mux21 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix181 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_8), .A0 (
          nx6487), .A1 (nx6489), .S0 (nx8295)) ;
    inv01 ix6486 (.Y (nx6487), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_9)) ;
    inv01 ix6488 (.Y (nx6489), .A (CacheWindow_4__3__7)) ;
    nor02_2x CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix89 (.Y (
             CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_9), .A0 (
             nx8295), .A1 (nx6491)) ;
    inv01 ix6490 (.Y (nx6491), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_10)) ;
    nor02_2x CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix93 (.Y (
             CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_10), .A0 (
             nx8295), .A1 (nx6493)) ;
    inv01 ix6492 (.Y (nx6493), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_11)) ;
    nor02_2x CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix97 (.Y (
             CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_11), .A0 (
             nx8295), .A1 (nx6495)) ;
    inv01 ix6494 (.Y (nx6495), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_12)) ;
    nor02_2x CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix101 (.Y (
             CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_12), .A0 (
             nx8295), .A1 (nx6497)) ;
    inv01 ix6496 (.Y (nx6497), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_13)) ;
    nor02_2x CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix105 (.Y (
             CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_13), .A0 (
             nx8295), .A1 (nx6499)) ;
    inv01 ix6498 (.Y (nx6499), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_14)) ;
    nor02_2x CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix109 (.Y (
             CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_14), .A0 (
             nx8297), .A1 (nx6501)) ;
    inv01 ix6500 (.Y (nx6501), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_15)) ;
    nor02_2x CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix113 (.Y (
             CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_15), .A0 (
             nx8297), .A1 (nx6503)) ;
    inv01 ix6502 (.Y (nx6503), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_16)) ;
    nor02_2x CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix117 (.Y (
             CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_16), .A0 (
             nx8297), .A1 (nx6503)) ;
    mux21 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix189 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothOperand_0), .A0 (nx6505), .A1 (
          nx6507), .S0 (nx8285)) ;
    inv01 ix6504 (.Y (nx6505), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_0)) ;
    inv01 ix6506 (.Y (nx6507), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_0)) ;
    mux21 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix197 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothOperand_1), .A0 (nx6509), .A1 (
          nx6511), .S0 (nx8285)) ;
    inv01 ix6508 (.Y (nx6509), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_1)) ;
    inv01 ix6510 (.Y (nx6511), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_1)) ;
    mux21 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix205 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothOperand_2), .A0 (nx6513), .A1 (
          nx6515), .S0 (nx8285)) ;
    inv01 ix6512 (.Y (nx6513), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_2)) ;
    inv01 ix6514 (.Y (nx6515), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_2)) ;
    mux21 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix213 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothOperand_3), .A0 (nx6517), .A1 (
          nx6519), .S0 (nx8285)) ;
    inv01 ix6516 (.Y (nx6517), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_3)) ;
    inv01 ix6518 (.Y (nx6519), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_3)) ;
    mux21 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix221 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothOperand_4), .A0 (nx6521), .A1 (
          nx6523), .S0 (nx8285)) ;
    inv01 ix6520 (.Y (nx6521), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_4)) ;
    inv01 ix6522 (.Y (nx6523), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_4)) ;
    mux21 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix229 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothOperand_5), .A0 (nx6525), .A1 (
          nx6527), .S0 (nx8287)) ;
    inv01 ix6524 (.Y (nx6525), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_5)) ;
    inv01 ix6526 (.Y (nx6527), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_5)) ;
    mux21 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix237 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothOperand_6), .A0 (nx6529), .A1 (
          nx6531), .S0 (nx8287)) ;
    inv01 ix6528 (.Y (nx6529), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_6)) ;
    inv01 ix6530 (.Y (nx6531), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_6)) ;
    mux21 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix245 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothOperand_7), .A0 (nx6533), .A1 (
          nx6535), .S0 (nx8287)) ;
    inv01 ix6532 (.Y (nx6533), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_7)) ;
    inv01 ix6534 (.Y (nx6535), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_7)) ;
    mux21 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix253 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothOperand_8), .A0 (nx6537), .A1 (
          nx6539), .S0 (nx8287)) ;
    inv01 ix6536 (.Y (nx6537), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_8)) ;
    inv01 ix6538 (.Y (nx6539), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_8)) ;
    mux21 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix261 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothOperand_9), .A0 (nx6541), .A1 (
          nx6543), .S0 (nx8287)) ;
    inv01 ix6540 (.Y (nx6541), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_9)) ;
    inv01 ix6542 (.Y (nx6543), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_9)) ;
    mux21 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix269 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothOperand_10), .A0 (nx6545), .A1 (
          nx6547), .S0 (nx8287)) ;
    inv01 ix6544 (.Y (nx6545), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_10)) ;
    inv01 ix6546 (.Y (nx6547), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_10)) ;
    mux21 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix277 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothOperand_11), .A0 (nx6549), .A1 (
          nx6551), .S0 (nx8287)) ;
    inv01 ix6548 (.Y (nx6549), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_11)) ;
    inv01 ix6550 (.Y (nx6551), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_11)) ;
    mux21 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix285 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothOperand_12), .A0 (nx6553), .A1 (
          nx6555), .S0 (nx8289)) ;
    inv01 ix6552 (.Y (nx6553), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_12)) ;
    inv01 ix6554 (.Y (nx6555), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_12)) ;
    mux21 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix293 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothOperand_13), .A0 (nx6557), .A1 (
          nx6559), .S0 (nx8289)) ;
    inv01 ix6556 (.Y (nx6557), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_13)) ;
    inv01 ix6558 (.Y (nx6559), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_13)) ;
    mux21 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix301 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothOperand_14), .A0 (nx6561), .A1 (
          nx6563), .S0 (nx8289)) ;
    inv01 ix6560 (.Y (nx6561), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_14)) ;
    inv01 ix6562 (.Y (nx6563), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_14)) ;
    mux21 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix309 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothOperand_15), .A0 (nx6565), .A1 (
          nx6567), .S0 (nx8289)) ;
    inv01 ix6564 (.Y (nx6565), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_15)) ;
    inv01 ix6566 (.Y (nx6567), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_15)) ;
    mux21 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix317 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BoothOperand_16), .A0 (nx6569), .A1 (
          nx6571), .S0 (nx8289)) ;
    inv01 ix6568 (.Y (nx6569), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_16)) ;
    inv01 ix6570 (.Y (nx6571), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_16)) ;
    xnor2 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix321 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_AddPToBoothOperand), .A0 (nx8289), .A1 (
          nx6437)) ;
    oai32 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix393 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .A0 (
          nx8617), .A1 (RST), .A2 (nx8299), .B0 (nx6507), .B1 (nx6575)) ;
    oai32 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix403 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .A0 (
          nx8617), .A1 (RST), .A2 (nx8299), .B0 (nx6511), .B1 (nx6575)) ;
    oai32 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix413 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .A0 (
          nx8617), .A1 (RST), .A2 (nx8299), .B0 (nx6515), .B1 (nx6575)) ;
    oai32 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix423 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .A0 (
          nx8617), .A1 (RST), .A2 (nx8299), .B0 (nx6519), .B1 (nx6575)) ;
    oai32 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix433 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .A0 (
          nx8617), .A1 (RST), .A2 (nx8299), .B0 (nx6523), .B1 (nx6575)) ;
    oai32 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix443 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .A0 (
          nx8617), .A1 (RST), .A2 (nx8299), .B0 (nx6527), .B1 (nx6575)) ;
    oai32 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix453 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .A0 (
          nx8617), .A1 (RST), .A2 (nx8301), .B0 (nx6531), .B1 (nx6575)) ;
    oai32 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix463 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .A0 (
          nx8619), .A1 (RST), .A2 (nx8301), .B0 (nx6535), .B1 (nx6577)) ;
    oai32 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix473 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .A0 (
          nx8619), .A1 (RST), .A2 (nx8301), .B0 (nx6539), .B1 (nx6577)) ;
    oai32 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix483 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .A0 (
          nx6579), .A1 (RST), .A2 (nx8301), .B0 (nx6543), .B1 (nx6577)) ;
    inv01 ix6578 (.Y (nx6579), .A (CacheFilter_4__3__0)) ;
    oai32 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix493 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .A0 (
          nx6581), .A1 (RST), .A2 (nx8301), .B0 (nx6547), .B1 (nx6577)) ;
    inv01 ix6580 (.Y (nx6581), .A (CacheFilter_4__3__1)) ;
    oai32 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix503 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .A0 (
          nx6583), .A1 (RST), .A2 (nx8301), .B0 (nx6551), .B1 (nx6577)) ;
    inv01 ix6582 (.Y (nx6583), .A (CacheFilter_4__3__2)) ;
    oai32 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix513 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .A0 (
          nx6585), .A1 (RST), .A2 (nx8301), .B0 (nx6555), .B1 (nx6577)) ;
    inv01 ix6584 (.Y (nx6585), .A (CacheFilter_4__3__3)) ;
    oai32 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix523 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .A0 (
          nx6587), .A1 (RST), .A2 (nx8303), .B0 (nx6559), .B1 (nx6577)) ;
    inv01 ix6586 (.Y (nx6587), .A (CacheFilter_4__3__4)) ;
    oai32 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix533 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .A0 (
          nx6589), .A1 (RST), .A2 (nx8303), .B0 (nx6563), .B1 (nx6591)) ;
    inv01 ix6588 (.Y (nx6589), .A (CacheFilter_4__3__5)) ;
    inv01 ix6590 (.Y (nx6591), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566)) ;
    oai32 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix543 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .A0 (
          nx6593), .A1 (RST), .A2 (nx8303), .B0 (nx6567), .B1 (nx6591)) ;
    inv01 ix6592 (.Y (nx6593), .A (CacheFilter_4__3__6)) ;
    oai32 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix553 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .A0 (
          nx6595), .A1 (RST), .A2 (nx8303), .B0 (nx6571), .B1 (nx6591)) ;
    inv01 ix6594 (.Y (nx6595), .A (CacheFilter_4__3__7)) ;
    nand02_2x CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix633 (.Y (
              nx6575), .A0 (nx7375), .A1 (nx8303)) ;
    nand02_2x CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix635 (.Y (
              nx6577), .A0 (nx7377), .A1 (nx8303)) ;
    oai32 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix393 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .A0 (
          nx8619), .A1 (RST), .A2 (nx8305), .B0 (nx6505), .B1 (nx6597)) ;
    oai32 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix403 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .A0 (
          nx8619), .A1 (RST), .A2 (nx8305), .B0 (nx6509), .B1 (nx6597)) ;
    oai32 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix413 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .A0 (
          nx8619), .A1 (RST), .A2 (nx8305), .B0 (nx6513), .B1 (nx6597)) ;
    oai32 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix423 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .A0 (
          nx8619), .A1 (RST), .A2 (nx8305), .B0 (nx6517), .B1 (nx6597)) ;
    oai32 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix433 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .A0 (
          nx8619), .A1 (RST), .A2 (nx8305), .B0 (nx6521), .B1 (nx6597)) ;
    oai32 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix443 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .A0 (
          nx8621), .A1 (RST), .A2 (nx8305), .B0 (nx6525), .B1 (nx6597)) ;
    oai32 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix453 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .A0 (
          nx8621), .A1 (RST), .A2 (nx8307), .B0 (nx6529), .B1 (nx6597)) ;
    oai32 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix463 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .A0 (
          nx8621), .A1 (RST), .A2 (nx8307), .B0 (nx6533), .B1 (nx6599)) ;
    oai32 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix473 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .A0 (
          nx8621), .A1 (RST), .A2 (nx8307), .B0 (nx6537), .B1 (nx6599)) ;
    oai32 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix483 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .A0 (
          nx6579), .A1 (RST), .A2 (nx8307), .B0 (nx6541), .B1 (nx6599)) ;
    oai32 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix493 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .A0 (
          nx6601), .A1 (RST), .A2 (nx8307), .B0 (nx6545), .B1 (nx6599)) ;
    inv01 ix6600 (.Y (nx6601), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_10)) ;
    oai32 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix503 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .A0 (
          nx6603), .A1 (RST), .A2 (nx8307), .B0 (nx6549), .B1 (nx6599)) ;
    inv01 ix6602 (.Y (nx6603), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_11)) ;
    oai32 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix513 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .A0 (
          nx6605), .A1 (RST), .A2 (nx8307), .B0 (nx6553), .B1 (nx6599)) ;
    inv01 ix6604 (.Y (nx6605), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_12)) ;
    oai32 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix523 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .A0 (
          nx6607), .A1 (RST), .A2 (nx8309), .B0 (nx6557), .B1 (nx6599)) ;
    inv01 ix6606 (.Y (nx6607), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_13)) ;
    oai32 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix533 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .A0 (
          nx6609), .A1 (RST), .A2 (nx8309), .B0 (nx6561), .B1 (nx6611)) ;
    inv01 ix6608 (.Y (nx6609), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_14)) ;
    inv01 ix6610 (.Y (nx6611), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566)) ;
    oai32 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix543 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .A0 (
          nx6613), .A1 (RST), .A2 (nx8309), .B0 (nx6565), .B1 (nx6611)) ;
    inv01 ix6612 (.Y (nx6613), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_15)) ;
    oai32 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix553 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .A0 (
          nx6615), .A1 (RST), .A2 (nx8309), .B0 (nx6569), .B1 (nx6611)) ;
    inv01 ix6614 (.Y (nx6615), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_16)) ;
    nand02_2x CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix633 (.Y (
              nx6597), .A0 (nx7377), .A1 (nx8309)) ;
    nand02_2x CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix635 (.Y (
              nx6599), .A0 (nx7377), .A1 (nx8309)) ;
    oai32 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix393 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .A0 (
          nx6617), .A1 (RST), .A2 (nx8311), .B0 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_nx384), .B1 (nx6619)) ;
    inv01 ix6616 (.Y (nx6617), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_0)) ;
    oai32 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix403 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .A0 (
          nx6621), .A1 (RST), .A2 (nx8311), .B0 (nx6437), .B1 (nx6619)) ;
    inv01 ix6620 (.Y (nx6621), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_1)) ;
    oai32 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix413 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .A0 (
          nx6623), .A1 (RST), .A2 (nx8311), .B0 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx387), .B1 (nx6619)) ;
    inv01 ix6622 (.Y (nx6623), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_2)) ;
    oai32 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix423 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .A0 (
          nx6625), .A1 (RST), .A2 (nx8311), .B0 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx399), .B1 (nx6619)) ;
    inv01 ix6624 (.Y (nx6625), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_3)) ;
    oai32 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix433 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .A0 (
          nx6627), .A1 (RST), .A2 (nx8311), .B0 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx409), .B1 (nx6619)) ;
    inv01 ix6626 (.Y (nx6627), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_4)) ;
    oai32 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix443 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .A0 (
          nx6629), .A1 (RST), .A2 (nx8311), .B0 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx419), .B1 (nx6619)) ;
    inv01 ix6628 (.Y (nx6629), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_5)) ;
    oai32 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix453 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .A0 (
          nx6631), .A1 (RST), .A2 (nx8311), .B0 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx429), .B1 (nx6619)) ;
    inv01 ix6630 (.Y (nx6631), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_6)) ;
    oai32 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix463 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .A0 (
          nx6633), .A1 (RST), .A2 (nx8313), .B0 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx439), .B1 (nx6635)) ;
    inv01 ix6632 (.Y (nx6633), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_7)) ;
    oai32 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix473 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .A0 (
          nx6637), .A1 (RST), .A2 (nx8313), .B0 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx449), .B1 (nx6635)) ;
    inv01 ix6636 (.Y (nx6637), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_8)) ;
    oai32 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix483 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .A0 (
          nx6639), .A1 (RST), .A2 (nx8313), .B0 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx469), .B1 (nx6635)) ;
    inv01 ix6638 (.Y (nx6639), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_9)) ;
    oai32 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix493 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .A0 (
          nx6641), .A1 (RST), .A2 (nx8313), .B0 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx477), .B1 (nx6635)) ;
    inv01 ix6640 (.Y (nx6641), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_10)) ;
    oai32 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix503 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .A0 (
          nx6643), .A1 (RST), .A2 (nx8313), .B0 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx485), .B1 (nx6635)) ;
    inv01 ix6642 (.Y (nx6643), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_11)) ;
    oai32 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix513 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .A0 (
          nx6645), .A1 (RST), .A2 (nx8313), .B0 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx493), .B1 (nx6635)) ;
    inv01 ix6644 (.Y (nx6645), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_12)) ;
    oai32 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix523 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .A0 (
          nx6647), .A1 (RST), .A2 (nx8313), .B0 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx501), .B1 (nx6635)) ;
    inv01 ix6646 (.Y (nx6647), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_13)) ;
    oai32 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix533 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .A0 (
          nx6649), .A1 (RST), .A2 (nx8315), .B0 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx509), .B1 (nx6651)) ;
    inv01 ix6648 (.Y (nx6649), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_14)) ;
    inv01 ix6650 (.Y (nx6651), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566)) ;
    oai32 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix543 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .A0 (
          nx6653), .A1 (RST), .A2 (nx8315), .B0 (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_nx517), .B1 (nx6651)) ;
    inv01 ix6652 (.Y (nx6653), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_15)) ;
    oai32 CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix553 (.Y (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .A0 (
          nx6655), .A1 (RST), .A2 (nx8315), .B0 (nx6453), .B1 (nx6651)) ;
    inv01 ix6654 (.Y (nx6655), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_16)) ;
    nand02_2x CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix633 (.Y (
              nx6619), .A0 (nx7377), .A1 (nx8315)) ;
    nand02_2x CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix635 (.Y (
              nx6635), .A0 (nx7377), .A1 (nx8315)) ;
    mux21 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix404 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx403), .A0 (nx6657), .A1 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_2), .S0 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx395)) ;
    inv01 ix6656 (.Y (nx6657), .A (CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx391)) ;
    mux21 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix414 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx413), .A0 (nx6659), .A1 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_3), .S0 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx405)) ;
    inv01 ix6658 (.Y (nx6659), .A (CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx403)) ;
    mux21 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix424 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx423), .A0 (nx6661), .A1 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_4), .S0 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx415)) ;
    inv01 ix6660 (.Y (nx6661), .A (CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx413)) ;
    mux21 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix434 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx433), .A0 (nx6663), .A1 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_5), .S0 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx425)) ;
    inv01 ix6662 (.Y (nx6663), .A (CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx423)) ;
    mux21 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix444 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx443), .A0 (nx6665), .A1 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_6), .S0 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx435)) ;
    inv01 ix6664 (.Y (nx6665), .A (CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx433)) ;
    mux21 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix454 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx453), .A0 (nx6667), .A1 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_7), .S0 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx445)) ;
    inv01 ix6666 (.Y (nx6667), .A (CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx443)) ;
    mux21 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix462 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx461), .A0 (nx6669), .A1 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_8), .S0 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx455)) ;
    inv01 ix6668 (.Y (nx6669), .A (CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx453)) ;
    mux21 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix468 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx467), .A0 (nx6671), .A1 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_9), .S0 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx463)) ;
    inv01 ix6670 (.Y (nx6671), .A (CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx461)) ;
    mux21 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix476 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx475), .A0 (nx6673), .A1 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_10), .S0 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx471)) ;
    inv01 ix6672 (.Y (nx6673), .A (CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx467)) ;
    mux21 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix484 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx483), .A0 (nx6675), .A1 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_11), .S0 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx479)) ;
    inv01 ix6674 (.Y (nx6675), .A (CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx475)) ;
    mux21 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix492 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx491), .A0 (nx6677), .A1 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_12), .S0 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx487)) ;
    inv01 ix6676 (.Y (nx6677), .A (CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx483)) ;
    mux21 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix500 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx499), .A0 (nx6679), .A1 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_13), .S0 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx495)) ;
    inv01 ix6678 (.Y (nx6679), .A (CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx491)) ;
    mux21 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix508 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx507), .A0 (nx6681), .A1 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_14), .S0 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx503)) ;
    inv01 ix6680 (.Y (nx6681), .A (CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx499)) ;
    mux21 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix516 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx515), .A0 (nx6683), .A1 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_15), .S0 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx511)) ;
    inv01 ix6682 (.Y (nx6683), .A (CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx507)) ;
    mux21 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix161 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_1), .A0 (nx6685), .A1 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx379), .S0 (nx8319)) ;
    inv01 ix6684 (.Y (nx6685), .A (CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_1)) ;
    mux21 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix181 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_2), .A0 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx387), .A1 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx389), .S0 (nx8319)) ;
    mux21 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix201 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_3), .A0 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx399), .A1 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx401), .S0 (nx8319)) ;
    mux21 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix221 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_4), .A0 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx409), .A1 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx411), .S0 (nx8319)) ;
    mux21 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix241 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_5), .A0 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx419), .A1 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx421), .S0 (nx8319)) ;
    mux21 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix261 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_6), .A0 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx429), .A1 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx431), .S0 (nx8319)) ;
    mux21 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix281 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_7), .A0 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx439), .A1 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx441), .S0 (nx8319)) ;
    mux21 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix301 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_8), .A0 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx449), .A1 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx451), .S0 (nx8321)) ;
    mux21 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix321 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_9), .A0 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx469), .A1 (nx6687), .S0 (nx8321)) ;
    inv01 ix6686 (.Y (nx6687), .A (CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx316)) ;
    mux21 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix341 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_10), .A0 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx477), .A1 (nx6689), .S0 (nx8321)) ;
    inv01 ix6688 (.Y (nx6689), .A (CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx336)) ;
    mux21 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix361 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_11), .A0 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx485), .A1 (nx6691), .S0 (nx8321)) ;
    inv01 ix6690 (.Y (nx6691), .A (CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx356)) ;
    mux21 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix381 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_12), .A0 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx493), .A1 (nx6693), .S0 (nx8321)) ;
    inv01 ix6692 (.Y (nx6693), .A (CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx376)) ;
    mux21 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix401 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_13), .A0 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx501), .A1 (nx6695), .S0 (nx8321)) ;
    inv01 ix6694 (.Y (nx6695), .A (CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx396)) ;
    mux21 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix421 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_14), .A0 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx509), .A1 (nx6697), .S0 (nx8321)) ;
    inv01 ix6696 (.Y (nx6697), .A (CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx416)) ;
    mux21 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix441 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_15), .A0 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx517), .A1 (nx6699), .S0 (nx8323)) ;
    inv01 ix6698 (.Y (nx6699), .A (CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx436)) ;
    mux21 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_ix461 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_16), .A0 (nx6701), 
          .A1 (nx6703), .S0 (nx8323)) ;
    inv01 ix6700 (.Y (nx6701), .A (CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothP_16)
          ) ;
    inv01 ix6702 (.Y (nx6703), .A (CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx456)) ;
    nor02_2x CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix81 (.Y (
             CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_nx80), .A0 (Instr), .A1 (
             nx7301)) ;
    nor02_2x CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix319 (.Y (
             CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642), .A0 (
             CALCULATOR_Start_dup_1352), .A1 (
             CALCULATOR_CalculatingBooth_dup_1315)) ;
    nor02_2x CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix85 (.Y (
             CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_0), .A0 (
             nx8333), .A1 (nx6705)) ;
    inv01 ix6704 (.Y (nx6705), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_1)) ;
    mux21 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix125 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_1), .A0 (
          nx6707), .A1 (nx6709), .S0 (nx8333)) ;
    inv01 ix6706 (.Y (nx6707), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_2)) ;
    inv01 ix6708 (.Y (nx6709), .A (CacheWindow_4__4__0)) ;
    mux21 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix133 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_2), .A0 (
          nx6711), .A1 (nx6713), .S0 (nx8333)) ;
    inv01 ix6710 (.Y (nx6711), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_3)) ;
    inv01 ix6712 (.Y (nx6713), .A (CacheWindow_4__4__1)) ;
    mux21 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix141 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_3), .A0 (
          nx6715), .A1 (nx6717), .S0 (nx8333)) ;
    inv01 ix6714 (.Y (nx6715), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_4)) ;
    inv01 ix6716 (.Y (nx6717), .A (CacheWindow_4__4__2)) ;
    mux21 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix149 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_4), .A0 (
          nx6719), .A1 (nx6721), .S0 (nx8333)) ;
    inv01 ix6718 (.Y (nx6719), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_5)) ;
    inv01 ix6720 (.Y (nx6721), .A (CacheWindow_4__4__3)) ;
    mux21 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix157 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_5), .A0 (
          nx6723), .A1 (nx6725), .S0 (nx8333)) ;
    inv01 ix6722 (.Y (nx6723), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_6)) ;
    inv01 ix6724 (.Y (nx6725), .A (CacheWindow_4__4__4)) ;
    mux21 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix165 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_6), .A0 (
          nx6727), .A1 (nx6729), .S0 (nx8333)) ;
    inv01 ix6726 (.Y (nx6727), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_7)) ;
    inv01 ix6728 (.Y (nx6729), .A (CacheWindow_4__4__5)) ;
    mux21 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix173 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_7), .A0 (
          nx6731), .A1 (nx6733), .S0 (nx8335)) ;
    inv01 ix6730 (.Y (nx6731), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_8)) ;
    inv01 ix6732 (.Y (nx6733), .A (CacheWindow_4__4__6)) ;
    mux21 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix181 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_8), .A0 (
          nx6735), .A1 (nx6737), .S0 (nx8335)) ;
    inv01 ix6734 (.Y (nx6735), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_9)) ;
    inv01 ix6736 (.Y (nx6737), .A (CacheWindow_4__4__7)) ;
    nor02_2x CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix89 (.Y (
             CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_9), .A0 (
             nx8335), .A1 (nx6739)) ;
    inv01 ix6738 (.Y (nx6739), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_10)) ;
    nor02_2x CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix93 (.Y (
             CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_10), .A0 (
             nx8335), .A1 (nx6741)) ;
    inv01 ix6740 (.Y (nx6741), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_11)) ;
    nor02_2x CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix97 (.Y (
             CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_11), .A0 (
             nx8335), .A1 (nx6743)) ;
    inv01 ix6742 (.Y (nx6743), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_12)) ;
    nor02_2x CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix101 (.Y (
             CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_12), .A0 (
             nx8335), .A1 (nx6745)) ;
    inv01 ix6744 (.Y (nx6745), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_13)) ;
    nor02_2x CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix105 (.Y (
             CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_13), .A0 (
             nx8335), .A1 (nx6747)) ;
    inv01 ix6746 (.Y (nx6747), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_14)) ;
    nor02_2x CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix109 (.Y (
             CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_14), .A0 (
             nx8337), .A1 (nx6749)) ;
    inv01 ix6748 (.Y (nx6749), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_15)) ;
    nor02_2x CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix113 (.Y (
             CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_15), .A0 (
             nx8337), .A1 (nx6751)) ;
    inv01 ix6750 (.Y (nx6751), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_16)) ;
    nor02_2x CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix117 (.Y (
             CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_16), .A0 (
             nx8337), .A1 (nx6751)) ;
    mux21 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix189 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothOperand_0), .A0 (nx6753), .A1 (
          nx6755), .S0 (nx8325)) ;
    inv01 ix6752 (.Y (nx6753), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_0)) ;
    inv01 ix6754 (.Y (nx6755), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_0)) ;
    mux21 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix197 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothOperand_1), .A0 (nx6757), .A1 (
          nx6759), .S0 (nx8325)) ;
    inv01 ix6756 (.Y (nx6757), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_1)) ;
    inv01 ix6758 (.Y (nx6759), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_1)) ;
    mux21 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix205 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothOperand_2), .A0 (nx6761), .A1 (
          nx6763), .S0 (nx8325)) ;
    inv01 ix6760 (.Y (nx6761), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_2)) ;
    inv01 ix6762 (.Y (nx6763), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_2)) ;
    mux21 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix213 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothOperand_3), .A0 (nx6765), .A1 (
          nx6767), .S0 (nx8325)) ;
    inv01 ix6764 (.Y (nx6765), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_3)) ;
    inv01 ix6766 (.Y (nx6767), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_3)) ;
    mux21 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix221 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothOperand_4), .A0 (nx6769), .A1 (
          nx6771), .S0 (nx8325)) ;
    inv01 ix6768 (.Y (nx6769), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_4)) ;
    inv01 ix6770 (.Y (nx6771), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_4)) ;
    mux21 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix229 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothOperand_5), .A0 (nx6773), .A1 (
          nx6775), .S0 (nx8327)) ;
    inv01 ix6772 (.Y (nx6773), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_5)) ;
    inv01 ix6774 (.Y (nx6775), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_5)) ;
    mux21 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix237 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothOperand_6), .A0 (nx6777), .A1 (
          nx6779), .S0 (nx8327)) ;
    inv01 ix6776 (.Y (nx6777), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_6)) ;
    inv01 ix6778 (.Y (nx6779), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_6)) ;
    mux21 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix245 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothOperand_7), .A0 (nx6781), .A1 (
          nx6783), .S0 (nx8327)) ;
    inv01 ix6780 (.Y (nx6781), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_7)) ;
    inv01 ix6782 (.Y (nx6783), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_7)) ;
    mux21 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix253 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothOperand_8), .A0 (nx6785), .A1 (
          nx6787), .S0 (nx8327)) ;
    inv01 ix6784 (.Y (nx6785), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_8)) ;
    inv01 ix6786 (.Y (nx6787), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_8)) ;
    mux21 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix261 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothOperand_9), .A0 (nx6789), .A1 (
          nx6791), .S0 (nx8327)) ;
    inv01 ix6788 (.Y (nx6789), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_9)) ;
    inv01 ix6790 (.Y (nx6791), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_9)) ;
    mux21 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix269 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothOperand_10), .A0 (nx6793), .A1 (
          nx6795), .S0 (nx8327)) ;
    inv01 ix6792 (.Y (nx6793), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_10)) ;
    inv01 ix6794 (.Y (nx6795), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_10)) ;
    mux21 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix277 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothOperand_11), .A0 (nx6797), .A1 (
          nx6799), .S0 (nx8327)) ;
    inv01 ix6796 (.Y (nx6797), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_11)) ;
    inv01 ix6798 (.Y (nx6799), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_11)) ;
    mux21 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix285 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothOperand_12), .A0 (nx6801), .A1 (
          nx6803), .S0 (nx8329)) ;
    inv01 ix6800 (.Y (nx6801), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_12)) ;
    inv01 ix6802 (.Y (nx6803), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_12)) ;
    mux21 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix293 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothOperand_13), .A0 (nx6805), .A1 (
          nx6807), .S0 (nx8329)) ;
    inv01 ix6804 (.Y (nx6805), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_13)) ;
    inv01 ix6806 (.Y (nx6807), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_13)) ;
    mux21 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix301 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothOperand_14), .A0 (nx6809), .A1 (
          nx6811), .S0 (nx8329)) ;
    inv01 ix6808 (.Y (nx6809), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_14)) ;
    inv01 ix6810 (.Y (nx6811), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_14)) ;
    mux21 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix309 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothOperand_15), .A0 (nx6813), .A1 (
          nx6815), .S0 (nx8329)) ;
    inv01 ix6812 (.Y (nx6813), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_15)) ;
    inv01 ix6814 (.Y (nx6815), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_15)) ;
    mux21 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix317 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BoothOperand_16), .A0 (nx6817), .A1 (
          nx6819), .S0 (nx8329)) ;
    inv01 ix6816 (.Y (nx6817), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_16)) ;
    inv01 ix6818 (.Y (nx6819), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_16)) ;
    xnor2 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix321 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_AddPToBoothOperand), .A0 (nx8329), .A1 (
          nx6685)) ;
    oai32 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix393 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .A0 (
          nx8623), .A1 (RST), .A2 (nx8339), .B0 (nx6755), .B1 (nx6823)) ;
    oai32 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix403 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .A0 (
          nx8623), .A1 (RST), .A2 (nx8339), .B0 (nx6759), .B1 (nx6823)) ;
    oai32 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix413 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .A0 (
          nx8623), .A1 (RST), .A2 (nx8339), .B0 (nx6763), .B1 (nx6823)) ;
    oai32 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix423 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .A0 (
          nx8623), .A1 (RST), .A2 (nx8339), .B0 (nx6767), .B1 (nx6823)) ;
    oai32 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix433 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .A0 (
          nx8623), .A1 (RST), .A2 (nx8339), .B0 (nx6771), .B1 (nx6823)) ;
    oai32 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix443 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .A0 (
          nx8623), .A1 (RST), .A2 (nx8339), .B0 (nx6775), .B1 (nx6823)) ;
    oai32 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix453 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .A0 (
          nx8623), .A1 (RST), .A2 (nx8341), .B0 (nx6779), .B1 (nx6823)) ;
    oai32 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix463 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .A0 (
          nx8625), .A1 (RST), .A2 (nx8341), .B0 (nx6783), .B1 (nx6825)) ;
    oai32 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix473 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .A0 (
          nx8625), .A1 (RST), .A2 (nx8341), .B0 (nx6787), .B1 (nx6825)) ;
    oai32 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix483 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .A0 (
          nx6827), .A1 (RST), .A2 (nx8341), .B0 (nx6791), .B1 (nx6825)) ;
    inv01 ix6826 (.Y (nx6827), .A (CacheFilter_4__4__0)) ;
    oai32 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix493 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .A0 (
          nx6829), .A1 (RST), .A2 (nx8341), .B0 (nx6795), .B1 (nx6825)) ;
    inv01 ix6828 (.Y (nx6829), .A (CacheFilter_4__4__1)) ;
    oai32 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix503 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .A0 (
          nx6831), .A1 (RST), .A2 (nx8341), .B0 (nx6799), .B1 (nx6825)) ;
    inv01 ix6830 (.Y (nx6831), .A (CacheFilter_4__4__2)) ;
    oai32 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix513 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .A0 (
          nx6833), .A1 (RST), .A2 (nx8341), .B0 (nx6803), .B1 (nx6825)) ;
    inv01 ix6832 (.Y (nx6833), .A (CacheFilter_4__4__3)) ;
    oai32 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix523 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .A0 (
          nx6835), .A1 (RST), .A2 (nx8343), .B0 (nx6807), .B1 (nx6825)) ;
    inv01 ix6834 (.Y (nx6835), .A (CacheFilter_4__4__4)) ;
    oai32 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix533 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .A0 (
          nx6837), .A1 (RST), .A2 (nx8343), .B0 (nx6811), .B1 (nx6839)) ;
    inv01 ix6836 (.Y (nx6837), .A (CacheFilter_4__4__5)) ;
    inv01 ix6838 (.Y (nx6839), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566)) ;
    oai32 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix543 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .A0 (
          nx6841), .A1 (RST), .A2 (nx8343), .B0 (nx6815), .B1 (nx6839)) ;
    inv01 ix6840 (.Y (nx6841), .A (CacheFilter_4__4__6)) ;
    oai32 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix553 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .A0 (
          nx6843), .A1 (RST), .A2 (nx8343), .B0 (nx6819), .B1 (nx6839)) ;
    inv01 ix6842 (.Y (nx6843), .A (CacheFilter_4__4__7)) ;
    nand02_2x CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix633 (.Y (
              nx6823), .A0 (nx7377), .A1 (nx8343)) ;
    nand02_2x CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix635 (.Y (
              nx6825), .A0 (nx7377), .A1 (nx8343)) ;
    oai32 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix393 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .A0 (
          nx8625), .A1 (RST), .A2 (nx8345), .B0 (nx6753), .B1 (nx6845)) ;
    oai32 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix403 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .A0 (
          nx8625), .A1 (RST), .A2 (nx8345), .B0 (nx6757), .B1 (nx6845)) ;
    oai32 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix413 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .A0 (
          nx8625), .A1 (RST), .A2 (nx8345), .B0 (nx6761), .B1 (nx6845)) ;
    oai32 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix423 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .A0 (
          nx8625), .A1 (RST), .A2 (nx8345), .B0 (nx6765), .B1 (nx6845)) ;
    oai32 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix433 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .A0 (
          nx8625), .A1 (RST), .A2 (nx8345), .B0 (nx6769), .B1 (nx6845)) ;
    oai32 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix443 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .A0 (
          nx8627), .A1 (RST), .A2 (nx8345), .B0 (nx6773), .B1 (nx6845)) ;
    oai32 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix453 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .A0 (
          nx8627), .A1 (RST), .A2 (nx8347), .B0 (nx6777), .B1 (nx6845)) ;
    oai32 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix463 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .A0 (
          nx8627), .A1 (RST), .A2 (nx8347), .B0 (nx6781), .B1 (nx6847)) ;
    oai32 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix473 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .A0 (
          nx8627), .A1 (RST), .A2 (nx8347), .B0 (nx6785), .B1 (nx6847)) ;
    oai32 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix483 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .A0 (
          nx6827), .A1 (RST), .A2 (nx8347), .B0 (nx6789), .B1 (nx6847)) ;
    oai32 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix493 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .A0 (
          nx6849), .A1 (RST), .A2 (nx8347), .B0 (nx6793), .B1 (nx6847)) ;
    inv01 ix6848 (.Y (nx6849), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_10)) ;
    oai32 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix503 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .A0 (
          nx6851), .A1 (RST), .A2 (nx8347), .B0 (nx6797), .B1 (nx6847)) ;
    inv01 ix6850 (.Y (nx6851), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_11)) ;
    oai32 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix513 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .A0 (
          nx6853), .A1 (RST), .A2 (nx8347), .B0 (nx6801), .B1 (nx6847)) ;
    inv01 ix6852 (.Y (nx6853), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_12)) ;
    oai32 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix523 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .A0 (
          nx6855), .A1 (RST), .A2 (nx8349), .B0 (nx6805), .B1 (nx6847)) ;
    inv01 ix6854 (.Y (nx6855), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_13)) ;
    oai32 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix533 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .A0 (
          nx6857), .A1 (RST), .A2 (nx8349), .B0 (nx6809), .B1 (nx6859)) ;
    inv01 ix6856 (.Y (nx6857), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_14)) ;
    inv01 ix6858 (.Y (nx6859), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566)) ;
    oai32 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix543 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .A0 (
          nx6861), .A1 (RST), .A2 (nx8349), .B0 (nx6813), .B1 (nx6859)) ;
    inv01 ix6860 (.Y (nx6861), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_15)) ;
    oai32 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix553 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .A0 (
          nx6863), .A1 (RST), .A2 (nx8349), .B0 (nx6817), .B1 (nx6859)) ;
    inv01 ix6862 (.Y (nx6863), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_16)) ;
    nand02_2x CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix633 (.Y (
              nx6845), .A0 (
              CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx564), .A1 (
              nx8349)) ;
    nand02_2x CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix635 (.Y (
              nx6847), .A0 (
              CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx564), .A1 (
              nx8349)) ;
    oai32 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix393 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .A0 (
          nx6865), .A1 (RST), .A2 (nx8351), .B0 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_nx384), .B1 (nx6867)) ;
    inv01 ix6864 (.Y (nx6865), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_0)) ;
    oai32 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix403 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .A0 (
          nx6869), .A1 (RST), .A2 (nx8351), .B0 (nx6685), .B1 (nx6867)) ;
    inv01 ix6868 (.Y (nx6869), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_1)) ;
    oai32 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix413 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .A0 (
          nx6871), .A1 (RST), .A2 (nx8351), .B0 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx387), .B1 (nx6867)) ;
    inv01 ix6870 (.Y (nx6871), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_2)) ;
    oai32 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix423 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .A0 (
          nx6873), .A1 (RST), .A2 (nx8351), .B0 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx399), .B1 (nx6867)) ;
    inv01 ix6872 (.Y (nx6873), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_3)) ;
    oai32 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix433 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .A0 (
          nx6875), .A1 (RST), .A2 (nx8351), .B0 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx409), .B1 (nx6867)) ;
    inv01 ix6874 (.Y (nx6875), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_4)) ;
    oai32 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix443 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .A0 (
          nx6877), .A1 (RST), .A2 (nx8351), .B0 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx419), .B1 (nx6867)) ;
    inv01 ix6876 (.Y (nx6877), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_5)) ;
    oai32 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix453 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .A0 (
          nx6879), .A1 (RST), .A2 (nx8351), .B0 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx429), .B1 (nx6867)) ;
    inv01 ix6878 (.Y (nx6879), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_6)) ;
    oai32 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix463 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .A0 (
          nx6881), .A1 (RST), .A2 (nx8353), .B0 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx439), .B1 (nx6883)) ;
    inv01 ix6880 (.Y (nx6881), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_7)) ;
    oai32 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix473 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .A0 (
          nx6885), .A1 (RST), .A2 (nx8353), .B0 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx449), .B1 (nx6883)) ;
    inv01 ix6884 (.Y (nx6885), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_8)) ;
    oai32 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix483 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .A0 (
          nx6887), .A1 (RST), .A2 (nx8353), .B0 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx469), .B1 (nx6883)) ;
    inv01 ix6886 (.Y (nx6887), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_9)) ;
    oai32 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix493 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .A0 (
          nx6889), .A1 (RST), .A2 (nx8353), .B0 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx477), .B1 (nx6883)) ;
    inv01 ix6888 (.Y (nx6889), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_10)) ;
    oai32 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix503 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .A0 (
          nx6891), .A1 (RST), .A2 (nx8353), .B0 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx485), .B1 (nx6883)) ;
    inv01 ix6890 (.Y (nx6891), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_11)) ;
    oai32 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix513 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .A0 (
          nx6893), .A1 (RST), .A2 (nx8353), .B0 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx493), .B1 (nx6883)) ;
    inv01 ix6892 (.Y (nx6893), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_12)) ;
    oai32 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix523 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .A0 (
          nx6895), .A1 (RST), .A2 (nx8353), .B0 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx501), .B1 (nx6883)) ;
    inv01 ix6894 (.Y (nx6895), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_13)) ;
    oai32 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix533 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .A0 (
          nx6897), .A1 (RST), .A2 (nx8355), .B0 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx509), .B1 (nx6899)) ;
    inv01 ix6896 (.Y (nx6897), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_14)) ;
    inv01 ix6898 (.Y (nx6899), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566)) ;
    oai32 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix543 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .A0 (
          nx6901), .A1 (RST), .A2 (nx8355), .B0 (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_nx517), .B1 (nx6899)) ;
    inv01 ix6900 (.Y (nx6901), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_15)) ;
    oai32 CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix553 (.Y (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .A0 (
          nx6903), .A1 (RST), .A2 (nx8355), .B0 (nx6701), .B1 (nx6899)) ;
    inv01 ix6902 (.Y (nx6903), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_16)) ;
    nand02_2x CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix633 (.Y (
              nx6867), .A0 (
              CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx564), .A1 (
              nx8355)) ;
    nand02_2x CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix635 (.Y (
              nx6883), .A0 (
              CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx564), .A1 (
              nx8355)) ;
    nand02 CACHE_ix1 (.Y (CACHE_nx955), .A0 (CACHE_EN_dup_1304), .A1 (FilterSize
           )) ;
    nand02 CACHE_ix3 (.Y (CACHE_nx941), .A0 (FilterSize), .A1 (CACHE_EN_dup_1293
           )) ;
    oai32 CACHE_L0_0_L1_0_Fij_ix213 (.Y (CACHE_L0_0_L1_0_Fij_nx212), .A0 (nx2115
          ), .A1 (nx8357), .A2 (nx6905), .B0 (nx875), .B1 (nx8629)) ;
    inv02 ix6904 (.Y (nx6905), .A (CACHE_L0_0_L1_0_Fij_nx331)) ;
    oai32 CACHE_L0_0_L1_0_Fij_ix223 (.Y (CACHE_L0_0_L1_0_Fij_nx222), .A0 (nx2117
          ), .A1 (nx8357), .A2 (nx6905), .B0 (nx877), .B1 (nx8629)) ;
    oai32 CACHE_L0_0_L1_0_Fij_ix233 (.Y (CACHE_L0_0_L1_0_Fij_nx232), .A0 (nx2119
          ), .A1 (nx8357), .A2 (nx6905), .B0 (nx879), .B1 (nx8629)) ;
    oai32 CACHE_L0_0_L1_0_Fij_ix243 (.Y (CACHE_L0_0_L1_0_Fij_nx242), .A0 (nx2121
          ), .A1 (nx8357), .A2 (nx6905), .B0 (nx881), .B1 (nx8629)) ;
    oai32 CACHE_L0_0_L1_0_Fij_ix253 (.Y (CACHE_L0_0_L1_0_Fij_nx252), .A0 (nx2123
          ), .A1 (nx8357), .A2 (nx6905), .B0 (nx883), .B1 (nx8629)) ;
    oai32 CACHE_L0_0_L1_0_Fij_ix263 (.Y (CACHE_L0_0_L1_0_Fij_nx262), .A0 (nx2125
          ), .A1 (nx8359), .A2 (nx6905), .B0 (nx885), .B1 (nx8629)) ;
    oai32 CACHE_L0_0_L1_0_Fij_ix273 (.Y (CACHE_L0_0_L1_0_Fij_nx272), .A0 (nx2129
          ), .A1 (nx8359), .A2 (nx6909), .B0 (nx889), .B1 (nx8629)) ;
    inv01 ix6908 (.Y (nx6909), .A (CACHE_L0_0_L1_0_Fij_nx333)) ;
    oai32 CACHE_L0_0_L1_0_Fij_ix283 (.Y (CACHE_L0_0_L1_0_Fij_nx282), .A0 (nx2131
          ), .A1 (nx8359), .A2 (nx6909), .B0 (nx891), .B1 (nx8631)) ;
    oai32 CACHE_L0_0_L1_0_Wij_ix213 (.Y (CACHE_L0_0_L1_0_Wij_nx212), .A0 (nx1997
          ), .A1 (nx8359), .A2 (nx6911), .B0 (nx757), .B1 (nx8633)) ;
    inv02 ix6910 (.Y (nx6911), .A (CACHE_L0_0_L1_0_Wij_nx331)) ;
    oai32 CACHE_L0_0_L1_0_Wij_ix223 (.Y (CACHE_L0_0_L1_0_Wij_nx222), .A0 (nx2001
          ), .A1 (nx8359), .A2 (nx6911), .B0 (nx761), .B1 (nx8633)) ;
    oai32 CACHE_L0_0_L1_0_Wij_ix233 (.Y (CACHE_L0_0_L1_0_Wij_nx232), .A0 (nx2005
          ), .A1 (nx8359), .A2 (nx6911), .B0 (nx765), .B1 (nx8633)) ;
    oai32 CACHE_L0_0_L1_0_Wij_ix243 (.Y (CACHE_L0_0_L1_0_Wij_nx242), .A0 (nx2009
          ), .A1 (nx8359), .A2 (nx6911), .B0 (nx769), .B1 (nx8633)) ;
    oai32 CACHE_L0_0_L1_0_Wij_ix253 (.Y (CACHE_L0_0_L1_0_Wij_nx252), .A0 (nx2013
          ), .A1 (CACHE_RST_dup_1073), .A2 (nx6911), .B0 (nx773), .B1 (nx8633)
          ) ;
    oai32 CACHE_L0_0_L1_0_Wij_ix263 (.Y (CACHE_L0_0_L1_0_Wij_nx262), .A0 (nx2017
          ), .A1 (CACHE_RST_dup_1073), .A2 (nx6911), .B0 (nx777), .B1 (nx8633)
          ) ;
    oai32 CACHE_L0_0_L1_0_Wij_ix273 (.Y (CACHE_L0_0_L1_0_Wij_nx272), .A0 (nx2021
          ), .A1 (CACHE_RST_dup_1073), .A2 (nx6915), .B0 (nx781), .B1 (nx8633)
          ) ;
    inv01 ix6914 (.Y (nx6915), .A (CACHE_L0_0_L1_0_Wij_nx333)) ;
    oai32 CACHE_L0_0_L1_0_Wij_ix283 (.Y (CACHE_L0_0_L1_0_Wij_nx282), .A0 (nx2025
          ), .A1 (CACHE_RST_dup_1073), .A2 (nx6915), .B0 (nx785), .B1 (nx8635)
          ) ;
    oai32 CACHE_L0_0_L1_1_Fij_ix213 (.Y (CACHE_L0_0_L1_1_Fij_nx212), .A0 (nx2363
          ), .A1 (nx8361), .A2 (nx6917), .B0 (nx1123), .B1 (nx8637)) ;
    inv02 ix6916 (.Y (nx6917), .A (CACHE_L0_0_L1_1_Fij_nx331)) ;
    oai32 CACHE_L0_0_L1_1_Fij_ix223 (.Y (CACHE_L0_0_L1_1_Fij_nx222), .A0 (nx2365
          ), .A1 (nx8361), .A2 (nx6917), .B0 (nx1125), .B1 (nx8637)) ;
    oai32 CACHE_L0_0_L1_1_Fij_ix233 (.Y (CACHE_L0_0_L1_1_Fij_nx232), .A0 (nx2367
          ), .A1 (nx8361), .A2 (nx6917), .B0 (nx1127), .B1 (nx8637)) ;
    oai32 CACHE_L0_0_L1_1_Fij_ix243 (.Y (CACHE_L0_0_L1_1_Fij_nx242), .A0 (nx2369
          ), .A1 (nx8361), .A2 (nx6917), .B0 (nx1129), .B1 (nx8637)) ;
    oai32 CACHE_L0_0_L1_1_Fij_ix253 (.Y (CACHE_L0_0_L1_1_Fij_nx252), .A0 (nx2371
          ), .A1 (nx8361), .A2 (nx6917), .B0 (nx1131), .B1 (nx8637)) ;
    oai32 CACHE_L0_0_L1_1_Fij_ix263 (.Y (CACHE_L0_0_L1_1_Fij_nx262), .A0 (nx2373
          ), .A1 (nx8363), .A2 (nx6917), .B0 (nx1133), .B1 (nx8637)) ;
    oai32 CACHE_L0_0_L1_1_Fij_ix273 (.Y (CACHE_L0_0_L1_1_Fij_nx272), .A0 (nx2377
          ), .A1 (nx8363), .A2 (nx6921), .B0 (nx1137), .B1 (nx8637)) ;
    inv01 ix6920 (.Y (nx6921), .A (CACHE_L0_0_L1_1_Fij_nx333)) ;
    oai32 CACHE_L0_0_L1_1_Fij_ix283 (.Y (CACHE_L0_0_L1_1_Fij_nx282), .A0 (nx2379
          ), .A1 (nx8363), .A2 (nx6921), .B0 (nx1139), .B1 (nx8639)) ;
    oai32 CACHE_L0_0_L1_1_Wij_ix213 (.Y (CACHE_L0_0_L1_1_Wij_nx212), .A0 (nx2245
          ), .A1 (nx8363), .A2 (nx6923), .B0 (nx1005), .B1 (nx8641)) ;
    inv02 ix6922 (.Y (nx6923), .A (CACHE_L0_0_L1_1_Wij_nx331)) ;
    oai32 CACHE_L0_0_L1_1_Wij_ix223 (.Y (CACHE_L0_0_L1_1_Wij_nx222), .A0 (nx2249
          ), .A1 (nx8363), .A2 (nx6923), .B0 (nx1009), .B1 (nx8641)) ;
    oai32 CACHE_L0_0_L1_1_Wij_ix233 (.Y (CACHE_L0_0_L1_1_Wij_nx232), .A0 (nx2253
          ), .A1 (nx8363), .A2 (nx6923), .B0 (nx1013), .B1 (nx8641)) ;
    oai32 CACHE_L0_0_L1_1_Wij_ix243 (.Y (CACHE_L0_0_L1_1_Wij_nx242), .A0 (nx2257
          ), .A1 (nx8363), .A2 (nx6923), .B0 (nx1017), .B1 (nx8641)) ;
    oai32 CACHE_L0_0_L1_1_Wij_ix253 (.Y (CACHE_L0_0_L1_1_Wij_nx252), .A0 (nx2261
          ), .A1 (CACHE_RST_dup_1094), .A2 (nx6923), .B0 (nx1021), .B1 (nx8641)
          ) ;
    oai32 CACHE_L0_0_L1_1_Wij_ix263 (.Y (CACHE_L0_0_L1_1_Wij_nx262), .A0 (nx2265
          ), .A1 (CACHE_RST_dup_1094), .A2 (nx6923), .B0 (nx1025), .B1 (nx8641)
          ) ;
    oai32 CACHE_L0_0_L1_1_Wij_ix273 (.Y (CACHE_L0_0_L1_1_Wij_nx272), .A0 (nx2269
          ), .A1 (CACHE_RST_dup_1094), .A2 (nx6927), .B0 (nx1029), .B1 (nx8641)
          ) ;
    inv01 ix6926 (.Y (nx6927), .A (CACHE_L0_0_L1_1_Wij_nx333)) ;
    oai32 CACHE_L0_0_L1_1_Wij_ix283 (.Y (CACHE_L0_0_L1_1_Wij_nx282), .A0 (nx2273
          ), .A1 (CACHE_RST_dup_1094), .A2 (nx6927), .B0 (nx1033), .B1 (nx8643)
          ) ;
    oai32 CACHE_L0_0_L1_2_Fij_ix213 (.Y (CACHE_L0_0_L1_2_Fij_nx212), .A0 (nx2611
          ), .A1 (nx8365), .A2 (nx6929), .B0 (nx1371), .B1 (nx8645)) ;
    inv02 ix6928 (.Y (nx6929), .A (CACHE_L0_0_L1_2_Fij_nx331)) ;
    oai32 CACHE_L0_0_L1_2_Fij_ix223 (.Y (CACHE_L0_0_L1_2_Fij_nx222), .A0 (nx2613
          ), .A1 (nx8365), .A2 (nx6929), .B0 (nx1373), .B1 (nx8645)) ;
    oai32 CACHE_L0_0_L1_2_Fij_ix233 (.Y (CACHE_L0_0_L1_2_Fij_nx232), .A0 (nx2615
          ), .A1 (nx8365), .A2 (nx6929), .B0 (nx1375), .B1 (nx8645)) ;
    oai32 CACHE_L0_0_L1_2_Fij_ix243 (.Y (CACHE_L0_0_L1_2_Fij_nx242), .A0 (nx2617
          ), .A1 (nx8365), .A2 (nx6929), .B0 (nx1377), .B1 (nx8645)) ;
    oai32 CACHE_L0_0_L1_2_Fij_ix253 (.Y (CACHE_L0_0_L1_2_Fij_nx252), .A0 (nx2619
          ), .A1 (nx8365), .A2 (nx6929), .B0 (nx1379), .B1 (nx8645)) ;
    oai32 CACHE_L0_0_L1_2_Fij_ix263 (.Y (CACHE_L0_0_L1_2_Fij_nx262), .A0 (nx2621
          ), .A1 (nx8367), .A2 (nx6929), .B0 (nx1381), .B1 (nx8645)) ;
    oai32 CACHE_L0_0_L1_2_Fij_ix273 (.Y (CACHE_L0_0_L1_2_Fij_nx272), .A0 (nx2625
          ), .A1 (nx8367), .A2 (nx6933), .B0 (nx1385), .B1 (nx8645)) ;
    inv01 ix6932 (.Y (nx6933), .A (CACHE_L0_0_L1_2_Fij_nx333)) ;
    oai32 CACHE_L0_0_L1_2_Fij_ix283 (.Y (CACHE_L0_0_L1_2_Fij_nx282), .A0 (nx2627
          ), .A1 (nx8367), .A2 (nx6933), .B0 (nx1387), .B1 (nx8647)) ;
    oai32 CACHE_L0_0_L1_2_Wij_ix213 (.Y (CACHE_L0_0_L1_2_Wij_nx212), .A0 (nx2493
          ), .A1 (nx8367), .A2 (nx6935), .B0 (nx1253), .B1 (nx8649)) ;
    inv02 ix6934 (.Y (nx6935), .A (CACHE_L0_0_L1_2_Wij_nx331)) ;
    oai32 CACHE_L0_0_L1_2_Wij_ix223 (.Y (CACHE_L0_0_L1_2_Wij_nx222), .A0 (nx2497
          ), .A1 (nx8367), .A2 (nx6935), .B0 (nx1257), .B1 (nx8649)) ;
    oai32 CACHE_L0_0_L1_2_Wij_ix233 (.Y (CACHE_L0_0_L1_2_Wij_nx232), .A0 (nx2501
          ), .A1 (nx8367), .A2 (nx6935), .B0 (nx1261), .B1 (nx8649)) ;
    oai32 CACHE_L0_0_L1_2_Wij_ix243 (.Y (CACHE_L0_0_L1_2_Wij_nx242), .A0 (nx2505
          ), .A1 (nx8367), .A2 (nx6935), .B0 (nx1265), .B1 (nx8649)) ;
    oai32 CACHE_L0_0_L1_2_Wij_ix253 (.Y (CACHE_L0_0_L1_2_Wij_nx252), .A0 (nx2509
          ), .A1 (CACHE_RST_dup_1116), .A2 (nx6935), .B0 (nx1269), .B1 (nx8649)
          ) ;
    oai32 CACHE_L0_0_L1_2_Wij_ix263 (.Y (CACHE_L0_0_L1_2_Wij_nx262), .A0 (nx2513
          ), .A1 (CACHE_RST_dup_1116), .A2 (nx6935), .B0 (nx1273), .B1 (nx8649)
          ) ;
    oai32 CACHE_L0_0_L1_2_Wij_ix273 (.Y (CACHE_L0_0_L1_2_Wij_nx272), .A0 (nx2517
          ), .A1 (CACHE_RST_dup_1116), .A2 (nx6939), .B0 (nx1277), .B1 (nx8649)
          ) ;
    inv01 ix6938 (.Y (nx6939), .A (CACHE_L0_0_L1_2_Wij_nx333)) ;
    oai32 CACHE_L0_0_L1_2_Wij_ix283 (.Y (CACHE_L0_0_L1_2_Wij_nx282), .A0 (nx2521
          ), .A1 (CACHE_RST_dup_1116), .A2 (nx6939), .B0 (nx1281), .B1 (nx8651)
          ) ;
    oai32 CACHE_L0_0_L1_3_Fij_ix213 (.Y (CACHE_L0_0_L1_3_Fij_nx212), .A0 (nx2859
          ), .A1 (nx8369), .A2 (nx6941), .B0 (nx1619), .B1 (nx8653)) ;
    inv02 ix6940 (.Y (nx6941), .A (CACHE_L0_0_L1_3_Fij_nx331)) ;
    oai32 CACHE_L0_0_L1_3_Fij_ix223 (.Y (CACHE_L0_0_L1_3_Fij_nx222), .A0 (nx2861
          ), .A1 (nx8369), .A2 (nx6941), .B0 (nx1621), .B1 (nx8653)) ;
    oai32 CACHE_L0_0_L1_3_Fij_ix233 (.Y (CACHE_L0_0_L1_3_Fij_nx232), .A0 (nx2863
          ), .A1 (nx8369), .A2 (nx6941), .B0 (nx1623), .B1 (nx8653)) ;
    oai32 CACHE_L0_0_L1_3_Fij_ix243 (.Y (CACHE_L0_0_L1_3_Fij_nx242), .A0 (nx2865
          ), .A1 (nx8369), .A2 (nx6941), .B0 (nx1625), .B1 (nx8653)) ;
    oai32 CACHE_L0_0_L1_3_Fij_ix253 (.Y (CACHE_L0_0_L1_3_Fij_nx252), .A0 (nx2867
          ), .A1 (nx8369), .A2 (nx6941), .B0 (nx1627), .B1 (nx8653)) ;
    oai32 CACHE_L0_0_L1_3_Fij_ix263 (.Y (CACHE_L0_0_L1_3_Fij_nx262), .A0 (nx2869
          ), .A1 (nx8371), .A2 (nx6941), .B0 (nx1629), .B1 (nx8653)) ;
    oai32 CACHE_L0_0_L1_3_Fij_ix273 (.Y (CACHE_L0_0_L1_3_Fij_nx272), .A0 (nx2873
          ), .A1 (nx8371), .A2 (nx6945), .B0 (nx1633), .B1 (nx8653)) ;
    inv01 ix6944 (.Y (nx6945), .A (CACHE_L0_0_L1_3_Fij_nx333)) ;
    oai32 CACHE_L0_0_L1_3_Fij_ix283 (.Y (CACHE_L0_0_L1_3_Fij_nx282), .A0 (nx2875
          ), .A1 (nx8371), .A2 (nx6945), .B0 (nx1635), .B1 (nx8655)) ;
    oai32 CACHE_L0_0_L1_3_Wij_ix213 (.Y (CACHE_L0_0_L1_3_Wij_nx212), .A0 (nx2741
          ), .A1 (nx8371), .A2 (nx6947), .B0 (nx1501), .B1 (nx8657)) ;
    inv02 ix6946 (.Y (nx6947), .A (CACHE_L0_0_L1_3_Wij_nx331)) ;
    oai32 CACHE_L0_0_L1_3_Wij_ix223 (.Y (CACHE_L0_0_L1_3_Wij_nx222), .A0 (nx2745
          ), .A1 (nx8371), .A2 (nx6947), .B0 (nx1505), .B1 (nx8657)) ;
    oai32 CACHE_L0_0_L1_3_Wij_ix233 (.Y (CACHE_L0_0_L1_3_Wij_nx232), .A0 (nx2749
          ), .A1 (nx8371), .A2 (nx6947), .B0 (nx1509), .B1 (nx8657)) ;
    oai32 CACHE_L0_0_L1_3_Wij_ix243 (.Y (CACHE_L0_0_L1_3_Wij_nx242), .A0 (nx2753
          ), .A1 (nx8371), .A2 (nx6947), .B0 (nx1513), .B1 (nx8657)) ;
    oai32 CACHE_L0_0_L1_3_Wij_ix253 (.Y (CACHE_L0_0_L1_3_Wij_nx252), .A0 (nx2757
          ), .A1 (CACHE_RST_dup_1138), .A2 (nx6947), .B0 (nx1517), .B1 (nx8657)
          ) ;
    oai32 CACHE_L0_0_L1_3_Wij_ix263 (.Y (CACHE_L0_0_L1_3_Wij_nx262), .A0 (nx2761
          ), .A1 (CACHE_RST_dup_1138), .A2 (nx6947), .B0 (nx1521), .B1 (nx8657)
          ) ;
    oai32 CACHE_L0_0_L1_3_Wij_ix273 (.Y (CACHE_L0_0_L1_3_Wij_nx272), .A0 (nx2765
          ), .A1 (CACHE_RST_dup_1138), .A2 (nx6951), .B0 (nx1525), .B1 (nx8657)
          ) ;
    inv01 ix6950 (.Y (nx6951), .A (CACHE_L0_0_L1_3_Wij_nx333)) ;
    oai32 CACHE_L0_0_L1_3_Wij_ix283 (.Y (CACHE_L0_0_L1_3_Wij_nx282), .A0 (nx2769
          ), .A1 (CACHE_RST_dup_1138), .A2 (nx6951), .B0 (nx1529), .B1 (nx8659)
          ) ;
    oai32 CACHE_L0_0_L1_4_Fij_ix213 (.Y (CACHE_L0_0_L1_4_Fij_nx212), .A0 (nx3107
          ), .A1 (nx8373), .A2 (nx6953), .B0 (nx1867), .B1 (nx8661)) ;
    inv02 ix6952 (.Y (nx6953), .A (CACHE_L0_0_L1_4_Fij_nx331)) ;
    oai32 CACHE_L0_0_L1_4_Fij_ix223 (.Y (CACHE_L0_0_L1_4_Fij_nx222), .A0 (nx3109
          ), .A1 (nx8373), .A2 (nx6953), .B0 (nx1869), .B1 (nx8661)) ;
    oai32 CACHE_L0_0_L1_4_Fij_ix233 (.Y (CACHE_L0_0_L1_4_Fij_nx232), .A0 (nx3111
          ), .A1 (nx8373), .A2 (nx6953), .B0 (nx1871), .B1 (nx8661)) ;
    oai32 CACHE_L0_0_L1_4_Fij_ix243 (.Y (CACHE_L0_0_L1_4_Fij_nx242), .A0 (nx3113
          ), .A1 (nx8373), .A2 (nx6953), .B0 (nx1873), .B1 (nx8661)) ;
    oai32 CACHE_L0_0_L1_4_Fij_ix253 (.Y (CACHE_L0_0_L1_4_Fij_nx252), .A0 (nx3115
          ), .A1 (nx8373), .A2 (nx6953), .B0 (nx1875), .B1 (nx8661)) ;
    oai32 CACHE_L0_0_L1_4_Fij_ix263 (.Y (CACHE_L0_0_L1_4_Fij_nx262), .A0 (nx3117
          ), .A1 (nx8375), .A2 (nx6953), .B0 (nx1877), .B1 (nx8661)) ;
    oai32 CACHE_L0_0_L1_4_Fij_ix273 (.Y (CACHE_L0_0_L1_4_Fij_nx272), .A0 (nx3121
          ), .A1 (nx8375), .A2 (nx6957), .B0 (nx1881), .B1 (nx8661)) ;
    inv01 ix6956 (.Y (nx6957), .A (CACHE_L0_0_L1_4_Fij_nx333)) ;
    oai32 CACHE_L0_0_L1_4_Fij_ix283 (.Y (CACHE_L0_0_L1_4_Fij_nx282), .A0 (nx3123
          ), .A1 (nx8375), .A2 (nx6957), .B0 (nx1883), .B1 (nx8663)) ;
    oai32 CACHE_L0_0_L1_4_Wij_ix213 (.Y (CACHE_L0_0_L1_4_Wij_nx212), .A0 (nx2989
          ), .A1 (nx8375), .A2 (nx6959), .B0 (nx1749), .B1 (nx8665)) ;
    inv02 ix6958 (.Y (nx6959), .A (CACHE_L0_0_L1_4_Wij_nx331)) ;
    oai32 CACHE_L0_0_L1_4_Wij_ix223 (.Y (CACHE_L0_0_L1_4_Wij_nx222), .A0 (nx2993
          ), .A1 (nx8375), .A2 (nx6959), .B0 (nx1753), .B1 (nx8665)) ;
    oai32 CACHE_L0_0_L1_4_Wij_ix233 (.Y (CACHE_L0_0_L1_4_Wij_nx232), .A0 (nx2997
          ), .A1 (nx8375), .A2 (nx6959), .B0 (nx1757), .B1 (nx8665)) ;
    oai32 CACHE_L0_0_L1_4_Wij_ix243 (.Y (CACHE_L0_0_L1_4_Wij_nx242), .A0 (nx3001
          ), .A1 (nx8375), .A2 (nx6959), .B0 (nx1761), .B1 (nx8665)) ;
    oai32 CACHE_L0_0_L1_4_Wij_ix253 (.Y (CACHE_L0_0_L1_4_Wij_nx252), .A0 (nx3005
          ), .A1 (CACHE_RST_dup_1160), .A2 (nx6959), .B0 (nx1765), .B1 (nx8665)
          ) ;
    oai32 CACHE_L0_0_L1_4_Wij_ix263 (.Y (CACHE_L0_0_L1_4_Wij_nx262), .A0 (nx3009
          ), .A1 (CACHE_RST_dup_1160), .A2 (nx6959), .B0 (nx1769), .B1 (nx8665)
          ) ;
    oai32 CACHE_L0_0_L1_4_Wij_ix273 (.Y (CACHE_L0_0_L1_4_Wij_nx272), .A0 (nx3013
          ), .A1 (CACHE_RST_dup_1160), .A2 (nx6963), .B0 (nx1773), .B1 (nx8665)
          ) ;
    inv01 ix6962 (.Y (nx6963), .A (CACHE_L0_0_L1_4_Wij_nx333)) ;
    oai32 CACHE_L0_0_L1_4_Wij_ix283 (.Y (CACHE_L0_0_L1_4_Wij_nx282), .A0 (nx3017
          ), .A1 (CACHE_RST_dup_1160), .A2 (nx6963), .B0 (nx1777), .B1 (nx8667)
          ) ;
    oai32 CACHE_L0_1_L1_0_Fij_ix213 (.Y (CACHE_L0_1_L1_0_Fij_nx212), .A0 (nx3355
          ), .A1 (nx8377), .A2 (nx6965), .B0 (nx2115), .B1 (nx8669)) ;
    inv02 ix6964 (.Y (nx6965), .A (CACHE_L0_1_L1_0_Fij_nx331)) ;
    oai32 CACHE_L0_1_L1_0_Fij_ix223 (.Y (CACHE_L0_1_L1_0_Fij_nx222), .A0 (nx3357
          ), .A1 (nx8377), .A2 (nx6965), .B0 (nx2117), .B1 (nx8669)) ;
    oai32 CACHE_L0_1_L1_0_Fij_ix233 (.Y (CACHE_L0_1_L1_0_Fij_nx232), .A0 (nx3359
          ), .A1 (nx8377), .A2 (nx6965), .B0 (nx2119), .B1 (nx8669)) ;
    oai32 CACHE_L0_1_L1_0_Fij_ix243 (.Y (CACHE_L0_1_L1_0_Fij_nx242), .A0 (nx3361
          ), .A1 (nx8377), .A2 (nx6965), .B0 (nx2121), .B1 (nx8669)) ;
    oai32 CACHE_L0_1_L1_0_Fij_ix253 (.Y (CACHE_L0_1_L1_0_Fij_nx252), .A0 (nx3363
          ), .A1 (nx8377), .A2 (nx6965), .B0 (nx2123), .B1 (nx8669)) ;
    oai32 CACHE_L0_1_L1_0_Fij_ix263 (.Y (CACHE_L0_1_L1_0_Fij_nx262), .A0 (nx3365
          ), .A1 (nx8379), .A2 (nx6965), .B0 (nx2125), .B1 (nx8669)) ;
    oai32 CACHE_L0_1_L1_0_Fij_ix273 (.Y (CACHE_L0_1_L1_0_Fij_nx272), .A0 (nx3369
          ), .A1 (nx8379), .A2 (nx6969), .B0 (nx2129), .B1 (nx8669)) ;
    inv01 ix6968 (.Y (nx6969), .A (CACHE_L0_1_L1_0_Fij_nx333)) ;
    oai32 CACHE_L0_1_L1_0_Fij_ix283 (.Y (CACHE_L0_1_L1_0_Fij_nx282), .A0 (nx3371
          ), .A1 (nx8379), .A2 (nx6969), .B0 (nx2131), .B1 (nx8671)) ;
    oai32 CACHE_L0_1_L1_0_Wij_ix213 (.Y (CACHE_L0_1_L1_0_Wij_nx212), .A0 (nx3237
          ), .A1 (nx8379), .A2 (nx6971), .B0 (nx1997), .B1 (nx8673)) ;
    inv02 ix6970 (.Y (nx6971), .A (CACHE_L0_1_L1_0_Wij_nx331)) ;
    oai32 CACHE_L0_1_L1_0_Wij_ix223 (.Y (CACHE_L0_1_L1_0_Wij_nx222), .A0 (nx3241
          ), .A1 (nx8379), .A2 (nx6971), .B0 (nx2001), .B1 (nx8673)) ;
    oai32 CACHE_L0_1_L1_0_Wij_ix233 (.Y (CACHE_L0_1_L1_0_Wij_nx232), .A0 (nx3245
          ), .A1 (nx8379), .A2 (nx6971), .B0 (nx2005), .B1 (nx8673)) ;
    oai32 CACHE_L0_1_L1_0_Wij_ix243 (.Y (CACHE_L0_1_L1_0_Wij_nx242), .A0 (nx3249
          ), .A1 (nx8379), .A2 (nx6971), .B0 (nx2009), .B1 (nx8673)) ;
    oai32 CACHE_L0_1_L1_0_Wij_ix253 (.Y (CACHE_L0_1_L1_0_Wij_nx252), .A0 (nx3253
          ), .A1 (CACHE_RST_dup_1182), .A2 (nx6971), .B0 (nx2013), .B1 (nx8673)
          ) ;
    oai32 CACHE_L0_1_L1_0_Wij_ix263 (.Y (CACHE_L0_1_L1_0_Wij_nx262), .A0 (nx3257
          ), .A1 (CACHE_RST_dup_1182), .A2 (nx6971), .B0 (nx2017), .B1 (nx8673)
          ) ;
    oai32 CACHE_L0_1_L1_0_Wij_ix273 (.Y (CACHE_L0_1_L1_0_Wij_nx272), .A0 (nx3261
          ), .A1 (CACHE_RST_dup_1182), .A2 (nx6975), .B0 (nx2021), .B1 (nx8673)
          ) ;
    inv01 ix6974 (.Y (nx6975), .A (CACHE_L0_1_L1_0_Wij_nx333)) ;
    oai32 CACHE_L0_1_L1_0_Wij_ix283 (.Y (CACHE_L0_1_L1_0_Wij_nx282), .A0 (nx3265
          ), .A1 (CACHE_RST_dup_1182), .A2 (nx6975), .B0 (nx2025), .B1 (nx8675)
          ) ;
    oai32 CACHE_L0_1_L1_1_Fij_ix213 (.Y (CACHE_L0_1_L1_1_Fij_nx212), .A0 (nx3603
          ), .A1 (nx8381), .A2 (nx6977), .B0 (nx2363), .B1 (nx8677)) ;
    inv02 ix6976 (.Y (nx6977), .A (CACHE_L0_1_L1_1_Fij_nx331)) ;
    oai32 CACHE_L0_1_L1_1_Fij_ix223 (.Y (CACHE_L0_1_L1_1_Fij_nx222), .A0 (nx3605
          ), .A1 (nx8381), .A2 (nx6977), .B0 (nx2365), .B1 (nx8677)) ;
    oai32 CACHE_L0_1_L1_1_Fij_ix233 (.Y (CACHE_L0_1_L1_1_Fij_nx232), .A0 (nx3607
          ), .A1 (nx8381), .A2 (nx6977), .B0 (nx2367), .B1 (nx8677)) ;
    oai32 CACHE_L0_1_L1_1_Fij_ix243 (.Y (CACHE_L0_1_L1_1_Fij_nx242), .A0 (nx3609
          ), .A1 (nx8381), .A2 (nx6977), .B0 (nx2369), .B1 (nx8677)) ;
    oai32 CACHE_L0_1_L1_1_Fij_ix253 (.Y (CACHE_L0_1_L1_1_Fij_nx252), .A0 (nx3611
          ), .A1 (nx8381), .A2 (nx6977), .B0 (nx2371), .B1 (nx8677)) ;
    oai32 CACHE_L0_1_L1_1_Fij_ix263 (.Y (CACHE_L0_1_L1_1_Fij_nx262), .A0 (nx3613
          ), .A1 (nx8383), .A2 (nx6977), .B0 (nx2373), .B1 (nx8677)) ;
    oai32 CACHE_L0_1_L1_1_Fij_ix273 (.Y (CACHE_L0_1_L1_1_Fij_nx272), .A0 (nx3617
          ), .A1 (nx8383), .A2 (nx6981), .B0 (nx2377), .B1 (nx8677)) ;
    inv01 ix6980 (.Y (nx6981), .A (CACHE_L0_1_L1_1_Fij_nx333)) ;
    oai32 CACHE_L0_1_L1_1_Fij_ix283 (.Y (CACHE_L0_1_L1_1_Fij_nx282), .A0 (nx3619
          ), .A1 (nx8383), .A2 (nx6981), .B0 (nx2379), .B1 (nx8679)) ;
    oai32 CACHE_L0_1_L1_1_Wij_ix213 (.Y (CACHE_L0_1_L1_1_Wij_nx212), .A0 (nx3485
          ), .A1 (nx8383), .A2 (nx6983), .B0 (nx2245), .B1 (nx8681)) ;
    inv02 ix6982 (.Y (nx6983), .A (CACHE_L0_1_L1_1_Wij_nx331)) ;
    oai32 CACHE_L0_1_L1_1_Wij_ix223 (.Y (CACHE_L0_1_L1_1_Wij_nx222), .A0 (nx3489
          ), .A1 (nx8383), .A2 (nx6983), .B0 (nx2249), .B1 (nx8681)) ;
    oai32 CACHE_L0_1_L1_1_Wij_ix233 (.Y (CACHE_L0_1_L1_1_Wij_nx232), .A0 (nx3493
          ), .A1 (nx8383), .A2 (nx6983), .B0 (nx2253), .B1 (nx8681)) ;
    oai32 CACHE_L0_1_L1_1_Wij_ix243 (.Y (CACHE_L0_1_L1_1_Wij_nx242), .A0 (nx3497
          ), .A1 (nx8383), .A2 (nx6983), .B0 (nx2257), .B1 (nx8681)) ;
    oai32 CACHE_L0_1_L1_1_Wij_ix253 (.Y (CACHE_L0_1_L1_1_Wij_nx252), .A0 (nx3501
          ), .A1 (CACHE_RST_dup_1204), .A2 (nx6983), .B0 (nx2261), .B1 (nx8681)
          ) ;
    oai32 CACHE_L0_1_L1_1_Wij_ix263 (.Y (CACHE_L0_1_L1_1_Wij_nx262), .A0 (nx3505
          ), .A1 (CACHE_RST_dup_1204), .A2 (nx6983), .B0 (nx2265), .B1 (nx8681)
          ) ;
    oai32 CACHE_L0_1_L1_1_Wij_ix273 (.Y (CACHE_L0_1_L1_1_Wij_nx272), .A0 (nx3509
          ), .A1 (CACHE_RST_dup_1204), .A2 (nx6987), .B0 (nx2269), .B1 (nx8681)
          ) ;
    inv01 ix6986 (.Y (nx6987), .A (CACHE_L0_1_L1_1_Wij_nx333)) ;
    oai32 CACHE_L0_1_L1_1_Wij_ix283 (.Y (CACHE_L0_1_L1_1_Wij_nx282), .A0 (nx3513
          ), .A1 (CACHE_RST_dup_1204), .A2 (nx6987), .B0 (nx2273), .B1 (nx8683)
          ) ;
    oai32 CACHE_L0_1_L1_2_Fij_ix213 (.Y (CACHE_L0_1_L1_2_Fij_nx212), .A0 (nx3851
          ), .A1 (nx8385), .A2 (nx6989), .B0 (nx2611), .B1 (nx8685)) ;
    inv02 ix6988 (.Y (nx6989), .A (CACHE_L0_1_L1_2_Fij_nx331)) ;
    oai32 CACHE_L0_1_L1_2_Fij_ix223 (.Y (CACHE_L0_1_L1_2_Fij_nx222), .A0 (nx3853
          ), .A1 (nx8385), .A2 (nx6989), .B0 (nx2613), .B1 (nx8685)) ;
    oai32 CACHE_L0_1_L1_2_Fij_ix233 (.Y (CACHE_L0_1_L1_2_Fij_nx232), .A0 (nx3855
          ), .A1 (nx8385), .A2 (nx6989), .B0 (nx2615), .B1 (nx8685)) ;
    oai32 CACHE_L0_1_L1_2_Fij_ix243 (.Y (CACHE_L0_1_L1_2_Fij_nx242), .A0 (nx3857
          ), .A1 (nx8385), .A2 (nx6989), .B0 (nx2617), .B1 (nx8685)) ;
    oai32 CACHE_L0_1_L1_2_Fij_ix253 (.Y (CACHE_L0_1_L1_2_Fij_nx252), .A0 (nx3859
          ), .A1 (nx8385), .A2 (nx6989), .B0 (nx2619), .B1 (nx8685)) ;
    oai32 CACHE_L0_1_L1_2_Fij_ix263 (.Y (CACHE_L0_1_L1_2_Fij_nx262), .A0 (nx3861
          ), .A1 (nx8387), .A2 (nx6989), .B0 (nx2621), .B1 (nx8685)) ;
    oai32 CACHE_L0_1_L1_2_Fij_ix273 (.Y (CACHE_L0_1_L1_2_Fij_nx272), .A0 (nx3865
          ), .A1 (nx8387), .A2 (nx6993), .B0 (nx2625), .B1 (nx8685)) ;
    inv01 ix6992 (.Y (nx6993), .A (CACHE_L0_1_L1_2_Fij_nx333)) ;
    oai32 CACHE_L0_1_L1_2_Fij_ix283 (.Y (CACHE_L0_1_L1_2_Fij_nx282), .A0 (nx3867
          ), .A1 (nx8387), .A2 (nx6993), .B0 (nx2627), .B1 (nx8687)) ;
    oai32 CACHE_L0_1_L1_2_Wij_ix213 (.Y (CACHE_L0_1_L1_2_Wij_nx212), .A0 (nx3733
          ), .A1 (nx8387), .A2 (nx6995), .B0 (nx2493), .B1 (nx8689)) ;
    inv02 ix6994 (.Y (nx6995), .A (CACHE_L0_1_L1_2_Wij_nx331)) ;
    oai32 CACHE_L0_1_L1_2_Wij_ix223 (.Y (CACHE_L0_1_L1_2_Wij_nx222), .A0 (nx3737
          ), .A1 (nx8387), .A2 (nx6995), .B0 (nx2497), .B1 (nx8689)) ;
    oai32 CACHE_L0_1_L1_2_Wij_ix233 (.Y (CACHE_L0_1_L1_2_Wij_nx232), .A0 (nx3741
          ), .A1 (nx8387), .A2 (nx6995), .B0 (nx2501), .B1 (nx8689)) ;
    oai32 CACHE_L0_1_L1_2_Wij_ix243 (.Y (CACHE_L0_1_L1_2_Wij_nx242), .A0 (nx3745
          ), .A1 (nx8387), .A2 (nx6995), .B0 (nx2505), .B1 (nx8689)) ;
    oai32 CACHE_L0_1_L1_2_Wij_ix253 (.Y (CACHE_L0_1_L1_2_Wij_nx252), .A0 (nx3749
          ), .A1 (CACHE_RST_dup_1226), .A2 (nx6995), .B0 (nx2509), .B1 (nx8689)
          ) ;
    oai32 CACHE_L0_1_L1_2_Wij_ix263 (.Y (CACHE_L0_1_L1_2_Wij_nx262), .A0 (nx3753
          ), .A1 (CACHE_RST_dup_1226), .A2 (nx6995), .B0 (nx2513), .B1 (nx8689)
          ) ;
    oai32 CACHE_L0_1_L1_2_Wij_ix273 (.Y (CACHE_L0_1_L1_2_Wij_nx272), .A0 (nx3757
          ), .A1 (CACHE_RST_dup_1226), .A2 (nx6999), .B0 (nx2517), .B1 (nx8689)
          ) ;
    inv01 ix6998 (.Y (nx6999), .A (CACHE_L0_1_L1_2_Wij_nx333)) ;
    oai32 CACHE_L0_1_L1_2_Wij_ix283 (.Y (CACHE_L0_1_L1_2_Wij_nx282), .A0 (nx3761
          ), .A1 (CACHE_RST_dup_1226), .A2 (nx6999), .B0 (nx2521), .B1 (nx8691)
          ) ;
    oai32 CACHE_L0_1_L1_3_Fij_ix213 (.Y (CACHE_L0_1_L1_3_Fij_nx212), .A0 (nx4099
          ), .A1 (nx8389), .A2 (nx7001), .B0 (nx2859), .B1 (nx8693)) ;
    inv02 ix7000 (.Y (nx7001), .A (CACHE_L0_1_L1_3_Fij_nx331)) ;
    oai32 CACHE_L0_1_L1_3_Fij_ix223 (.Y (CACHE_L0_1_L1_3_Fij_nx222), .A0 (nx4101
          ), .A1 (nx8389), .A2 (nx7001), .B0 (nx2861), .B1 (nx8693)) ;
    oai32 CACHE_L0_1_L1_3_Fij_ix233 (.Y (CACHE_L0_1_L1_3_Fij_nx232), .A0 (nx4103
          ), .A1 (nx8389), .A2 (nx7001), .B0 (nx2863), .B1 (nx8693)) ;
    oai32 CACHE_L0_1_L1_3_Fij_ix243 (.Y (CACHE_L0_1_L1_3_Fij_nx242), .A0 (nx4105
          ), .A1 (nx8389), .A2 (nx7001), .B0 (nx2865), .B1 (nx8693)) ;
    oai32 CACHE_L0_1_L1_3_Fij_ix253 (.Y (CACHE_L0_1_L1_3_Fij_nx252), .A0 (nx4107
          ), .A1 (nx8389), .A2 (nx7001), .B0 (nx2867), .B1 (nx8693)) ;
    oai32 CACHE_L0_1_L1_3_Fij_ix263 (.Y (CACHE_L0_1_L1_3_Fij_nx262), .A0 (nx4109
          ), .A1 (nx8391), .A2 (nx7001), .B0 (nx2869), .B1 (nx8693)) ;
    oai32 CACHE_L0_1_L1_3_Fij_ix273 (.Y (CACHE_L0_1_L1_3_Fij_nx272), .A0 (nx4113
          ), .A1 (nx8391), .A2 (nx7005), .B0 (nx2873), .B1 (nx8693)) ;
    inv01 ix7004 (.Y (nx7005), .A (CACHE_L0_1_L1_3_Fij_nx333)) ;
    oai32 CACHE_L0_1_L1_3_Fij_ix283 (.Y (CACHE_L0_1_L1_3_Fij_nx282), .A0 (nx4115
          ), .A1 (nx8391), .A2 (nx7005), .B0 (nx2875), .B1 (nx8695)) ;
    oai32 CACHE_L0_1_L1_3_Wij_ix213 (.Y (CACHE_L0_1_L1_3_Wij_nx212), .A0 (nx3981
          ), .A1 (nx8391), .A2 (nx7007), .B0 (nx2741), .B1 (nx8697)) ;
    inv02 ix7006 (.Y (nx7007), .A (CACHE_L0_1_L1_3_Wij_nx331)) ;
    oai32 CACHE_L0_1_L1_3_Wij_ix223 (.Y (CACHE_L0_1_L1_3_Wij_nx222), .A0 (nx3985
          ), .A1 (nx8391), .A2 (nx7007), .B0 (nx2745), .B1 (nx8697)) ;
    oai32 CACHE_L0_1_L1_3_Wij_ix233 (.Y (CACHE_L0_1_L1_3_Wij_nx232), .A0 (nx3989
          ), .A1 (nx8391), .A2 (nx7007), .B0 (nx2749), .B1 (nx8697)) ;
    oai32 CACHE_L0_1_L1_3_Wij_ix243 (.Y (CACHE_L0_1_L1_3_Wij_nx242), .A0 (nx3993
          ), .A1 (nx8391), .A2 (nx7007), .B0 (nx2753), .B1 (nx8697)) ;
    oai32 CACHE_L0_1_L1_3_Wij_ix253 (.Y (CACHE_L0_1_L1_3_Wij_nx252), .A0 (nx3997
          ), .A1 (CACHE_RST_dup_1248), .A2 (nx7007), .B0 (nx2757), .B1 (nx8697)
          ) ;
    oai32 CACHE_L0_1_L1_3_Wij_ix263 (.Y (CACHE_L0_1_L1_3_Wij_nx262), .A0 (nx4001
          ), .A1 (CACHE_RST_dup_1248), .A2 (nx7007), .B0 (nx2761), .B1 (nx8697)
          ) ;
    oai32 CACHE_L0_1_L1_3_Wij_ix273 (.Y (CACHE_L0_1_L1_3_Wij_nx272), .A0 (nx4005
          ), .A1 (CACHE_RST_dup_1248), .A2 (nx7011), .B0 (nx2765), .B1 (nx8697)
          ) ;
    inv01 ix7010 (.Y (nx7011), .A (CACHE_L0_1_L1_3_Wij_nx333)) ;
    oai32 CACHE_L0_1_L1_3_Wij_ix283 (.Y (CACHE_L0_1_L1_3_Wij_nx282), .A0 (nx4009
          ), .A1 (CACHE_RST_dup_1248), .A2 (nx7011), .B0 (nx2769), .B1 (nx8699)
          ) ;
    oai32 CACHE_L0_1_L1_4_Fij_ix213 (.Y (CACHE_L0_1_L1_4_Fij_nx212), .A0 (nx4347
          ), .A1 (nx8393), .A2 (nx7013), .B0 (nx3107), .B1 (nx8701)) ;
    inv02 ix7012 (.Y (nx7013), .A (CACHE_L0_1_L1_4_Fij_nx331)) ;
    oai32 CACHE_L0_1_L1_4_Fij_ix223 (.Y (CACHE_L0_1_L1_4_Fij_nx222), .A0 (nx4349
          ), .A1 (nx8393), .A2 (nx7013), .B0 (nx3109), .B1 (nx8701)) ;
    oai32 CACHE_L0_1_L1_4_Fij_ix233 (.Y (CACHE_L0_1_L1_4_Fij_nx232), .A0 (nx4351
          ), .A1 (nx8393), .A2 (nx7013), .B0 (nx3111), .B1 (nx8701)) ;
    oai32 CACHE_L0_1_L1_4_Fij_ix243 (.Y (CACHE_L0_1_L1_4_Fij_nx242), .A0 (nx4353
          ), .A1 (nx8393), .A2 (nx7013), .B0 (nx3113), .B1 (nx8701)) ;
    oai32 CACHE_L0_1_L1_4_Fij_ix253 (.Y (CACHE_L0_1_L1_4_Fij_nx252), .A0 (nx4355
          ), .A1 (nx8393), .A2 (nx7013), .B0 (nx3115), .B1 (nx8701)) ;
    oai32 CACHE_L0_1_L1_4_Fij_ix263 (.Y (CACHE_L0_1_L1_4_Fij_nx262), .A0 (nx4357
          ), .A1 (nx8395), .A2 (nx7013), .B0 (nx3117), .B1 (nx8701)) ;
    oai32 CACHE_L0_1_L1_4_Fij_ix273 (.Y (CACHE_L0_1_L1_4_Fij_nx272), .A0 (nx4361
          ), .A1 (nx8395), .A2 (nx7017), .B0 (nx3121), .B1 (nx8701)) ;
    inv01 ix7016 (.Y (nx7017), .A (CACHE_L0_1_L1_4_Fij_nx333)) ;
    oai32 CACHE_L0_1_L1_4_Fij_ix283 (.Y (CACHE_L0_1_L1_4_Fij_nx282), .A0 (nx4363
          ), .A1 (nx8395), .A2 (nx7017), .B0 (nx3123), .B1 (nx8703)) ;
    oai32 CACHE_L0_1_L1_4_Wij_ix213 (.Y (CACHE_L0_1_L1_4_Wij_nx212), .A0 (nx4229
          ), .A1 (nx8395), .A2 (nx7019), .B0 (nx2989), .B1 (nx8705)) ;
    inv02 ix7018 (.Y (nx7019), .A (CACHE_L0_1_L1_4_Wij_nx331)) ;
    oai32 CACHE_L0_1_L1_4_Wij_ix223 (.Y (CACHE_L0_1_L1_4_Wij_nx222), .A0 (nx4233
          ), .A1 (nx8395), .A2 (nx7019), .B0 (nx2993), .B1 (nx8705)) ;
    oai32 CACHE_L0_1_L1_4_Wij_ix233 (.Y (CACHE_L0_1_L1_4_Wij_nx232), .A0 (nx4237
          ), .A1 (nx8395), .A2 (nx7019), .B0 (nx2997), .B1 (nx8705)) ;
    oai32 CACHE_L0_1_L1_4_Wij_ix243 (.Y (CACHE_L0_1_L1_4_Wij_nx242), .A0 (nx4241
          ), .A1 (nx8395), .A2 (nx7019), .B0 (nx3001), .B1 (nx8705)) ;
    oai32 CACHE_L0_1_L1_4_Wij_ix253 (.Y (CACHE_L0_1_L1_4_Wij_nx252), .A0 (nx4245
          ), .A1 (CACHE_RST_dup_1270), .A2 (nx7019), .B0 (nx3005), .B1 (nx8705)
          ) ;
    oai32 CACHE_L0_1_L1_4_Wij_ix263 (.Y (CACHE_L0_1_L1_4_Wij_nx262), .A0 (nx4249
          ), .A1 (CACHE_RST_dup_1270), .A2 (nx7019), .B0 (nx3009), .B1 (nx8705)
          ) ;
    oai32 CACHE_L0_1_L1_4_Wij_ix273 (.Y (CACHE_L0_1_L1_4_Wij_nx272), .A0 (nx4253
          ), .A1 (CACHE_RST_dup_1270), .A2 (nx7023), .B0 (nx3013), .B1 (nx8705)
          ) ;
    inv01 ix7022 (.Y (nx7023), .A (CACHE_L0_1_L1_4_Wij_nx333)) ;
    oai32 CACHE_L0_1_L1_4_Wij_ix283 (.Y (CACHE_L0_1_L1_4_Wij_nx282), .A0 (nx4257
          ), .A1 (CACHE_RST_dup_1270), .A2 (nx7023), .B0 (nx3017), .B1 (nx8707)
          ) ;
    oai32 CACHE_L0_2_L1_0_Fij_ix213 (.Y (CACHE_L0_2_L1_0_Fij_nx212), .A0 (nx4595
          ), .A1 (nx8397), .A2 (nx7025), .B0 (nx3355), .B1 (nx8709)) ;
    inv02 ix7024 (.Y (nx7025), .A (CACHE_L0_2_L1_0_Fij_nx331)) ;
    oai32 CACHE_L0_2_L1_0_Fij_ix223 (.Y (CACHE_L0_2_L1_0_Fij_nx222), .A0 (nx4597
          ), .A1 (nx8397), .A2 (nx7025), .B0 (nx3357), .B1 (nx8709)) ;
    oai32 CACHE_L0_2_L1_0_Fij_ix233 (.Y (CACHE_L0_2_L1_0_Fij_nx232), .A0 (nx4599
          ), .A1 (nx8397), .A2 (nx7025), .B0 (nx3359), .B1 (nx8709)) ;
    oai32 CACHE_L0_2_L1_0_Fij_ix243 (.Y (CACHE_L0_2_L1_0_Fij_nx242), .A0 (nx4601
          ), .A1 (nx8397), .A2 (nx7025), .B0 (nx3361), .B1 (nx8709)) ;
    oai32 CACHE_L0_2_L1_0_Fij_ix253 (.Y (CACHE_L0_2_L1_0_Fij_nx252), .A0 (nx4603
          ), .A1 (nx8397), .A2 (nx7025), .B0 (nx3363), .B1 (nx8709)) ;
    oai32 CACHE_L0_2_L1_0_Fij_ix263 (.Y (CACHE_L0_2_L1_0_Fij_nx262), .A0 (nx4605
          ), .A1 (nx8399), .A2 (nx7025), .B0 (nx3365), .B1 (nx8709)) ;
    oai32 CACHE_L0_2_L1_0_Fij_ix273 (.Y (CACHE_L0_2_L1_0_Fij_nx272), .A0 (nx4609
          ), .A1 (nx8399), .A2 (nx7029), .B0 (nx3369), .B1 (nx8709)) ;
    inv01 ix7028 (.Y (nx7029), .A (CACHE_L0_2_L1_0_Fij_nx333)) ;
    oai32 CACHE_L0_2_L1_0_Fij_ix283 (.Y (CACHE_L0_2_L1_0_Fij_nx282), .A0 (nx4611
          ), .A1 (nx8399), .A2 (nx7029), .B0 (nx3371), .B1 (nx8711)) ;
    oai32 CACHE_L0_2_L1_0_Wij_ix213 (.Y (CACHE_L0_2_L1_0_Wij_nx212), .A0 (nx4477
          ), .A1 (nx8399), .A2 (nx7031), .B0 (nx3237), .B1 (nx8713)) ;
    inv02 ix7030 (.Y (nx7031), .A (CACHE_L0_2_L1_0_Wij_nx331)) ;
    oai32 CACHE_L0_2_L1_0_Wij_ix223 (.Y (CACHE_L0_2_L1_0_Wij_nx222), .A0 (nx4481
          ), .A1 (nx8399), .A2 (nx7031), .B0 (nx3241), .B1 (nx8713)) ;
    oai32 CACHE_L0_2_L1_0_Wij_ix233 (.Y (CACHE_L0_2_L1_0_Wij_nx232), .A0 (nx4485
          ), .A1 (nx8399), .A2 (nx7031), .B0 (nx3245), .B1 (nx8713)) ;
    oai32 CACHE_L0_2_L1_0_Wij_ix243 (.Y (CACHE_L0_2_L1_0_Wij_nx242), .A0 (nx4489
          ), .A1 (nx8399), .A2 (nx7031), .B0 (nx3249), .B1 (nx8713)) ;
    oai32 CACHE_L0_2_L1_0_Wij_ix253 (.Y (CACHE_L0_2_L1_0_Wij_nx252), .A0 (nx4493
          ), .A1 (CACHE_RST_dup_1292), .A2 (nx7031), .B0 (nx3253), .B1 (nx8713)
          ) ;
    oai32 CACHE_L0_2_L1_0_Wij_ix263 (.Y (CACHE_L0_2_L1_0_Wij_nx262), .A0 (nx4497
          ), .A1 (CACHE_RST_dup_1292), .A2 (nx7031), .B0 (nx3257), .B1 (nx8713)
          ) ;
    oai32 CACHE_L0_2_L1_0_Wij_ix273 (.Y (CACHE_L0_2_L1_0_Wij_nx272), .A0 (nx4501
          ), .A1 (CACHE_RST_dup_1292), .A2 (nx7035), .B0 (nx3261), .B1 (nx8713)
          ) ;
    inv01 ix7034 (.Y (nx7035), .A (CACHE_L0_2_L1_0_Wij_nx333)) ;
    oai32 CACHE_L0_2_L1_0_Wij_ix283 (.Y (CACHE_L0_2_L1_0_Wij_nx282), .A0 (nx4505
          ), .A1 (CACHE_RST_dup_1292), .A2 (nx7035), .B0 (nx3265), .B1 (nx8715)
          ) ;
    oai32 CACHE_L0_2_L1_1_Fij_ix213 (.Y (CACHE_L0_2_L1_1_Fij_nx212), .A0 (nx4843
          ), .A1 (nx8401), .A2 (nx7037), .B0 (nx3603), .B1 (nx8717)) ;
    inv02 ix7036 (.Y (nx7037), .A (CACHE_L0_2_L1_1_Fij_nx331)) ;
    oai32 CACHE_L0_2_L1_1_Fij_ix223 (.Y (CACHE_L0_2_L1_1_Fij_nx222), .A0 (nx4845
          ), .A1 (nx8401), .A2 (nx7037), .B0 (nx3605), .B1 (nx8717)) ;
    oai32 CACHE_L0_2_L1_1_Fij_ix233 (.Y (CACHE_L0_2_L1_1_Fij_nx232), .A0 (nx4847
          ), .A1 (nx8401), .A2 (nx7037), .B0 (nx3607), .B1 (nx8717)) ;
    oai32 CACHE_L0_2_L1_1_Fij_ix243 (.Y (CACHE_L0_2_L1_1_Fij_nx242), .A0 (nx4849
          ), .A1 (nx8401), .A2 (nx7037), .B0 (nx3609), .B1 (nx8717)) ;
    oai32 CACHE_L0_2_L1_1_Fij_ix253 (.Y (CACHE_L0_2_L1_1_Fij_nx252), .A0 (nx4851
          ), .A1 (nx8401), .A2 (nx7037), .B0 (nx3611), .B1 (nx8717)) ;
    oai32 CACHE_L0_2_L1_1_Fij_ix263 (.Y (CACHE_L0_2_L1_1_Fij_nx262), .A0 (nx4853
          ), .A1 (nx8403), .A2 (nx7037), .B0 (nx3613), .B1 (nx8717)) ;
    oai32 CACHE_L0_2_L1_1_Fij_ix273 (.Y (CACHE_L0_2_L1_1_Fij_nx272), .A0 (nx4857
          ), .A1 (nx8403), .A2 (nx7041), .B0 (nx3617), .B1 (nx8717)) ;
    inv01 ix7040 (.Y (nx7041), .A (CACHE_L0_2_L1_1_Fij_nx333)) ;
    oai32 CACHE_L0_2_L1_1_Fij_ix283 (.Y (CACHE_L0_2_L1_1_Fij_nx282), .A0 (nx4859
          ), .A1 (nx8403), .A2 (nx7041), .B0 (nx3619), .B1 (nx8719)) ;
    oai32 CACHE_L0_2_L1_1_Wij_ix213 (.Y (CACHE_L0_2_L1_1_Wij_nx212), .A0 (nx4725
          ), .A1 (nx8403), .A2 (nx7043), .B0 (nx3485), .B1 (nx8721)) ;
    inv02 ix7042 (.Y (nx7043), .A (CACHE_L0_2_L1_1_Wij_nx331)) ;
    oai32 CACHE_L0_2_L1_1_Wij_ix223 (.Y (CACHE_L0_2_L1_1_Wij_nx222), .A0 (nx4729
          ), .A1 (nx8403), .A2 (nx7043), .B0 (nx3489), .B1 (nx8721)) ;
    oai32 CACHE_L0_2_L1_1_Wij_ix233 (.Y (CACHE_L0_2_L1_1_Wij_nx232), .A0 (nx4733
          ), .A1 (nx8403), .A2 (nx7043), .B0 (nx3493), .B1 (nx8721)) ;
    oai32 CACHE_L0_2_L1_1_Wij_ix243 (.Y (CACHE_L0_2_L1_1_Wij_nx242), .A0 (nx4737
          ), .A1 (nx8403), .A2 (nx7043), .B0 (nx3497), .B1 (nx8721)) ;
    oai32 CACHE_L0_2_L1_1_Wij_ix253 (.Y (CACHE_L0_2_L1_1_Wij_nx252), .A0 (nx4741
          ), .A1 (CACHE_RST_dup_1314), .A2 (nx7043), .B0 (nx3501), .B1 (nx8721)
          ) ;
    oai32 CACHE_L0_2_L1_1_Wij_ix263 (.Y (CACHE_L0_2_L1_1_Wij_nx262), .A0 (nx4745
          ), .A1 (CACHE_RST_dup_1314), .A2 (nx7043), .B0 (nx3505), .B1 (nx8721)
          ) ;
    oai32 CACHE_L0_2_L1_1_Wij_ix273 (.Y (CACHE_L0_2_L1_1_Wij_nx272), .A0 (nx4749
          ), .A1 (CACHE_RST_dup_1314), .A2 (nx7047), .B0 (nx3509), .B1 (nx8721)
          ) ;
    inv01 ix7046 (.Y (nx7047), .A (CACHE_L0_2_L1_1_Wij_nx333)) ;
    oai32 CACHE_L0_2_L1_1_Wij_ix283 (.Y (CACHE_L0_2_L1_1_Wij_nx282), .A0 (nx4753
          ), .A1 (CACHE_RST_dup_1314), .A2 (nx7047), .B0 (nx3513), .B1 (nx8723)
          ) ;
    oai32 CACHE_L0_2_L1_2_Fij_ix213 (.Y (CACHE_L0_2_L1_2_Fij_nx212), .A0 (nx5091
          ), .A1 (nx8405), .A2 (nx7049), .B0 (nx3851), .B1 (nx8725)) ;
    inv02 ix7048 (.Y (nx7049), .A (CACHE_L0_2_L1_2_Fij_nx331)) ;
    oai32 CACHE_L0_2_L1_2_Fij_ix223 (.Y (CACHE_L0_2_L1_2_Fij_nx222), .A0 (nx5093
          ), .A1 (nx8405), .A2 (nx7049), .B0 (nx3853), .B1 (nx8725)) ;
    oai32 CACHE_L0_2_L1_2_Fij_ix233 (.Y (CACHE_L0_2_L1_2_Fij_nx232), .A0 (nx5095
          ), .A1 (nx8405), .A2 (nx7049), .B0 (nx3855), .B1 (nx8725)) ;
    oai32 CACHE_L0_2_L1_2_Fij_ix243 (.Y (CACHE_L0_2_L1_2_Fij_nx242), .A0 (nx5097
          ), .A1 (nx8405), .A2 (nx7049), .B0 (nx3857), .B1 (nx8725)) ;
    oai32 CACHE_L0_2_L1_2_Fij_ix253 (.Y (CACHE_L0_2_L1_2_Fij_nx252), .A0 (nx5099
          ), .A1 (nx8405), .A2 (nx7049), .B0 (nx3859), .B1 (nx8725)) ;
    oai32 CACHE_L0_2_L1_2_Fij_ix263 (.Y (CACHE_L0_2_L1_2_Fij_nx262), .A0 (nx5101
          ), .A1 (nx8407), .A2 (nx7049), .B0 (nx3861), .B1 (nx8725)) ;
    oai32 CACHE_L0_2_L1_2_Fij_ix273 (.Y (CACHE_L0_2_L1_2_Fij_nx272), .A0 (nx5105
          ), .A1 (nx8407), .A2 (nx7053), .B0 (nx3865), .B1 (nx8725)) ;
    inv01 ix7052 (.Y (nx7053), .A (CACHE_L0_2_L1_2_Fij_nx333)) ;
    oai32 CACHE_L0_2_L1_2_Fij_ix283 (.Y (CACHE_L0_2_L1_2_Fij_nx282), .A0 (nx5107
          ), .A1 (nx8407), .A2 (nx7053), .B0 (nx3867), .B1 (nx8727)) ;
    oai32 CACHE_L0_2_L1_2_Wij_ix213 (.Y (CACHE_L0_2_L1_2_Wij_nx212), .A0 (nx4973
          ), .A1 (nx8407), .A2 (nx7055), .B0 (nx3733), .B1 (nx8729)) ;
    inv02 ix7054 (.Y (nx7055), .A (CACHE_L0_2_L1_2_Wij_nx331)) ;
    oai32 CACHE_L0_2_L1_2_Wij_ix223 (.Y (CACHE_L0_2_L1_2_Wij_nx222), .A0 (nx4977
          ), .A1 (nx8407), .A2 (nx7055), .B0 (nx3737), .B1 (nx8729)) ;
    oai32 CACHE_L0_2_L1_2_Wij_ix233 (.Y (CACHE_L0_2_L1_2_Wij_nx232), .A0 (nx4981
          ), .A1 (nx8407), .A2 (nx7055), .B0 (nx3741), .B1 (nx8729)) ;
    oai32 CACHE_L0_2_L1_2_Wij_ix243 (.Y (CACHE_L0_2_L1_2_Wij_nx242), .A0 (nx4985
          ), .A1 (nx8407), .A2 (nx7055), .B0 (nx3745), .B1 (nx8729)) ;
    oai32 CACHE_L0_2_L1_2_Wij_ix253 (.Y (CACHE_L0_2_L1_2_Wij_nx252), .A0 (nx4989
          ), .A1 (CACHE_RST_dup_1336), .A2 (nx7055), .B0 (nx3749), .B1 (nx8729)
          ) ;
    oai32 CACHE_L0_2_L1_2_Wij_ix263 (.Y (CACHE_L0_2_L1_2_Wij_nx262), .A0 (nx4993
          ), .A1 (CACHE_RST_dup_1336), .A2 (nx7055), .B0 (nx3753), .B1 (nx8729)
          ) ;
    oai32 CACHE_L0_2_L1_2_Wij_ix273 (.Y (CACHE_L0_2_L1_2_Wij_nx272), .A0 (nx4997
          ), .A1 (CACHE_RST_dup_1336), .A2 (nx7059), .B0 (nx3757), .B1 (nx8729)
          ) ;
    inv01 ix7058 (.Y (nx7059), .A (CACHE_L0_2_L1_2_Wij_nx333)) ;
    oai32 CACHE_L0_2_L1_2_Wij_ix283 (.Y (CACHE_L0_2_L1_2_Wij_nx282), .A0 (nx5001
          ), .A1 (CACHE_RST_dup_1336), .A2 (nx7059), .B0 (nx3761), .B1 (nx8731)
          ) ;
    oai32 CACHE_L0_2_L1_3_Fij_ix213 (.Y (CACHE_L0_2_L1_3_Fij_nx212), .A0 (nx5339
          ), .A1 (nx8409), .A2 (nx7061), .B0 (nx4099), .B1 (nx8733)) ;
    inv02 ix7060 (.Y (nx7061), .A (CACHE_L0_2_L1_3_Fij_nx331)) ;
    oai32 CACHE_L0_2_L1_3_Fij_ix223 (.Y (CACHE_L0_2_L1_3_Fij_nx222), .A0 (nx5341
          ), .A1 (nx8409), .A2 (nx7061), .B0 (nx4101), .B1 (nx8733)) ;
    oai32 CACHE_L0_2_L1_3_Fij_ix233 (.Y (CACHE_L0_2_L1_3_Fij_nx232), .A0 (nx5343
          ), .A1 (nx8409), .A2 (nx7061), .B0 (nx4103), .B1 (nx8733)) ;
    oai32 CACHE_L0_2_L1_3_Fij_ix243 (.Y (CACHE_L0_2_L1_3_Fij_nx242), .A0 (nx5345
          ), .A1 (nx8409), .A2 (nx7061), .B0 (nx4105), .B1 (nx8733)) ;
    oai32 CACHE_L0_2_L1_3_Fij_ix253 (.Y (CACHE_L0_2_L1_3_Fij_nx252), .A0 (nx5347
          ), .A1 (nx8409), .A2 (nx7061), .B0 (nx4107), .B1 (nx8733)) ;
    oai32 CACHE_L0_2_L1_3_Fij_ix263 (.Y (CACHE_L0_2_L1_3_Fij_nx262), .A0 (nx5349
          ), .A1 (nx8411), .A2 (nx7061), .B0 (nx4109), .B1 (nx8733)) ;
    oai32 CACHE_L0_2_L1_3_Fij_ix273 (.Y (CACHE_L0_2_L1_3_Fij_nx272), .A0 (nx5353
          ), .A1 (nx8411), .A2 (nx7065), .B0 (nx4113), .B1 (nx8733)) ;
    inv01 ix7064 (.Y (nx7065), .A (CACHE_L0_2_L1_3_Fij_nx333)) ;
    oai32 CACHE_L0_2_L1_3_Fij_ix283 (.Y (CACHE_L0_2_L1_3_Fij_nx282), .A0 (nx5355
          ), .A1 (nx8411), .A2 (nx7065), .B0 (nx4115), .B1 (nx8735)) ;
    oai32 CACHE_L0_2_L1_3_Wij_ix213 (.Y (CACHE_L0_2_L1_3_Wij_nx212), .A0 (nx5221
          ), .A1 (nx8411), .A2 (nx7067), .B0 (nx3981), .B1 (nx8737)) ;
    inv02 ix7066 (.Y (nx7067), .A (CACHE_L0_2_L1_3_Wij_nx331)) ;
    oai32 CACHE_L0_2_L1_3_Wij_ix223 (.Y (CACHE_L0_2_L1_3_Wij_nx222), .A0 (nx5225
          ), .A1 (nx8411), .A2 (nx7067), .B0 (nx3985), .B1 (nx8737)) ;
    oai32 CACHE_L0_2_L1_3_Wij_ix233 (.Y (CACHE_L0_2_L1_3_Wij_nx232), .A0 (nx5229
          ), .A1 (nx8411), .A2 (nx7067), .B0 (nx3989), .B1 (nx8737)) ;
    oai32 CACHE_L0_2_L1_3_Wij_ix243 (.Y (CACHE_L0_2_L1_3_Wij_nx242), .A0 (nx5233
          ), .A1 (nx8411), .A2 (nx7067), .B0 (nx3993), .B1 (nx8737)) ;
    oai32 CACHE_L0_2_L1_3_Wij_ix253 (.Y (CACHE_L0_2_L1_3_Wij_nx252), .A0 (nx5237
          ), .A1 (CACHE_RST_dup_1358), .A2 (nx7067), .B0 (nx3997), .B1 (nx8737)
          ) ;
    oai32 CACHE_L0_2_L1_3_Wij_ix263 (.Y (CACHE_L0_2_L1_3_Wij_nx262), .A0 (nx5241
          ), .A1 (CACHE_RST_dup_1358), .A2 (nx7067), .B0 (nx4001), .B1 (nx8737)
          ) ;
    oai32 CACHE_L0_2_L1_3_Wij_ix273 (.Y (CACHE_L0_2_L1_3_Wij_nx272), .A0 (nx5245
          ), .A1 (CACHE_RST_dup_1358), .A2 (nx7071), .B0 (nx4005), .B1 (nx8737)
          ) ;
    inv01 ix7070 (.Y (nx7071), .A (CACHE_L0_2_L1_3_Wij_nx333)) ;
    oai32 CACHE_L0_2_L1_3_Wij_ix283 (.Y (CACHE_L0_2_L1_3_Wij_nx282), .A0 (nx5249
          ), .A1 (CACHE_RST_dup_1358), .A2 (nx7071), .B0 (nx4009), .B1 (nx8739)
          ) ;
    oai32 CACHE_L0_2_L1_4_Fij_ix213 (.Y (CACHE_L0_2_L1_4_Fij_nx212), .A0 (nx5587
          ), .A1 (nx8413), .A2 (nx7073), .B0 (nx4347), .B1 (nx8741)) ;
    inv02 ix7072 (.Y (nx7073), .A (CACHE_L0_2_L1_4_Fij_nx331)) ;
    oai32 CACHE_L0_2_L1_4_Fij_ix223 (.Y (CACHE_L0_2_L1_4_Fij_nx222), .A0 (nx5589
          ), .A1 (nx8413), .A2 (nx7073), .B0 (nx4349), .B1 (nx8741)) ;
    oai32 CACHE_L0_2_L1_4_Fij_ix233 (.Y (CACHE_L0_2_L1_4_Fij_nx232), .A0 (nx5591
          ), .A1 (nx8413), .A2 (nx7073), .B0 (nx4351), .B1 (nx8741)) ;
    oai32 CACHE_L0_2_L1_4_Fij_ix243 (.Y (CACHE_L0_2_L1_4_Fij_nx242), .A0 (nx5593
          ), .A1 (nx8413), .A2 (nx7073), .B0 (nx4353), .B1 (nx8741)) ;
    oai32 CACHE_L0_2_L1_4_Fij_ix253 (.Y (CACHE_L0_2_L1_4_Fij_nx252), .A0 (nx5595
          ), .A1 (nx8413), .A2 (nx7073), .B0 (nx4355), .B1 (nx8741)) ;
    oai32 CACHE_L0_2_L1_4_Fij_ix263 (.Y (CACHE_L0_2_L1_4_Fij_nx262), .A0 (nx5597
          ), .A1 (nx8415), .A2 (nx7073), .B0 (nx4357), .B1 (nx8741)) ;
    oai32 CACHE_L0_2_L1_4_Fij_ix273 (.Y (CACHE_L0_2_L1_4_Fij_nx272), .A0 (nx5601
          ), .A1 (nx8415), .A2 (nx7077), .B0 (nx4361), .B1 (nx8741)) ;
    inv01 ix7076 (.Y (nx7077), .A (CACHE_L0_2_L1_4_Fij_nx333)) ;
    oai32 CACHE_L0_2_L1_4_Fij_ix283 (.Y (CACHE_L0_2_L1_4_Fij_nx282), .A0 (nx5603
          ), .A1 (nx8415), .A2 (nx7077), .B0 (nx4363), .B1 (nx8743)) ;
    oai32 CACHE_L0_2_L1_4_Wij_ix213 (.Y (CACHE_L0_2_L1_4_Wij_nx212), .A0 (nx5469
          ), .A1 (nx8415), .A2 (nx7079), .B0 (nx4229), .B1 (nx8745)) ;
    inv02 ix7078 (.Y (nx7079), .A (CACHE_L0_2_L1_4_Wij_nx331)) ;
    oai32 CACHE_L0_2_L1_4_Wij_ix223 (.Y (CACHE_L0_2_L1_4_Wij_nx222), .A0 (nx5473
          ), .A1 (nx8415), .A2 (nx7079), .B0 (nx4233), .B1 (nx8745)) ;
    oai32 CACHE_L0_2_L1_4_Wij_ix233 (.Y (CACHE_L0_2_L1_4_Wij_nx232), .A0 (nx5477
          ), .A1 (nx8415), .A2 (nx7079), .B0 (nx4237), .B1 (nx8745)) ;
    oai32 CACHE_L0_2_L1_4_Wij_ix243 (.Y (CACHE_L0_2_L1_4_Wij_nx242), .A0 (nx5481
          ), .A1 (nx8415), .A2 (nx7079), .B0 (nx4241), .B1 (nx8745)) ;
    oai32 CACHE_L0_2_L1_4_Wij_ix253 (.Y (CACHE_L0_2_L1_4_Wij_nx252), .A0 (nx5485
          ), .A1 (CACHE_RST_dup_1380), .A2 (nx7079), .B0 (nx4245), .B1 (nx8745)
          ) ;
    oai32 CACHE_L0_2_L1_4_Wij_ix263 (.Y (CACHE_L0_2_L1_4_Wij_nx262), .A0 (nx5489
          ), .A1 (CACHE_RST_dup_1380), .A2 (nx7079), .B0 (nx4249), .B1 (nx8745)
          ) ;
    oai32 CACHE_L0_2_L1_4_Wij_ix273 (.Y (CACHE_L0_2_L1_4_Wij_nx272), .A0 (nx5493
          ), .A1 (CACHE_RST_dup_1380), .A2 (nx7083), .B0 (nx4253), .B1 (nx8745)
          ) ;
    inv01 ix7082 (.Y (nx7083), .A (CACHE_L0_2_L1_4_Wij_nx333)) ;
    oai32 CACHE_L0_2_L1_4_Wij_ix283 (.Y (CACHE_L0_2_L1_4_Wij_nx282), .A0 (nx5497
          ), .A1 (CACHE_RST_dup_1380), .A2 (nx7083), .B0 (nx4257), .B1 (nx8747)
          ) ;
    oai32 CACHE_L0_3_L1_0_Fij_ix213 (.Y (CACHE_L0_3_L1_0_Fij_nx212), .A0 (nx5835
          ), .A1 (nx8417), .A2 (nx7085), .B0 (nx4595), .B1 (nx8749)) ;
    inv02 ix7084 (.Y (nx7085), .A (CACHE_L0_3_L1_0_Fij_nx331)) ;
    oai32 CACHE_L0_3_L1_0_Fij_ix223 (.Y (CACHE_L0_3_L1_0_Fij_nx222), .A0 (nx5837
          ), .A1 (nx8417), .A2 (nx7085), .B0 (nx4597), .B1 (nx8749)) ;
    oai32 CACHE_L0_3_L1_0_Fij_ix233 (.Y (CACHE_L0_3_L1_0_Fij_nx232), .A0 (nx5839
          ), .A1 (nx8417), .A2 (nx7085), .B0 (nx4599), .B1 (nx8749)) ;
    oai32 CACHE_L0_3_L1_0_Fij_ix243 (.Y (CACHE_L0_3_L1_0_Fij_nx242), .A0 (nx5841
          ), .A1 (nx8417), .A2 (nx7085), .B0 (nx4601), .B1 (nx8749)) ;
    oai32 CACHE_L0_3_L1_0_Fij_ix253 (.Y (CACHE_L0_3_L1_0_Fij_nx252), .A0 (nx5843
          ), .A1 (nx8417), .A2 (nx7085), .B0 (nx4603), .B1 (nx8749)) ;
    oai32 CACHE_L0_3_L1_0_Fij_ix263 (.Y (CACHE_L0_3_L1_0_Fij_nx262), .A0 (nx5845
          ), .A1 (nx8419), .A2 (nx7085), .B0 (nx4605), .B1 (nx8749)) ;
    oai32 CACHE_L0_3_L1_0_Fij_ix273 (.Y (CACHE_L0_3_L1_0_Fij_nx272), .A0 (nx5849
          ), .A1 (nx8419), .A2 (nx7089), .B0 (nx4609), .B1 (nx8749)) ;
    inv01 ix7088 (.Y (nx7089), .A (CACHE_L0_3_L1_0_Fij_nx333)) ;
    oai32 CACHE_L0_3_L1_0_Fij_ix283 (.Y (CACHE_L0_3_L1_0_Fij_nx282), .A0 (nx5851
          ), .A1 (nx8419), .A2 (nx7089), .B0 (nx4611), .B1 (nx8751)) ;
    oai32 CACHE_L0_3_L1_0_Wij_ix213 (.Y (CACHE_L0_3_L1_0_Wij_nx212), .A0 (nx5717
          ), .A1 (nx8419), .A2 (nx7091), .B0 (nx4477), .B1 (nx8753)) ;
    inv02 ix7090 (.Y (nx7091), .A (CACHE_L0_3_L1_0_Wij_nx331)) ;
    oai32 CACHE_L0_3_L1_0_Wij_ix223 (.Y (CACHE_L0_3_L1_0_Wij_nx222), .A0 (nx5721
          ), .A1 (nx8419), .A2 (nx7091), .B0 (nx4481), .B1 (nx8753)) ;
    oai32 CACHE_L0_3_L1_0_Wij_ix233 (.Y (CACHE_L0_3_L1_0_Wij_nx232), .A0 (nx5725
          ), .A1 (nx8419), .A2 (nx7091), .B0 (nx4485), .B1 (nx8753)) ;
    oai32 CACHE_L0_3_L1_0_Wij_ix243 (.Y (CACHE_L0_3_L1_0_Wij_nx242), .A0 (nx5729
          ), .A1 (nx8419), .A2 (nx7091), .B0 (nx4489), .B1 (nx8753)) ;
    oai32 CACHE_L0_3_L1_0_Wij_ix253 (.Y (CACHE_L0_3_L1_0_Wij_nx252), .A0 (nx5733
          ), .A1 (CACHE_RST_dup_1402), .A2 (nx7091), .B0 (nx4493), .B1 (nx8753)
          ) ;
    oai32 CACHE_L0_3_L1_0_Wij_ix263 (.Y (CACHE_L0_3_L1_0_Wij_nx262), .A0 (nx5737
          ), .A1 (CACHE_RST_dup_1402), .A2 (nx7091), .B0 (nx4497), .B1 (nx8753)
          ) ;
    oai32 CACHE_L0_3_L1_0_Wij_ix273 (.Y (CACHE_L0_3_L1_0_Wij_nx272), .A0 (nx5741
          ), .A1 (CACHE_RST_dup_1402), .A2 (nx7095), .B0 (nx4501), .B1 (nx8753)
          ) ;
    inv01 ix7094 (.Y (nx7095), .A (CACHE_L0_3_L1_0_Wij_nx333)) ;
    oai32 CACHE_L0_3_L1_0_Wij_ix283 (.Y (CACHE_L0_3_L1_0_Wij_nx282), .A0 (nx5745
          ), .A1 (CACHE_RST_dup_1402), .A2 (nx7095), .B0 (nx4505), .B1 (nx8755)
          ) ;
    oai32 CACHE_L0_3_L1_1_Fij_ix213 (.Y (CACHE_L0_3_L1_1_Fij_nx212), .A0 (nx6083
          ), .A1 (nx8421), .A2 (nx7097), .B0 (nx4843), .B1 (nx8757)) ;
    inv02 ix7096 (.Y (nx7097), .A (CACHE_L0_3_L1_1_Fij_nx331)) ;
    oai32 CACHE_L0_3_L1_1_Fij_ix223 (.Y (CACHE_L0_3_L1_1_Fij_nx222), .A0 (nx6085
          ), .A1 (nx8421), .A2 (nx7097), .B0 (nx4845), .B1 (nx8757)) ;
    oai32 CACHE_L0_3_L1_1_Fij_ix233 (.Y (CACHE_L0_3_L1_1_Fij_nx232), .A0 (nx6087
          ), .A1 (nx8421), .A2 (nx7097), .B0 (nx4847), .B1 (nx8757)) ;
    oai32 CACHE_L0_3_L1_1_Fij_ix243 (.Y (CACHE_L0_3_L1_1_Fij_nx242), .A0 (nx6089
          ), .A1 (nx8421), .A2 (nx7097), .B0 (nx4849), .B1 (nx8757)) ;
    oai32 CACHE_L0_3_L1_1_Fij_ix253 (.Y (CACHE_L0_3_L1_1_Fij_nx252), .A0 (nx6091
          ), .A1 (nx8421), .A2 (nx7097), .B0 (nx4851), .B1 (nx8757)) ;
    oai32 CACHE_L0_3_L1_1_Fij_ix263 (.Y (CACHE_L0_3_L1_1_Fij_nx262), .A0 (nx6093
          ), .A1 (nx8423), .A2 (nx7097), .B0 (nx4853), .B1 (nx8757)) ;
    oai32 CACHE_L0_3_L1_1_Fij_ix273 (.Y (CACHE_L0_3_L1_1_Fij_nx272), .A0 (nx6097
          ), .A1 (nx8423), .A2 (nx7101), .B0 (nx4857), .B1 (nx8757)) ;
    inv01 ix7100 (.Y (nx7101), .A (CACHE_L0_3_L1_1_Fij_nx333)) ;
    oai32 CACHE_L0_3_L1_1_Fij_ix283 (.Y (CACHE_L0_3_L1_1_Fij_nx282), .A0 (nx6099
          ), .A1 (nx8423), .A2 (nx7101), .B0 (nx4859), .B1 (nx8759)) ;
    oai32 CACHE_L0_3_L1_1_Wij_ix213 (.Y (CACHE_L0_3_L1_1_Wij_nx212), .A0 (nx5965
          ), .A1 (nx8423), .A2 (nx7103), .B0 (nx4725), .B1 (nx8761)) ;
    inv02 ix7102 (.Y (nx7103), .A (CACHE_L0_3_L1_1_Wij_nx331)) ;
    oai32 CACHE_L0_3_L1_1_Wij_ix223 (.Y (CACHE_L0_3_L1_1_Wij_nx222), .A0 (nx5969
          ), .A1 (nx8423), .A2 (nx7103), .B0 (nx4729), .B1 (nx8761)) ;
    oai32 CACHE_L0_3_L1_1_Wij_ix233 (.Y (CACHE_L0_3_L1_1_Wij_nx232), .A0 (nx5973
          ), .A1 (nx8423), .A2 (nx7103), .B0 (nx4733), .B1 (nx8761)) ;
    oai32 CACHE_L0_3_L1_1_Wij_ix243 (.Y (CACHE_L0_3_L1_1_Wij_nx242), .A0 (nx5977
          ), .A1 (nx8423), .A2 (nx7103), .B0 (nx4737), .B1 (nx8761)) ;
    oai32 CACHE_L0_3_L1_1_Wij_ix253 (.Y (CACHE_L0_3_L1_1_Wij_nx252), .A0 (nx5981
          ), .A1 (CACHE_RST_dup_1424), .A2 (nx7103), .B0 (nx4741), .B1 (nx8761)
          ) ;
    oai32 CACHE_L0_3_L1_1_Wij_ix263 (.Y (CACHE_L0_3_L1_1_Wij_nx262), .A0 (nx5985
          ), .A1 (CACHE_RST_dup_1424), .A2 (nx7103), .B0 (nx4745), .B1 (nx8761)
          ) ;
    oai32 CACHE_L0_3_L1_1_Wij_ix273 (.Y (CACHE_L0_3_L1_1_Wij_nx272), .A0 (nx5989
          ), .A1 (CACHE_RST_dup_1424), .A2 (nx7107), .B0 (nx4749), .B1 (nx8761)
          ) ;
    inv01 ix7106 (.Y (nx7107), .A (CACHE_L0_3_L1_1_Wij_nx333)) ;
    oai32 CACHE_L0_3_L1_1_Wij_ix283 (.Y (CACHE_L0_3_L1_1_Wij_nx282), .A0 (nx5993
          ), .A1 (CACHE_RST_dup_1424), .A2 (nx7107), .B0 (nx4753), .B1 (nx8763)
          ) ;
    oai32 CACHE_L0_3_L1_2_Fij_ix213 (.Y (CACHE_L0_3_L1_2_Fij_nx212), .A0 (nx6331
          ), .A1 (nx8425), .A2 (nx7109), .B0 (nx5091), .B1 (nx8765)) ;
    inv02 ix7108 (.Y (nx7109), .A (CACHE_L0_3_L1_2_Fij_nx331)) ;
    oai32 CACHE_L0_3_L1_2_Fij_ix223 (.Y (CACHE_L0_3_L1_2_Fij_nx222), .A0 (nx6333
          ), .A1 (nx8425), .A2 (nx7109), .B0 (nx5093), .B1 (nx8765)) ;
    oai32 CACHE_L0_3_L1_2_Fij_ix233 (.Y (CACHE_L0_3_L1_2_Fij_nx232), .A0 (nx6335
          ), .A1 (nx8425), .A2 (nx7109), .B0 (nx5095), .B1 (nx8765)) ;
    oai32 CACHE_L0_3_L1_2_Fij_ix243 (.Y (CACHE_L0_3_L1_2_Fij_nx242), .A0 (nx6337
          ), .A1 (nx8425), .A2 (nx7109), .B0 (nx5097), .B1 (nx8765)) ;
    oai32 CACHE_L0_3_L1_2_Fij_ix253 (.Y (CACHE_L0_3_L1_2_Fij_nx252), .A0 (nx6339
          ), .A1 (nx8425), .A2 (nx7109), .B0 (nx5099), .B1 (nx8765)) ;
    oai32 CACHE_L0_3_L1_2_Fij_ix263 (.Y (CACHE_L0_3_L1_2_Fij_nx262), .A0 (nx6341
          ), .A1 (nx8427), .A2 (nx7109), .B0 (nx5101), .B1 (nx8765)) ;
    oai32 CACHE_L0_3_L1_2_Fij_ix273 (.Y (CACHE_L0_3_L1_2_Fij_nx272), .A0 (nx6345
          ), .A1 (nx8427), .A2 (nx7113), .B0 (nx5105), .B1 (nx8765)) ;
    inv01 ix7112 (.Y (nx7113), .A (CACHE_L0_3_L1_2_Fij_nx333)) ;
    oai32 CACHE_L0_3_L1_2_Fij_ix283 (.Y (CACHE_L0_3_L1_2_Fij_nx282), .A0 (nx6347
          ), .A1 (nx8427), .A2 (nx7113), .B0 (nx5107), .B1 (nx8767)) ;
    oai32 CACHE_L0_3_L1_2_Wij_ix213 (.Y (CACHE_L0_3_L1_2_Wij_nx212), .A0 (nx6213
          ), .A1 (nx8427), .A2 (nx7115), .B0 (nx4973), .B1 (nx8769)) ;
    inv02 ix7114 (.Y (nx7115), .A (CACHE_L0_3_L1_2_Wij_nx331)) ;
    oai32 CACHE_L0_3_L1_2_Wij_ix223 (.Y (CACHE_L0_3_L1_2_Wij_nx222), .A0 (nx6217
          ), .A1 (nx8427), .A2 (nx7115), .B0 (nx4977), .B1 (nx8769)) ;
    oai32 CACHE_L0_3_L1_2_Wij_ix233 (.Y (CACHE_L0_3_L1_2_Wij_nx232), .A0 (nx6221
          ), .A1 (nx8427), .A2 (nx7115), .B0 (nx4981), .B1 (nx8769)) ;
    oai32 CACHE_L0_3_L1_2_Wij_ix243 (.Y (CACHE_L0_3_L1_2_Wij_nx242), .A0 (nx6225
          ), .A1 (nx8427), .A2 (nx7115), .B0 (nx4985), .B1 (nx8769)) ;
    oai32 CACHE_L0_3_L1_2_Wij_ix253 (.Y (CACHE_L0_3_L1_2_Wij_nx252), .A0 (nx6229
          ), .A1 (CACHE_RST_dup_1446), .A2 (nx7115), .B0 (nx4989), .B1 (nx8769)
          ) ;
    oai32 CACHE_L0_3_L1_2_Wij_ix263 (.Y (CACHE_L0_3_L1_2_Wij_nx262), .A0 (nx6233
          ), .A1 (CACHE_RST_dup_1446), .A2 (nx7115), .B0 (nx4993), .B1 (nx8769)
          ) ;
    oai32 CACHE_L0_3_L1_2_Wij_ix273 (.Y (CACHE_L0_3_L1_2_Wij_nx272), .A0 (nx6237
          ), .A1 (CACHE_RST_dup_1446), .A2 (nx7119), .B0 (nx4997), .B1 (nx8769)
          ) ;
    inv01 ix7118 (.Y (nx7119), .A (CACHE_L0_3_L1_2_Wij_nx333)) ;
    oai32 CACHE_L0_3_L1_2_Wij_ix283 (.Y (CACHE_L0_3_L1_2_Wij_nx282), .A0 (nx6241
          ), .A1 (CACHE_RST_dup_1446), .A2 (nx7119), .B0 (nx5001), .B1 (nx8771)
          ) ;
    oai32 CACHE_L0_3_L1_3_Fij_ix213 (.Y (CACHE_L0_3_L1_3_Fij_nx212), .A0 (nx6579
          ), .A1 (nx8429), .A2 (nx7121), .B0 (nx5339), .B1 (nx8773)) ;
    inv02 ix7120 (.Y (nx7121), .A (CACHE_L0_3_L1_3_Fij_nx331)) ;
    oai32 CACHE_L0_3_L1_3_Fij_ix223 (.Y (CACHE_L0_3_L1_3_Fij_nx222), .A0 (nx6581
          ), .A1 (nx8429), .A2 (nx7121), .B0 (nx5341), .B1 (nx8773)) ;
    oai32 CACHE_L0_3_L1_3_Fij_ix233 (.Y (CACHE_L0_3_L1_3_Fij_nx232), .A0 (nx6583
          ), .A1 (nx8429), .A2 (nx7121), .B0 (nx5343), .B1 (nx8773)) ;
    oai32 CACHE_L0_3_L1_3_Fij_ix243 (.Y (CACHE_L0_3_L1_3_Fij_nx242), .A0 (nx6585
          ), .A1 (nx8429), .A2 (nx7121), .B0 (nx5345), .B1 (nx8773)) ;
    oai32 CACHE_L0_3_L1_3_Fij_ix253 (.Y (CACHE_L0_3_L1_3_Fij_nx252), .A0 (nx6587
          ), .A1 (nx8429), .A2 (nx7121), .B0 (nx5347), .B1 (nx8773)) ;
    oai32 CACHE_L0_3_L1_3_Fij_ix263 (.Y (CACHE_L0_3_L1_3_Fij_nx262), .A0 (nx6589
          ), .A1 (nx8431), .A2 (nx7121), .B0 (nx5349), .B1 (nx8773)) ;
    oai32 CACHE_L0_3_L1_3_Fij_ix273 (.Y (CACHE_L0_3_L1_3_Fij_nx272), .A0 (nx6593
          ), .A1 (nx8431), .A2 (nx7125), .B0 (nx5353), .B1 (nx8773)) ;
    inv01 ix7124 (.Y (nx7125), .A (CACHE_L0_3_L1_3_Fij_nx333)) ;
    oai32 CACHE_L0_3_L1_3_Fij_ix283 (.Y (CACHE_L0_3_L1_3_Fij_nx282), .A0 (nx6595
          ), .A1 (nx8431), .A2 (nx7125), .B0 (nx5355), .B1 (nx8775)) ;
    oai32 CACHE_L0_3_L1_3_Wij_ix213 (.Y (CACHE_L0_3_L1_3_Wij_nx212), .A0 (nx6461
          ), .A1 (nx8431), .A2 (nx7127), .B0 (nx5221), .B1 (nx8777)) ;
    inv02 ix7126 (.Y (nx7127), .A (CACHE_L0_3_L1_3_Wij_nx331)) ;
    oai32 CACHE_L0_3_L1_3_Wij_ix223 (.Y (CACHE_L0_3_L1_3_Wij_nx222), .A0 (nx6465
          ), .A1 (nx8431), .A2 (nx7127), .B0 (nx5225), .B1 (nx8777)) ;
    oai32 CACHE_L0_3_L1_3_Wij_ix233 (.Y (CACHE_L0_3_L1_3_Wij_nx232), .A0 (nx6469
          ), .A1 (nx8431), .A2 (nx7127), .B0 (nx5229), .B1 (nx8777)) ;
    oai32 CACHE_L0_3_L1_3_Wij_ix243 (.Y (CACHE_L0_3_L1_3_Wij_nx242), .A0 (nx6473
          ), .A1 (nx8431), .A2 (nx7127), .B0 (nx5233), .B1 (nx8777)) ;
    oai32 CACHE_L0_3_L1_3_Wij_ix253 (.Y (CACHE_L0_3_L1_3_Wij_nx252), .A0 (nx6477
          ), .A1 (CACHE_RST_dup_1468), .A2 (nx7127), .B0 (nx5237), .B1 (nx8777)
          ) ;
    oai32 CACHE_L0_3_L1_3_Wij_ix263 (.Y (CACHE_L0_3_L1_3_Wij_nx262), .A0 (nx6481
          ), .A1 (CACHE_RST_dup_1468), .A2 (nx7127), .B0 (nx5241), .B1 (nx8777)
          ) ;
    oai32 CACHE_L0_3_L1_3_Wij_ix273 (.Y (CACHE_L0_3_L1_3_Wij_nx272), .A0 (nx6485
          ), .A1 (CACHE_RST_dup_1468), .A2 (nx7131), .B0 (nx5245), .B1 (nx8777)
          ) ;
    inv01 ix7130 (.Y (nx7131), .A (CACHE_L0_3_L1_3_Wij_nx333)) ;
    oai32 CACHE_L0_3_L1_3_Wij_ix283 (.Y (CACHE_L0_3_L1_3_Wij_nx282), .A0 (nx6489
          ), .A1 (CACHE_RST_dup_1468), .A2 (nx7131), .B0 (nx5249), .B1 (nx8779)
          ) ;
    oai32 CACHE_L0_3_L1_4_Fij_ix213 (.Y (CACHE_L0_3_L1_4_Fij_nx212), .A0 (nx6827
          ), .A1 (nx8433), .A2 (nx7133), .B0 (nx5587), .B1 (nx8781)) ;
    inv02 ix7132 (.Y (nx7133), .A (CACHE_L0_3_L1_4_Fij_nx331)) ;
    oai32 CACHE_L0_3_L1_4_Fij_ix223 (.Y (CACHE_L0_3_L1_4_Fij_nx222), .A0 (nx6829
          ), .A1 (nx8433), .A2 (nx7133), .B0 (nx5589), .B1 (nx8781)) ;
    oai32 CACHE_L0_3_L1_4_Fij_ix233 (.Y (CACHE_L0_3_L1_4_Fij_nx232), .A0 (nx6831
          ), .A1 (nx8433), .A2 (nx7133), .B0 (nx5591), .B1 (nx8781)) ;
    oai32 CACHE_L0_3_L1_4_Fij_ix243 (.Y (CACHE_L0_3_L1_4_Fij_nx242), .A0 (nx6833
          ), .A1 (nx8433), .A2 (nx7133), .B0 (nx5593), .B1 (nx8781)) ;
    oai32 CACHE_L0_3_L1_4_Fij_ix253 (.Y (CACHE_L0_3_L1_4_Fij_nx252), .A0 (nx6835
          ), .A1 (nx8433), .A2 (nx7133), .B0 (nx5595), .B1 (nx8781)) ;
    oai32 CACHE_L0_3_L1_4_Fij_ix263 (.Y (CACHE_L0_3_L1_4_Fij_nx262), .A0 (nx6837
          ), .A1 (nx8435), .A2 (nx7133), .B0 (nx5597), .B1 (nx8781)) ;
    oai32 CACHE_L0_3_L1_4_Fij_ix273 (.Y (CACHE_L0_3_L1_4_Fij_nx272), .A0 (nx6841
          ), .A1 (nx8435), .A2 (nx7137), .B0 (nx5601), .B1 (nx8781)) ;
    inv01 ix7136 (.Y (nx7137), .A (CACHE_L0_3_L1_4_Fij_nx333)) ;
    oai32 CACHE_L0_3_L1_4_Fij_ix283 (.Y (CACHE_L0_3_L1_4_Fij_nx282), .A0 (nx6843
          ), .A1 (nx8435), .A2 (nx7137), .B0 (nx5603), .B1 (nx8783)) ;
    oai32 CACHE_L0_3_L1_4_Wij_ix213 (.Y (CACHE_L0_3_L1_4_Wij_nx212), .A0 (nx6709
          ), .A1 (nx8435), .A2 (nx7139), .B0 (nx5469), .B1 (nx8785)) ;
    inv02 ix7138 (.Y (nx7139), .A (CACHE_L0_3_L1_4_Wij_nx331)) ;
    oai32 CACHE_L0_3_L1_4_Wij_ix223 (.Y (CACHE_L0_3_L1_4_Wij_nx222), .A0 (nx6713
          ), .A1 (nx8435), .A2 (nx7139), .B0 (nx5473), .B1 (nx8785)) ;
    oai32 CACHE_L0_3_L1_4_Wij_ix233 (.Y (CACHE_L0_3_L1_4_Wij_nx232), .A0 (nx6717
          ), .A1 (nx8435), .A2 (nx7139), .B0 (nx5477), .B1 (nx8785)) ;
    oai32 CACHE_L0_3_L1_4_Wij_ix243 (.Y (CACHE_L0_3_L1_4_Wij_nx242), .A0 (nx6721
          ), .A1 (nx8435), .A2 (nx7139), .B0 (nx5481), .B1 (nx8785)) ;
    oai32 CACHE_L0_3_L1_4_Wij_ix253 (.Y (CACHE_L0_3_L1_4_Wij_nx252), .A0 (nx6725
          ), .A1 (CACHE_RST_dup_1490), .A2 (nx7139), .B0 (nx5485), .B1 (nx8785)
          ) ;
    oai32 CACHE_L0_3_L1_4_Wij_ix263 (.Y (CACHE_L0_3_L1_4_Wij_nx262), .A0 (nx6729
          ), .A1 (CACHE_RST_dup_1490), .A2 (nx7139), .B0 (nx5489), .B1 (nx8785)
          ) ;
    oai32 CACHE_L0_3_L1_4_Wij_ix273 (.Y (CACHE_L0_3_L1_4_Wij_nx272), .A0 (nx6733
          ), .A1 (CACHE_RST_dup_1490), .A2 (nx7143), .B0 (nx5493), .B1 (nx8785)
          ) ;
    inv01 ix7142 (.Y (nx7143), .A (CACHE_L0_3_L1_4_Wij_nx333)) ;
    oai32 CACHE_L0_3_L1_4_Wij_ix283 (.Y (CACHE_L0_3_L1_4_Wij_nx282), .A0 (nx6737
          ), .A1 (CACHE_RST_dup_1490), .A2 (nx7143), .B0 (nx5497), .B1 (nx8787)
          ) ;
    oai32 CACHE_L0_4_L1_0_Fij_ix213 (.Y (CACHE_L0_4_L1_0_Fij_nx212), .A0 (nx7145
          ), .A1 (nx8437), .A2 (nx7147), .B0 (nx5835), .B1 (nx8789)) ;
    inv01 ix7144 (.Y (nx7145), .A (MemDout[0])) ;
    inv02 ix7146 (.Y (nx7147), .A (CACHE_L0_4_L1_0_Fij_nx331)) ;
    oai32 CACHE_L0_4_L1_0_Fij_ix223 (.Y (CACHE_L0_4_L1_0_Fij_nx222), .A0 (nx7151
          ), .A1 (nx8437), .A2 (nx7147), .B0 (nx5837), .B1 (nx8789)) ;
    inv01 ix7150 (.Y (nx7151), .A (MemDout[1])) ;
    oai32 CACHE_L0_4_L1_0_Fij_ix233 (.Y (CACHE_L0_4_L1_0_Fij_nx232), .A0 (nx7153
          ), .A1 (nx8437), .A2 (nx7147), .B0 (nx5839), .B1 (nx8789)) ;
    inv01 ix7152 (.Y (nx7153), .A (MemDout[2])) ;
    oai32 CACHE_L0_4_L1_0_Fij_ix243 (.Y (CACHE_L0_4_L1_0_Fij_nx242), .A0 (nx7155
          ), .A1 (nx8437), .A2 (nx7147), .B0 (nx5841), .B1 (nx8789)) ;
    inv01 ix7154 (.Y (nx7155), .A (MemDout[3])) ;
    oai32 CACHE_L0_4_L1_0_Fij_ix253 (.Y (CACHE_L0_4_L1_0_Fij_nx252), .A0 (nx7157
          ), .A1 (nx8437), .A2 (nx7147), .B0 (nx5843), .B1 (nx8789)) ;
    inv01 ix7156 (.Y (nx7157), .A (MemDout[4])) ;
    oai32 CACHE_L0_4_L1_0_Fij_ix263 (.Y (CACHE_L0_4_L1_0_Fij_nx262), .A0 (nx7159
          ), .A1 (nx8439), .A2 (nx7147), .B0 (nx5845), .B1 (nx8789)) ;
    inv01 ix7158 (.Y (nx7159), .A (MemDout[5])) ;
    oai32 CACHE_L0_4_L1_0_Fij_ix273 (.Y (CACHE_L0_4_L1_0_Fij_nx272), .A0 (nx7161
          ), .A1 (nx8439), .A2 (nx7163), .B0 (nx5849), .B1 (nx8789)) ;
    inv01 ix7160 (.Y (nx7161), .A (MemDout[6])) ;
    inv01 ix7162 (.Y (nx7163), .A (CACHE_L0_4_L1_0_Fij_nx333)) ;
    oai32 CACHE_L0_4_L1_0_Fij_ix283 (.Y (CACHE_L0_4_L1_0_Fij_nx282), .A0 (nx7165
          ), .A1 (nx8439), .A2 (nx7163), .B0 (nx5851), .B1 (nx8791)) ;
    inv01 ix7164 (.Y (nx7165), .A (MemDout[7])) ;
    oai32 CACHE_L0_4_L1_0_Wij_ix213 (.Y (CACHE_L0_4_L1_0_Wij_nx212), .A0 (nx7145
          ), .A1 (nx8439), .A2 (nx7167), .B0 (nx5717), .B1 (nx8793)) ;
    inv02 ix7166 (.Y (nx7167), .A (CACHE_L0_4_L1_0_Wij_nx331)) ;
    oai32 CACHE_L0_4_L1_0_Wij_ix223 (.Y (CACHE_L0_4_L1_0_Wij_nx222), .A0 (nx7151
          ), .A1 (nx8439), .A2 (nx7167), .B0 (nx5721), .B1 (nx8793)) ;
    oai32 CACHE_L0_4_L1_0_Wij_ix233 (.Y (CACHE_L0_4_L1_0_Wij_nx232), .A0 (nx7153
          ), .A1 (nx8439), .A2 (nx7167), .B0 (nx5725), .B1 (nx8793)) ;
    oai32 CACHE_L0_4_L1_0_Wij_ix243 (.Y (CACHE_L0_4_L1_0_Wij_nx242), .A0 (nx7155
          ), .A1 (nx8439), .A2 (nx7167), .B0 (nx5729), .B1 (nx8793)) ;
    oai32 CACHE_L0_4_L1_0_Wij_ix253 (.Y (CACHE_L0_4_L1_0_Wij_nx252), .A0 (nx7157
          ), .A1 (CACHE_RST_dup_1512), .A2 (nx7167), .B0 (nx5733), .B1 (nx8793)
          ) ;
    oai32 CACHE_L0_4_L1_0_Wij_ix263 (.Y (CACHE_L0_4_L1_0_Wij_nx262), .A0 (nx7159
          ), .A1 (CACHE_RST_dup_1512), .A2 (nx7167), .B0 (nx5737), .B1 (nx8793)
          ) ;
    oai32 CACHE_L0_4_L1_0_Wij_ix273 (.Y (CACHE_L0_4_L1_0_Wij_nx272), .A0 (nx7161
          ), .A1 (CACHE_RST_dup_1512), .A2 (nx7171), .B0 (nx5741), .B1 (nx8793)
          ) ;
    inv01 ix7170 (.Y (nx7171), .A (CACHE_L0_4_L1_0_Wij_nx333)) ;
    oai32 CACHE_L0_4_L1_0_Wij_ix283 (.Y (CACHE_L0_4_L1_0_Wij_nx282), .A0 (nx7165
          ), .A1 (CACHE_RST_dup_1512), .A2 (nx7171), .B0 (nx5745), .B1 (nx8795)
          ) ;
    oai32 CACHE_L0_4_L1_1_Fij_ix213 (.Y (CACHE_L0_4_L1_1_Fij_nx212), .A0 (nx7173
          ), .A1 (nx8441), .A2 (nx7175), .B0 (nx6083), .B1 (nx8797)) ;
    inv01 ix7172 (.Y (nx7173), .A (MemDout[8])) ;
    inv02 ix7174 (.Y (nx7175), .A (CACHE_L0_4_L1_1_Fij_nx331)) ;
    oai32 CACHE_L0_4_L1_1_Fij_ix223 (.Y (CACHE_L0_4_L1_1_Fij_nx222), .A0 (nx7179
          ), .A1 (nx8441), .A2 (nx7175), .B0 (nx6085), .B1 (nx8797)) ;
    inv01 ix7178 (.Y (nx7179), .A (MemDout[9])) ;
    oai32 CACHE_L0_4_L1_1_Fij_ix233 (.Y (CACHE_L0_4_L1_1_Fij_nx232), .A0 (nx7181
          ), .A1 (nx8441), .A2 (nx7175), .B0 (nx6087), .B1 (nx8797)) ;
    inv01 ix7180 (.Y (nx7181), .A (MemDout[10])) ;
    oai32 CACHE_L0_4_L1_1_Fij_ix243 (.Y (CACHE_L0_4_L1_1_Fij_nx242), .A0 (nx7183
          ), .A1 (nx8441), .A2 (nx7175), .B0 (nx6089), .B1 (nx8797)) ;
    inv01 ix7182 (.Y (nx7183), .A (MemDout[11])) ;
    oai32 CACHE_L0_4_L1_1_Fij_ix253 (.Y (CACHE_L0_4_L1_1_Fij_nx252), .A0 (nx7185
          ), .A1 (nx8441), .A2 (nx7175), .B0 (nx6091), .B1 (nx8797)) ;
    inv01 ix7184 (.Y (nx7185), .A (MemDout[12])) ;
    oai32 CACHE_L0_4_L1_1_Fij_ix263 (.Y (CACHE_L0_4_L1_1_Fij_nx262), .A0 (nx7187
          ), .A1 (nx8443), .A2 (nx7175), .B0 (nx6093), .B1 (nx8797)) ;
    inv01 ix7186 (.Y (nx7187), .A (MemDout[13])) ;
    oai32 CACHE_L0_4_L1_1_Fij_ix273 (.Y (CACHE_L0_4_L1_1_Fij_nx272), .A0 (nx7189
          ), .A1 (nx8443), .A2 (nx7191), .B0 (nx6097), .B1 (nx8797)) ;
    inv01 ix7188 (.Y (nx7189), .A (MemDout[14])) ;
    inv01 ix7190 (.Y (nx7191), .A (CACHE_L0_4_L1_1_Fij_nx333)) ;
    oai32 CACHE_L0_4_L1_1_Fij_ix283 (.Y (CACHE_L0_4_L1_1_Fij_nx282), .A0 (nx7193
          ), .A1 (nx8443), .A2 (nx7191), .B0 (nx6099), .B1 (nx8799)) ;
    inv01 ix7192 (.Y (nx7193), .A (MemDout[15])) ;
    oai32 CACHE_L0_4_L1_1_Wij_ix213 (.Y (CACHE_L0_4_L1_1_Wij_nx212), .A0 (nx7173
          ), .A1 (nx8443), .A2 (nx7195), .B0 (nx5965), .B1 (nx8801)) ;
    inv02 ix7194 (.Y (nx7195), .A (CACHE_L0_4_L1_1_Wij_nx331)) ;
    oai32 CACHE_L0_4_L1_1_Wij_ix223 (.Y (CACHE_L0_4_L1_1_Wij_nx222), .A0 (nx7179
          ), .A1 (nx8443), .A2 (nx7195), .B0 (nx5969), .B1 (nx8801)) ;
    oai32 CACHE_L0_4_L1_1_Wij_ix233 (.Y (CACHE_L0_4_L1_1_Wij_nx232), .A0 (nx7181
          ), .A1 (nx8443), .A2 (nx7195), .B0 (nx5973), .B1 (nx8801)) ;
    oai32 CACHE_L0_4_L1_1_Wij_ix243 (.Y (CACHE_L0_4_L1_1_Wij_nx242), .A0 (nx7183
          ), .A1 (nx8443), .A2 (nx7195), .B0 (nx5977), .B1 (nx8801)) ;
    oai32 CACHE_L0_4_L1_1_Wij_ix253 (.Y (CACHE_L0_4_L1_1_Wij_nx252), .A0 (nx7185
          ), .A1 (CACHE_RST_dup_1534), .A2 (nx7195), .B0 (nx5981), .B1 (nx8801)
          ) ;
    oai32 CACHE_L0_4_L1_1_Wij_ix263 (.Y (CACHE_L0_4_L1_1_Wij_nx262), .A0 (nx7187
          ), .A1 (CACHE_RST_dup_1534), .A2 (nx7195), .B0 (nx5985), .B1 (nx8801)
          ) ;
    oai32 CACHE_L0_4_L1_1_Wij_ix273 (.Y (CACHE_L0_4_L1_1_Wij_nx272), .A0 (nx7189
          ), .A1 (CACHE_RST_dup_1534), .A2 (nx7199), .B0 (nx5989), .B1 (nx8801)
          ) ;
    inv01 ix7198 (.Y (nx7199), .A (CACHE_L0_4_L1_1_Wij_nx333)) ;
    oai32 CACHE_L0_4_L1_1_Wij_ix283 (.Y (CACHE_L0_4_L1_1_Wij_nx282), .A0 (nx7193
          ), .A1 (CACHE_RST_dup_1534), .A2 (nx7199), .B0 (nx5993), .B1 (nx8803)
          ) ;
    oai32 CACHE_L0_4_L1_2_Fij_ix213 (.Y (CACHE_L0_4_L1_2_Fij_nx212), .A0 (nx7201
          ), .A1 (nx8445), .A2 (nx7203), .B0 (nx6331), .B1 (nx8805)) ;
    inv01 ix7200 (.Y (nx7201), .A (MemDout[16])) ;
    inv02 ix7202 (.Y (nx7203), .A (CACHE_L0_4_L1_2_Fij_nx331)) ;
    oai32 CACHE_L0_4_L1_2_Fij_ix223 (.Y (CACHE_L0_4_L1_2_Fij_nx222), .A0 (nx7207
          ), .A1 (nx8445), .A2 (nx7203), .B0 (nx6333), .B1 (nx8805)) ;
    inv01 ix7206 (.Y (nx7207), .A (MemDout[17])) ;
    oai32 CACHE_L0_4_L1_2_Fij_ix233 (.Y (CACHE_L0_4_L1_2_Fij_nx232), .A0 (nx7209
          ), .A1 (nx8445), .A2 (nx7203), .B0 (nx6335), .B1 (nx8805)) ;
    inv01 ix7208 (.Y (nx7209), .A (MemDout[18])) ;
    oai32 CACHE_L0_4_L1_2_Fij_ix243 (.Y (CACHE_L0_4_L1_2_Fij_nx242), .A0 (nx7211
          ), .A1 (nx8445), .A2 (nx7203), .B0 (nx6337), .B1 (nx8805)) ;
    inv01 ix7210 (.Y (nx7211), .A (MemDout[19])) ;
    oai32 CACHE_L0_4_L1_2_Fij_ix253 (.Y (CACHE_L0_4_L1_2_Fij_nx252), .A0 (nx7213
          ), .A1 (nx8445), .A2 (nx7203), .B0 (nx6339), .B1 (nx8805)) ;
    inv01 ix7212 (.Y (nx7213), .A (MemDout[20])) ;
    oai32 CACHE_L0_4_L1_2_Fij_ix263 (.Y (CACHE_L0_4_L1_2_Fij_nx262), .A0 (nx7215
          ), .A1 (nx8447), .A2 (nx7203), .B0 (nx6341), .B1 (nx8805)) ;
    inv01 ix7214 (.Y (nx7215), .A (MemDout[21])) ;
    oai32 CACHE_L0_4_L1_2_Fij_ix273 (.Y (CACHE_L0_4_L1_2_Fij_nx272), .A0 (nx7217
          ), .A1 (nx8447), .A2 (nx7219), .B0 (nx6345), .B1 (nx8805)) ;
    inv01 ix7216 (.Y (nx7217), .A (MemDout[22])) ;
    inv01 ix7218 (.Y (nx7219), .A (CACHE_L0_4_L1_2_Fij_nx333)) ;
    oai32 CACHE_L0_4_L1_2_Fij_ix283 (.Y (CACHE_L0_4_L1_2_Fij_nx282), .A0 (nx7221
          ), .A1 (nx8447), .A2 (nx7219), .B0 (nx6347), .B1 (nx8807)) ;
    inv01 ix7220 (.Y (nx7221), .A (MemDout[23])) ;
    oai32 CACHE_L0_4_L1_2_Wij_ix213 (.Y (CACHE_L0_4_L1_2_Wij_nx212), .A0 (nx7201
          ), .A1 (nx8447), .A2 (nx7223), .B0 (nx6213), .B1 (nx8809)) ;
    inv02 ix7222 (.Y (nx7223), .A (CACHE_L0_4_L1_2_Wij_nx331)) ;
    oai32 CACHE_L0_4_L1_2_Wij_ix223 (.Y (CACHE_L0_4_L1_2_Wij_nx222), .A0 (nx7207
          ), .A1 (nx8447), .A2 (nx7223), .B0 (nx6217), .B1 (nx8809)) ;
    oai32 CACHE_L0_4_L1_2_Wij_ix233 (.Y (CACHE_L0_4_L1_2_Wij_nx232), .A0 (nx7209
          ), .A1 (nx8447), .A2 (nx7223), .B0 (nx6221), .B1 (nx8809)) ;
    oai32 CACHE_L0_4_L1_2_Wij_ix243 (.Y (CACHE_L0_4_L1_2_Wij_nx242), .A0 (nx7211
          ), .A1 (nx8447), .A2 (nx7223), .B0 (nx6225), .B1 (nx8809)) ;
    oai32 CACHE_L0_4_L1_2_Wij_ix253 (.Y (CACHE_L0_4_L1_2_Wij_nx252), .A0 (nx7213
          ), .A1 (CACHE_RST_dup_1556), .A2 (nx7223), .B0 (nx6229), .B1 (nx8809)
          ) ;
    oai32 CACHE_L0_4_L1_2_Wij_ix263 (.Y (CACHE_L0_4_L1_2_Wij_nx262), .A0 (nx7215
          ), .A1 (CACHE_RST_dup_1556), .A2 (nx7223), .B0 (nx6233), .B1 (nx8809)
          ) ;
    oai32 CACHE_L0_4_L1_2_Wij_ix273 (.Y (CACHE_L0_4_L1_2_Wij_nx272), .A0 (nx7217
          ), .A1 (CACHE_RST_dup_1556), .A2 (nx7227), .B0 (nx6237), .B1 (nx8809)
          ) ;
    inv01 ix7226 (.Y (nx7227), .A (CACHE_L0_4_L1_2_Wij_nx333)) ;
    oai32 CACHE_L0_4_L1_2_Wij_ix283 (.Y (CACHE_L0_4_L1_2_Wij_nx282), .A0 (nx7221
          ), .A1 (CACHE_RST_dup_1556), .A2 (nx7227), .B0 (nx6241), .B1 (nx8811)
          ) ;
    oai32 CACHE_L0_4_L1_3_Fij_ix213 (.Y (CACHE_L0_4_L1_3_Fij_nx212), .A0 (nx7229
          ), .A1 (nx8449), .A2 (nx7231), .B0 (nx6579), .B1 (nx8813)) ;
    inv01 ix7228 (.Y (nx7229), .A (MemDout[24])) ;
    inv02 ix7230 (.Y (nx7231), .A (CACHE_L0_4_L1_3_Fij_nx331)) ;
    oai32 CACHE_L0_4_L1_3_Fij_ix223 (.Y (CACHE_L0_4_L1_3_Fij_nx222), .A0 (nx7235
          ), .A1 (nx8449), .A2 (nx7231), .B0 (nx6581), .B1 (nx8813)) ;
    inv01 ix7234 (.Y (nx7235), .A (MemDout[25])) ;
    oai32 CACHE_L0_4_L1_3_Fij_ix233 (.Y (CACHE_L0_4_L1_3_Fij_nx232), .A0 (nx7237
          ), .A1 (nx8449), .A2 (nx7231), .B0 (nx6583), .B1 (nx8813)) ;
    inv01 ix7236 (.Y (nx7237), .A (MemDout[26])) ;
    oai32 CACHE_L0_4_L1_3_Fij_ix243 (.Y (CACHE_L0_4_L1_3_Fij_nx242), .A0 (nx7239
          ), .A1 (nx8449), .A2 (nx7231), .B0 (nx6585), .B1 (nx8813)) ;
    inv01 ix7238 (.Y (nx7239), .A (MemDout[27])) ;
    oai32 CACHE_L0_4_L1_3_Fij_ix253 (.Y (CACHE_L0_4_L1_3_Fij_nx252), .A0 (nx7241
          ), .A1 (nx8449), .A2 (nx7231), .B0 (nx6587), .B1 (nx8813)) ;
    inv01 ix7240 (.Y (nx7241), .A (MemDout[28])) ;
    oai32 CACHE_L0_4_L1_3_Fij_ix263 (.Y (CACHE_L0_4_L1_3_Fij_nx262), .A0 (nx7243
          ), .A1 (nx8451), .A2 (nx7231), .B0 (nx6589), .B1 (nx8813)) ;
    inv01 ix7242 (.Y (nx7243), .A (MemDout[29])) ;
    oai32 CACHE_L0_4_L1_3_Fij_ix273 (.Y (CACHE_L0_4_L1_3_Fij_nx272), .A0 (nx7245
          ), .A1 (nx8451), .A2 (nx7247), .B0 (nx6593), .B1 (nx8813)) ;
    inv01 ix7244 (.Y (nx7245), .A (MemDout[30])) ;
    inv01 ix7246 (.Y (nx7247), .A (CACHE_L0_4_L1_3_Fij_nx333)) ;
    oai32 CACHE_L0_4_L1_3_Fij_ix283 (.Y (CACHE_L0_4_L1_3_Fij_nx282), .A0 (nx7249
          ), .A1 (nx8451), .A2 (nx7247), .B0 (nx6595), .B1 (nx8815)) ;
    inv01 ix7248 (.Y (nx7249), .A (MemDout[31])) ;
    oai32 CACHE_L0_4_L1_3_Wij_ix213 (.Y (CACHE_L0_4_L1_3_Wij_nx212), .A0 (nx7229
          ), .A1 (nx8451), .A2 (nx7251), .B0 (nx6461), .B1 (nx8817)) ;
    inv02 ix7250 (.Y (nx7251), .A (CACHE_L0_4_L1_3_Wij_nx331)) ;
    oai32 CACHE_L0_4_L1_3_Wij_ix223 (.Y (CACHE_L0_4_L1_3_Wij_nx222), .A0 (nx7235
          ), .A1 (nx8451), .A2 (nx7251), .B0 (nx6465), .B1 (nx8817)) ;
    oai32 CACHE_L0_4_L1_3_Wij_ix233 (.Y (CACHE_L0_4_L1_3_Wij_nx232), .A0 (nx7237
          ), .A1 (nx8451), .A2 (nx7251), .B0 (nx6469), .B1 (nx8817)) ;
    oai32 CACHE_L0_4_L1_3_Wij_ix243 (.Y (CACHE_L0_4_L1_3_Wij_nx242), .A0 (nx7239
          ), .A1 (nx8451), .A2 (nx7251), .B0 (nx6473), .B1 (nx8817)) ;
    oai32 CACHE_L0_4_L1_3_Wij_ix253 (.Y (CACHE_L0_4_L1_3_Wij_nx252), .A0 (nx7241
          ), .A1 (CACHE_RST_dup_1578), .A2 (nx7251), .B0 (nx6477), .B1 (nx8817)
          ) ;
    oai32 CACHE_L0_4_L1_3_Wij_ix263 (.Y (CACHE_L0_4_L1_3_Wij_nx262), .A0 (nx7243
          ), .A1 (CACHE_RST_dup_1578), .A2 (nx7251), .B0 (nx6481), .B1 (nx8817)
          ) ;
    oai32 CACHE_L0_4_L1_3_Wij_ix273 (.Y (CACHE_L0_4_L1_3_Wij_nx272), .A0 (nx7245
          ), .A1 (CACHE_RST_dup_1578), .A2 (nx7255), .B0 (nx6485), .B1 (nx8817)
          ) ;
    inv01 ix7254 (.Y (nx7255), .A (CACHE_L0_4_L1_3_Wij_nx333)) ;
    oai32 CACHE_L0_4_L1_3_Wij_ix283 (.Y (CACHE_L0_4_L1_3_Wij_nx282), .A0 (nx7249
          ), .A1 (CACHE_RST_dup_1578), .A2 (nx7255), .B0 (nx6489), .B1 (nx8819)
          ) ;
    oai32 CACHE_L0_4_L1_4_Fij_ix213 (.Y (CACHE_L0_4_L1_4_Fij_nx212), .A0 (nx7257
          ), .A1 (nx8453), .A2 (nx7259), .B0 (nx6827), .B1 (nx8821)) ;
    inv01 ix7256 (.Y (nx7257), .A (MemDout[32])) ;
    inv02 ix7258 (.Y (nx7259), .A (CACHE_L0_4_L1_4_Fij_nx331)) ;
    oai32 CACHE_L0_4_L1_4_Fij_ix223 (.Y (CACHE_L0_4_L1_4_Fij_nx222), .A0 (nx7263
          ), .A1 (nx8453), .A2 (nx7259), .B0 (nx6829), .B1 (nx8821)) ;
    inv01 ix7262 (.Y (nx7263), .A (MemDout[33])) ;
    oai32 CACHE_L0_4_L1_4_Fij_ix233 (.Y (CACHE_L0_4_L1_4_Fij_nx232), .A0 (nx7265
          ), .A1 (nx8453), .A2 (nx7259), .B0 (nx6831), .B1 (nx8821)) ;
    inv01 ix7264 (.Y (nx7265), .A (MemDout[34])) ;
    oai32 CACHE_L0_4_L1_4_Fij_ix243 (.Y (CACHE_L0_4_L1_4_Fij_nx242), .A0 (nx7267
          ), .A1 (nx8453), .A2 (nx7259), .B0 (nx6833), .B1 (nx8821)) ;
    inv01 ix7266 (.Y (nx7267), .A (MemDout[35])) ;
    oai32 CACHE_L0_4_L1_4_Fij_ix253 (.Y (CACHE_L0_4_L1_4_Fij_nx252), .A0 (nx7269
          ), .A1 (nx8453), .A2 (nx7259), .B0 (nx6835), .B1 (nx8821)) ;
    inv01 ix7268 (.Y (nx7269), .A (MemDout[36])) ;
    oai32 CACHE_L0_4_L1_4_Fij_ix263 (.Y (CACHE_L0_4_L1_4_Fij_nx262), .A0 (nx7271
          ), .A1 (nx8455), .A2 (nx7259), .B0 (nx6837), .B1 (nx8821)) ;
    inv01 ix7270 (.Y (nx7271), .A (MemDout[37])) ;
    oai32 CACHE_L0_4_L1_4_Fij_ix273 (.Y (CACHE_L0_4_L1_4_Fij_nx272), .A0 (nx7273
          ), .A1 (nx8455), .A2 (nx7275), .B0 (nx6841), .B1 (nx8821)) ;
    inv01 ix7272 (.Y (nx7273), .A (MemDout[38])) ;
    inv01 ix7274 (.Y (nx7275), .A (CACHE_L0_4_L1_4_Fij_nx333)) ;
    oai32 CACHE_L0_4_L1_4_Fij_ix283 (.Y (CACHE_L0_4_L1_4_Fij_nx282), .A0 (nx7277
          ), .A1 (nx8455), .A2 (nx7275), .B0 (nx6843), .B1 (nx8823)) ;
    inv01 ix7276 (.Y (nx7277), .A (MemDout[39])) ;
    oai32 CACHE_L0_4_L1_4_Wij_ix213 (.Y (CACHE_L0_4_L1_4_Wij_nx212), .A0 (nx7257
          ), .A1 (nx8455), .A2 (nx7279), .B0 (nx6709), .B1 (nx8825)) ;
    inv02 ix7278 (.Y (nx7279), .A (CACHE_L0_4_L1_4_Wij_nx331)) ;
    oai32 CACHE_L0_4_L1_4_Wij_ix223 (.Y (CACHE_L0_4_L1_4_Wij_nx222), .A0 (nx7263
          ), .A1 (nx8455), .A2 (nx7279), .B0 (nx6713), .B1 (nx8825)) ;
    oai32 CACHE_L0_4_L1_4_Wij_ix233 (.Y (CACHE_L0_4_L1_4_Wij_nx232), .A0 (nx7265
          ), .A1 (nx8455), .A2 (nx7279), .B0 (nx6717), .B1 (nx8825)) ;
    oai32 CACHE_L0_4_L1_4_Wij_ix243 (.Y (CACHE_L0_4_L1_4_Wij_nx242), .A0 (nx7267
          ), .A1 (nx8455), .A2 (nx7279), .B0 (nx6721), .B1 (nx8825)) ;
    oai32 CACHE_L0_4_L1_4_Wij_ix253 (.Y (CACHE_L0_4_L1_4_Wij_nx252), .A0 (nx7269
          ), .A1 (CACHE_RST_dup_1600), .A2 (nx7279), .B0 (nx6725), .B1 (nx8825)
          ) ;
    oai32 CACHE_L0_4_L1_4_Wij_ix263 (.Y (CACHE_L0_4_L1_4_Wij_nx262), .A0 (nx7271
          ), .A1 (CACHE_RST_dup_1600), .A2 (nx7279), .B0 (nx6729), .B1 (nx8825)
          ) ;
    oai32 CACHE_L0_4_L1_4_Wij_ix273 (.Y (CACHE_L0_4_L1_4_Wij_nx272), .A0 (nx7273
          ), .A1 (CACHE_RST_dup_1600), .A2 (nx7283), .B0 (nx6733), .B1 (nx8825)
          ) ;
    inv01 ix7282 (.Y (nx7283), .A (CACHE_L0_4_L1_4_Wij_nx333)) ;
    oai32 CACHE_L0_4_L1_4_Wij_ix283 (.Y (CACHE_L0_4_L1_4_Wij_nx282), .A0 (nx7277
          ), .A1 (CACHE_RST_dup_1600), .A2 (nx7283), .B0 (nx6737), .B1 (nx8827)
          ) ;
    buf02 ix7284 (.Y (nx7285), .A (CONTROLLER_Restart)) ;
    inv01 ix7286 (.Y (nx7287), .A (CONTROLLER_CntRST)) ;
    inv02 ix7288 (.Y (nx7289), .A (nx7287)) ;
    inv02 ix7290 (.Y (nx7291), .A (nx7287)) ;
    inv02 ix7292 (.Y (nx7293), .A (nx7287)) ;
    inv02 CONTROLLER_ix810_rep_1 (.Y (nx7295), .A (CONTROLLER_nx124)) ;
    inv02 CONTROLLER_ix814_rep_1 (.Y (nx7297), .A (CONTROLLER_nx138)) ;
    inv02 ix7298 (.Y (nx7299), .A (nx8837)) ;
    inv02 ix7300 (.Y (nx7301), .A (nx8837)) ;
    inv02 CALCULATOR_ix1110_rep_1 (.Y (nx7303), .A (nx8837)) ;
    inv01 CALCULATOR_ix1110_rep_2 (.Y (nx7305), .A (nx8837)) ;
    inv02 ix7306 (.Y (nx7307), .A (nx8837)) ;
    inv02 ix7308 (.Y (nx7309), .A (nx8839)) ;
    inv02 ix7310 (.Y (nx7311), .A (nx8839)) ;
    inv02 ix7312 (.Y (nx7313), .A (nx8839)) ;
    inv01 ix7314 (.Y (nx7315), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_AddPToBoothOperand)) ;
    inv02 ix7316 (.Y (nx7317), .A (nx7315)) ;
    inv02 ix7318 (.Y (nx7319), .A (nx7315)) ;
    inv02 ix7320 (.Y (nx7321), .A (nx7315)) ;
    inv02 ix7322 (.Y (nx7323), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix7324 (.Y (nx7325), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix7326 (.Y (nx7327), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv01 ix7328 (.Y (nx7329), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx80)) ;
    inv02 ix7330 (.Y (nx7331), .A (nx7329)) ;
    inv02 ix7332 (.Y (nx7333), .A (nx7329)) ;
    inv02 ix7334 (.Y (nx7335), .A (nx7329)) ;
    inv02 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix565_rep_1 (.Y (
          nx7337), .A (RST)) ;
    inv02 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix565_rep_2 (.Y (
          nx7339), .A (RST)) ;
    inv02 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix565_rep_3 (.Y (
          nx7341), .A (RST)) ;
    inv02 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix565_rep_4 (.Y (
          nx7343), .A (RST)) ;
    inv02 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix565_rep_5 (.Y (
          nx7345), .A (RST)) ;
    inv02 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix565_rep_6 (.Y (
          nx7347), .A (RST)) ;
    inv02 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix565_rep_7 (.Y (
          nx7349), .A (RST)) ;
    inv02 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix565_rep_8 (.Y (
          nx7351), .A (RST)) ;
    inv02 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix565_rep_9 (.Y (
          nx7353), .A (RST)) ;
    inv02 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix565_rep_10 (.Y (
          nx7355), .A (RST)) ;
    inv02 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix565_rep_11 (.Y (
          nx7357), .A (RST)) ;
    inv02 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix565_rep_12 (.Y (
          nx7359), .A (RST)) ;
    inv02 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix565_rep_13 (.Y (
          nx7361), .A (RST)) ;
    inv02 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix565_rep_14 (.Y (
          nx7363), .A (RST)) ;
    inv02 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix565_rep_15 (.Y (
          nx7365), .A (RST)) ;
    inv02 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix565_rep_16 (.Y (
          nx7367), .A (RST)) ;
    inv02 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix565_rep_17 (.Y (
          nx7369), .A (RST)) ;
    inv02 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix565_rep_18 (.Y (
          nx7371), .A (RST)) ;
    inv02 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix565_rep_19 (.Y (
          nx7373), .A (RST)) ;
    inv02 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix565_rep_20 (.Y (
          nx7375), .A (RST)) ;
    inv02 CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix565_rep_21 (.Y (
          nx7377), .A (RST)) ;
    inv02 ix7378 (.Y (nx7379), .A (CALCULATOR_Start_dup_1144)) ;
    inv02 ix7380 (.Y (nx7381), .A (CALCULATOR_Start_dup_1144)) ;
    inv02 ix7382 (.Y (nx7383), .A (CALCULATOR_Start_dup_1144)) ;
    inv02 ix7384 (.Y (nx7385), .A (CALCULATOR_Start_dup_1144)) ;
    inv02 ix7386 (.Y (nx7387), .A (CALCULATOR_Start_dup_1144)) ;
    inv02 ix7388 (.Y (nx7389), .A (CALCULATOR_Start_dup_1144)) ;
    inv02 ix7390 (.Y (nx7391), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix7392 (.Y (nx7393), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix7394 (.Y (nx7395), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv01 ix7396 (.Y (nx7397), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_AddPToBoothOperand)) ;
    inv02 ix7398 (.Y (nx7399), .A (nx7397)) ;
    inv02 ix7400 (.Y (nx7401), .A (nx7397)) ;
    inv02 ix7402 (.Y (nx7403), .A (nx7397)) ;
    inv02 ix7404 (.Y (nx7405), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix7406 (.Y (nx7407), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix7408 (.Y (nx7409), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv01 ix7410 (.Y (nx7411), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx80)) ;
    inv02 ix7412 (.Y (nx7413), .A (nx7411)) ;
    inv02 ix7414 (.Y (nx7415), .A (nx7411)) ;
    inv02 ix7416 (.Y (nx7417), .A (nx7411)) ;
    inv02 ix7418 (.Y (nx7419), .A (CALCULATOR_Start_dup_1149)) ;
    inv02 ix7420 (.Y (nx7421), .A (CALCULATOR_Start_dup_1149)) ;
    inv02 ix7422 (.Y (nx7423), .A (CALCULATOR_Start_dup_1149)) ;
    inv02 ix7424 (.Y (nx7425), .A (CALCULATOR_Start_dup_1149)) ;
    inv02 ix7426 (.Y (nx7427), .A (CALCULATOR_Start_dup_1149)) ;
    inv02 ix7428 (.Y (nx7429), .A (CALCULATOR_Start_dup_1149)) ;
    inv02 ix7430 (.Y (nx7431), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix7432 (.Y (nx7433), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix7434 (.Y (nx7435), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv01 ix7436 (.Y (nx7437), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_AddPToBoothOperand)) ;
    inv02 ix7438 (.Y (nx7439), .A (nx7437)) ;
    inv02 ix7440 (.Y (nx7441), .A (nx7437)) ;
    inv02 ix7442 (.Y (nx7443), .A (nx7437)) ;
    inv02 ix7444 (.Y (nx7445), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix7446 (.Y (nx7447), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix7448 (.Y (nx7449), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv01 ix7450 (.Y (nx7451), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx80)) ;
    inv02 ix7452 (.Y (nx7453), .A (nx7451)) ;
    inv02 ix7454 (.Y (nx7455), .A (nx7451)) ;
    inv02 ix7456 (.Y (nx7457), .A (nx7451)) ;
    inv02 ix7458 (.Y (nx7459), .A (CALCULATOR_Start_dup_1154)) ;
    inv02 ix7460 (.Y (nx7461), .A (CALCULATOR_Start_dup_1154)) ;
    inv02 ix7462 (.Y (nx7463), .A (CALCULATOR_Start_dup_1154)) ;
    inv02 ix7464 (.Y (nx7465), .A (CALCULATOR_Start_dup_1154)) ;
    inv02 ix7466 (.Y (nx7467), .A (CALCULATOR_Start_dup_1154)) ;
    inv02 ix7468 (.Y (nx7469), .A (CALCULATOR_Start_dup_1154)) ;
    inv02 ix7470 (.Y (nx7471), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix7472 (.Y (nx7473), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix7474 (.Y (nx7475), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv01 ix7476 (.Y (nx7477), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_AddPToBoothOperand)) ;
    inv02 ix7478 (.Y (nx7479), .A (nx7477)) ;
    inv02 ix7480 (.Y (nx7481), .A (nx7477)) ;
    inv02 ix7482 (.Y (nx7483), .A (nx7477)) ;
    inv02 ix7484 (.Y (nx7485), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix7486 (.Y (nx7487), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix7488 (.Y (nx7489), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv01 ix7490 (.Y (nx7491), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx80)) ;
    inv02 ix7492 (.Y (nx7493), .A (nx7491)) ;
    inv02 ix7494 (.Y (nx7495), .A (nx7491)) ;
    inv02 ix7496 (.Y (nx7497), .A (nx7491)) ;
    inv02 ix7498 (.Y (nx7499), .A (CALCULATOR_Start_dup_1159)) ;
    inv02 ix7500 (.Y (nx7501), .A (CALCULATOR_Start_dup_1159)) ;
    inv02 ix7502 (.Y (nx7503), .A (CALCULATOR_Start_dup_1159)) ;
    inv02 ix7504 (.Y (nx7505), .A (CALCULATOR_Start_dup_1159)) ;
    inv02 ix7506 (.Y (nx7507), .A (CALCULATOR_Start_dup_1159)) ;
    inv02 ix7508 (.Y (nx7509), .A (CALCULATOR_Start_dup_1159)) ;
    inv02 ix7510 (.Y (nx7511), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix7512 (.Y (nx7513), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix7514 (.Y (nx7515), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv01 ix7516 (.Y (nx7517), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_AddPToBoothOperand)) ;
    inv02 ix7518 (.Y (nx7519), .A (nx7517)) ;
    inv02 ix7520 (.Y (nx7521), .A (nx7517)) ;
    inv02 ix7522 (.Y (nx7523), .A (nx7517)) ;
    inv02 ix7524 (.Y (nx7525), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix7526 (.Y (nx7527), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix7528 (.Y (nx7529), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv01 ix7530 (.Y (nx7531), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx80)) ;
    inv02 ix7532 (.Y (nx7533), .A (nx7531)) ;
    inv02 ix7534 (.Y (nx7535), .A (nx7531)) ;
    inv02 ix7536 (.Y (nx7537), .A (nx7531)) ;
    inv02 ix7538 (.Y (nx7539), .A (CALCULATOR_Start_dup_1164)) ;
    inv02 ix7540 (.Y (nx7541), .A (CALCULATOR_Start_dup_1164)) ;
    inv02 ix7542 (.Y (nx7543), .A (CALCULATOR_Start_dup_1164)) ;
    inv02 ix7544 (.Y (nx7545), .A (CALCULATOR_Start_dup_1164)) ;
    inv02 ix7546 (.Y (nx7547), .A (CALCULATOR_Start_dup_1164)) ;
    inv02 ix7548 (.Y (nx7549), .A (CALCULATOR_Start_dup_1164)) ;
    inv02 ix7550 (.Y (nx7551), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix7552 (.Y (nx7553), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix7554 (.Y (nx7555), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv01 ix7556 (.Y (nx7557), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_AddPToBoothOperand)) ;
    inv02 ix7558 (.Y (nx7559), .A (nx7557)) ;
    inv02 ix7560 (.Y (nx7561), .A (nx7557)) ;
    inv02 ix7562 (.Y (nx7563), .A (nx7557)) ;
    inv02 ix7564 (.Y (nx7565), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix7566 (.Y (nx7567), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix7568 (.Y (nx7569), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv01 ix7570 (.Y (nx7571), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx80)) ;
    inv02 ix7572 (.Y (nx7573), .A (nx7571)) ;
    inv02 ix7574 (.Y (nx7575), .A (nx7571)) ;
    inv02 ix7576 (.Y (nx7577), .A (nx7571)) ;
    inv02 ix7578 (.Y (nx7579), .A (CALCULATOR_Start_dup_1169)) ;
    inv02 ix7580 (.Y (nx7581), .A (CALCULATOR_Start_dup_1169)) ;
    inv02 ix7582 (.Y (nx7583), .A (CALCULATOR_Start_dup_1169)) ;
    inv02 ix7584 (.Y (nx7585), .A (CALCULATOR_Start_dup_1169)) ;
    inv02 ix7586 (.Y (nx7587), .A (CALCULATOR_Start_dup_1169)) ;
    inv02 ix7588 (.Y (nx7589), .A (CALCULATOR_Start_dup_1169)) ;
    inv02 ix7590 (.Y (nx7591), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix7592 (.Y (nx7593), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix7594 (.Y (nx7595), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv01 ix7596 (.Y (nx7597), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_AddPToBoothOperand)) ;
    inv02 ix7598 (.Y (nx7599), .A (nx7597)) ;
    inv02 ix7600 (.Y (nx7601), .A (nx7597)) ;
    inv02 ix7602 (.Y (nx7603), .A (nx7597)) ;
    inv02 ix7604 (.Y (nx7605), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix7606 (.Y (nx7607), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix7608 (.Y (nx7609), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv01 ix7610 (.Y (nx7611), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx80)) ;
    inv02 ix7612 (.Y (nx7613), .A (nx7611)) ;
    inv02 ix7614 (.Y (nx7615), .A (nx7611)) ;
    inv02 ix7616 (.Y (nx7617), .A (nx7611)) ;
    inv02 ix7618 (.Y (nx7619), .A (CALCULATOR_Start_dup_1174)) ;
    inv02 ix7620 (.Y (nx7621), .A (CALCULATOR_Start_dup_1174)) ;
    inv02 ix7622 (.Y (nx7623), .A (CALCULATOR_Start_dup_1174)) ;
    inv02 ix7624 (.Y (nx7625), .A (CALCULATOR_Start_dup_1174)) ;
    inv02 ix7626 (.Y (nx7627), .A (CALCULATOR_Start_dup_1174)) ;
    inv02 ix7628 (.Y (nx7629), .A (CALCULATOR_Start_dup_1174)) ;
    inv02 ix7630 (.Y (nx7631), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix7632 (.Y (nx7633), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix7634 (.Y (nx7635), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv01 ix7636 (.Y (nx7637), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_AddPToBoothOperand)) ;
    inv02 ix7638 (.Y (nx7639), .A (nx7637)) ;
    inv02 ix7640 (.Y (nx7641), .A (nx7637)) ;
    inv02 ix7642 (.Y (nx7643), .A (nx7637)) ;
    inv02 ix7644 (.Y (nx7645), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix7646 (.Y (nx7647), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix7648 (.Y (nx7649), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv01 ix7650 (.Y (nx7651), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx80)) ;
    inv02 ix7652 (.Y (nx7653), .A (nx7651)) ;
    inv02 ix7654 (.Y (nx7655), .A (nx7651)) ;
    inv02 ix7656 (.Y (nx7657), .A (nx7651)) ;
    inv02 ix7658 (.Y (nx7659), .A (CALCULATOR_Start_dup_1179)) ;
    inv02 ix7660 (.Y (nx7661), .A (CALCULATOR_Start_dup_1179)) ;
    inv02 ix7662 (.Y (nx7663), .A (CALCULATOR_Start_dup_1179)) ;
    inv02 ix7664 (.Y (nx7665), .A (CALCULATOR_Start_dup_1179)) ;
    inv02 ix7666 (.Y (nx7667), .A (CALCULATOR_Start_dup_1179)) ;
    inv02 ix7668 (.Y (nx7669), .A (CALCULATOR_Start_dup_1179)) ;
    inv02 ix7670 (.Y (nx7671), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix7672 (.Y (nx7673), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix7674 (.Y (nx7675), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv01 ix7676 (.Y (nx7677), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_AddPToBoothOperand)) ;
    inv02 ix7678 (.Y (nx7679), .A (nx7677)) ;
    inv02 ix7680 (.Y (nx7681), .A (nx7677)) ;
    inv02 ix7682 (.Y (nx7683), .A (nx7677)) ;
    inv02 ix7684 (.Y (nx7685), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix7686 (.Y (nx7687), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix7688 (.Y (nx7689), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv01 ix7690 (.Y (nx7691), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx80)) ;
    inv02 ix7692 (.Y (nx7693), .A (nx7691)) ;
    inv02 ix7694 (.Y (nx7695), .A (nx7691)) ;
    inv02 ix7696 (.Y (nx7697), .A (nx7691)) ;
    inv02 ix7698 (.Y (nx7699), .A (CALCULATOR_Start_dup_1184)) ;
    inv02 ix7700 (.Y (nx7701), .A (CALCULATOR_Start_dup_1184)) ;
    inv02 ix7702 (.Y (nx7703), .A (CALCULATOR_Start_dup_1184)) ;
    inv02 ix7704 (.Y (nx7705), .A (CALCULATOR_Start_dup_1184)) ;
    inv02 ix7706 (.Y (nx7707), .A (CALCULATOR_Start_dup_1184)) ;
    inv02 ix7708 (.Y (nx7709), .A (CALCULATOR_Start_dup_1184)) ;
    inv02 ix7710 (.Y (nx7711), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix7712 (.Y (nx7713), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix7714 (.Y (nx7715), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv01 ix7716 (.Y (nx7717), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_AddPToBoothOperand)) ;
    inv02 ix7718 (.Y (nx7719), .A (nx7717)) ;
    inv02 ix7720 (.Y (nx7721), .A (nx7717)) ;
    inv02 ix7722 (.Y (nx7723), .A (nx7717)) ;
    inv02 ix7724 (.Y (nx7725), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix7726 (.Y (nx7727), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix7728 (.Y (nx7729), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv01 ix7730 (.Y (nx7731), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx80)) ;
    inv02 ix7732 (.Y (nx7733), .A (nx7731)) ;
    inv02 ix7734 (.Y (nx7735), .A (nx7731)) ;
    inv02 ix7736 (.Y (nx7737), .A (nx7731)) ;
    inv02 ix7738 (.Y (nx7739), .A (CALCULATOR_Start_dup_1189)) ;
    inv02 ix7740 (.Y (nx7741), .A (CALCULATOR_Start_dup_1189)) ;
    inv02 ix7742 (.Y (nx7743), .A (CALCULATOR_Start_dup_1189)) ;
    inv02 ix7744 (.Y (nx7745), .A (CALCULATOR_Start_dup_1189)) ;
    inv02 ix7746 (.Y (nx7747), .A (CALCULATOR_Start_dup_1189)) ;
    inv02 ix7748 (.Y (nx7749), .A (CALCULATOR_Start_dup_1189)) ;
    inv02 ix7750 (.Y (nx7751), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix7752 (.Y (nx7753), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix7754 (.Y (nx7755), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv01 ix7756 (.Y (nx7757), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_AddPToBoothOperand)) ;
    inv02 ix7758 (.Y (nx7759), .A (nx7757)) ;
    inv02 ix7760 (.Y (nx7761), .A (nx7757)) ;
    inv02 ix7762 (.Y (nx7763), .A (nx7757)) ;
    inv02 ix7764 (.Y (nx7765), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix7766 (.Y (nx7767), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix7768 (.Y (nx7769), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv01 ix7770 (.Y (nx7771), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx80)) ;
    inv02 ix7772 (.Y (nx7773), .A (nx7771)) ;
    inv02 ix7774 (.Y (nx7775), .A (nx7771)) ;
    inv02 ix7776 (.Y (nx7777), .A (nx7771)) ;
    inv02 ix7778 (.Y (nx7779), .A (CALCULATOR_Start_dup_1194)) ;
    inv02 ix7780 (.Y (nx7781), .A (CALCULATOR_Start_dup_1194)) ;
    inv02 ix7782 (.Y (nx7783), .A (CALCULATOR_Start_dup_1194)) ;
    inv02 ix7784 (.Y (nx7785), .A (CALCULATOR_Start_dup_1194)) ;
    inv02 ix7786 (.Y (nx7787), .A (CALCULATOR_Start_dup_1194)) ;
    inv02 ix7788 (.Y (nx7789), .A (CALCULATOR_Start_dup_1194)) ;
    inv02 ix7790 (.Y (nx7791), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix7792 (.Y (nx7793), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix7794 (.Y (nx7795), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv01 ix7796 (.Y (nx7797), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_AddPToBoothOperand)) ;
    inv02 ix7798 (.Y (nx7799), .A (nx7797)) ;
    inv02 ix7800 (.Y (nx7801), .A (nx7797)) ;
    inv02 ix7802 (.Y (nx7803), .A (nx7797)) ;
    inv02 ix7804 (.Y (nx7805), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix7806 (.Y (nx7807), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix7808 (.Y (nx7809), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv01 ix7810 (.Y (nx7811), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx80)) ;
    inv02 ix7812 (.Y (nx7813), .A (nx7811)) ;
    inv02 ix7814 (.Y (nx7815), .A (nx7811)) ;
    inv02 ix7816 (.Y (nx7817), .A (nx7811)) ;
    inv02 ix7818 (.Y (nx7819), .A (CALCULATOR_Start_dup_1199)) ;
    inv02 ix7820 (.Y (nx7821), .A (CALCULATOR_Start_dup_1199)) ;
    inv02 ix7822 (.Y (nx7823), .A (CALCULATOR_Start_dup_1199)) ;
    inv02 ix7824 (.Y (nx7825), .A (CALCULATOR_Start_dup_1199)) ;
    inv02 ix7826 (.Y (nx7827), .A (CALCULATOR_Start_dup_1199)) ;
    inv02 ix7828 (.Y (nx7829), .A (CALCULATOR_Start_dup_1199)) ;
    inv02 ix7830 (.Y (nx7831), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix7832 (.Y (nx7833), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix7834 (.Y (nx7835), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv01 ix7836 (.Y (nx7837), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_AddPToBoothOperand)) ;
    inv02 ix7838 (.Y (nx7839), .A (nx7837)) ;
    inv02 ix7840 (.Y (nx7841), .A (nx7837)) ;
    inv02 ix7842 (.Y (nx7843), .A (nx7837)) ;
    inv02 ix7844 (.Y (nx7845), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix7846 (.Y (nx7847), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix7848 (.Y (nx7849), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv01 ix7850 (.Y (nx7851), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx80)) ;
    inv02 ix7852 (.Y (nx7853), .A (nx7851)) ;
    inv02 ix7854 (.Y (nx7855), .A (nx7851)) ;
    inv02 ix7856 (.Y (nx7857), .A (nx7851)) ;
    inv02 ix7858 (.Y (nx7859), .A (CALCULATOR_Start_dup_1204)) ;
    inv02 ix7860 (.Y (nx7861), .A (CALCULATOR_Start_dup_1204)) ;
    inv02 ix7862 (.Y (nx7863), .A (CALCULATOR_Start_dup_1204)) ;
    inv02 ix7864 (.Y (nx7865), .A (CALCULATOR_Start_dup_1204)) ;
    inv02 ix7866 (.Y (nx7867), .A (CALCULATOR_Start_dup_1204)) ;
    inv02 ix7868 (.Y (nx7869), .A (CALCULATOR_Start_dup_1204)) ;
    inv02 ix7870 (.Y (nx7871), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix7872 (.Y (nx7873), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix7874 (.Y (nx7875), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv01 ix7876 (.Y (nx7877), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_AddPToBoothOperand)) ;
    inv02 ix7878 (.Y (nx7879), .A (nx7877)) ;
    inv02 ix7880 (.Y (nx7881), .A (nx7877)) ;
    inv02 ix7882 (.Y (nx7883), .A (nx7877)) ;
    inv02 ix7884 (.Y (nx7885), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix7886 (.Y (nx7887), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix7888 (.Y (nx7889), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv01 ix7890 (.Y (nx7891), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx80)) ;
    inv02 ix7892 (.Y (nx7893), .A (nx7891)) ;
    inv02 ix7894 (.Y (nx7895), .A (nx7891)) ;
    inv02 ix7896 (.Y (nx7897), .A (nx7891)) ;
    inv02 ix7898 (.Y (nx7899), .A (CALCULATOR_Start_dup_1209)) ;
    inv02 ix7900 (.Y (nx7901), .A (CALCULATOR_Start_dup_1209)) ;
    inv02 ix7902 (.Y (nx7903), .A (CALCULATOR_Start_dup_1209)) ;
    inv02 ix7904 (.Y (nx7905), .A (CALCULATOR_Start_dup_1209)) ;
    inv02 ix7906 (.Y (nx7907), .A (CALCULATOR_Start_dup_1209)) ;
    inv02 ix7908 (.Y (nx7909), .A (CALCULATOR_Start_dup_1209)) ;
    inv02 ix7910 (.Y (nx7911), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix7912 (.Y (nx7913), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix7914 (.Y (nx7915), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv01 ix7916 (.Y (nx7917), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_AddPToBoothOperand)) ;
    inv02 ix7918 (.Y (nx7919), .A (nx7917)) ;
    inv02 ix7920 (.Y (nx7921), .A (nx7917)) ;
    inv02 ix7922 (.Y (nx7923), .A (nx7917)) ;
    inv02 ix7924 (.Y (nx7925), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix7926 (.Y (nx7927), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix7928 (.Y (nx7929), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv01 ix7930 (.Y (nx7931), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_nx80)) ;
    inv02 ix7932 (.Y (nx7933), .A (nx7931)) ;
    inv02 ix7934 (.Y (nx7935), .A (nx7931)) ;
    inv02 ix7936 (.Y (nx7937), .A (nx7931)) ;
    inv02 ix7938 (.Y (nx7939), .A (CALCULATOR_Start_dup_1222)) ;
    inv02 ix7940 (.Y (nx7941), .A (CALCULATOR_Start_dup_1222)) ;
    inv02 ix7942 (.Y (nx7943), .A (CALCULATOR_Start_dup_1222)) ;
    inv02 ix7944 (.Y (nx7945), .A (CALCULATOR_Start_dup_1222)) ;
    inv02 ix7946 (.Y (nx7947), .A (CALCULATOR_Start_dup_1222)) ;
    inv02 ix7948 (.Y (nx7949), .A (CALCULATOR_Start_dup_1222)) ;
    inv02 ix7950 (.Y (nx7951), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix7952 (.Y (nx7953), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix7954 (.Y (nx7955), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv01 ix7956 (.Y (nx7957), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_AddPToBoothOperand)) ;
    inv02 ix7958 (.Y (nx7959), .A (nx7957)) ;
    inv02 ix7960 (.Y (nx7961), .A (nx7957)) ;
    inv02 ix7962 (.Y (nx7963), .A (nx7957)) ;
    inv02 ix7964 (.Y (nx7965), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix7966 (.Y (nx7967), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix7968 (.Y (nx7969), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv01 ix7970 (.Y (nx7971), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_nx80)) ;
    inv02 ix7972 (.Y (nx7973), .A (nx7971)) ;
    inv02 ix7974 (.Y (nx7975), .A (nx7971)) ;
    inv02 ix7976 (.Y (nx7977), .A (nx7971)) ;
    inv02 ix7978 (.Y (nx7979), .A (CALCULATOR_Start_dup_1235)) ;
    inv02 ix7980 (.Y (nx7981), .A (CALCULATOR_Start_dup_1235)) ;
    inv02 ix7982 (.Y (nx7983), .A (CALCULATOR_Start_dup_1235)) ;
    inv02 ix7984 (.Y (nx7985), .A (CALCULATOR_Start_dup_1235)) ;
    inv02 ix7986 (.Y (nx7987), .A (CALCULATOR_Start_dup_1235)) ;
    inv02 ix7988 (.Y (nx7989), .A (CALCULATOR_Start_dup_1235)) ;
    inv02 ix7990 (.Y (nx7991), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix7992 (.Y (nx7993), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix7994 (.Y (nx7995), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv01 ix7996 (.Y (nx7997), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_AddPToBoothOperand)) ;
    inv02 ix7998 (.Y (nx7999), .A (nx7997)) ;
    inv02 ix8000 (.Y (nx8001), .A (nx7997)) ;
    inv02 ix8002 (.Y (nx8003), .A (nx7997)) ;
    inv02 ix8004 (.Y (nx8005), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix8006 (.Y (nx8007), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix8008 (.Y (nx8009), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv01 ix8010 (.Y (nx8011), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_nx80)) ;
    inv02 ix8012 (.Y (nx8013), .A (nx8011)) ;
    inv02 ix8014 (.Y (nx8015), .A (nx8011)) ;
    inv02 ix8016 (.Y (nx8017), .A (nx8011)) ;
    inv02 ix8018 (.Y (nx8019), .A (CALCULATOR_Start_dup_1248)) ;
    inv02 ix8020 (.Y (nx8021), .A (CALCULATOR_Start_dup_1248)) ;
    inv02 ix8022 (.Y (nx8023), .A (CALCULATOR_Start_dup_1248)) ;
    inv02 ix8024 (.Y (nx8025), .A (CALCULATOR_Start_dup_1248)) ;
    inv02 ix8026 (.Y (nx8027), .A (CALCULATOR_Start_dup_1248)) ;
    inv02 ix8028 (.Y (nx8029), .A (CALCULATOR_Start_dup_1248)) ;
    inv02 ix8030 (.Y (nx8031), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix8032 (.Y (nx8033), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix8034 (.Y (nx8035), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv01 ix8036 (.Y (nx8037), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_AddPToBoothOperand)) ;
    inv02 ix8038 (.Y (nx8039), .A (nx8037)) ;
    inv02 ix8040 (.Y (nx8041), .A (nx8037)) ;
    inv02 ix8042 (.Y (nx8043), .A (nx8037)) ;
    inv02 ix8044 (.Y (nx8045), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix8046 (.Y (nx8047), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix8048 (.Y (nx8049), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv01 ix8050 (.Y (nx8051), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_nx80)) ;
    inv02 ix8052 (.Y (nx8053), .A (nx8051)) ;
    inv02 ix8054 (.Y (nx8055), .A (nx8051)) ;
    inv02 ix8056 (.Y (nx8057), .A (nx8051)) ;
    inv02 ix8058 (.Y (nx8059), .A (CALCULATOR_Start_dup_1261)) ;
    inv02 ix8060 (.Y (nx8061), .A (CALCULATOR_Start_dup_1261)) ;
    inv02 ix8062 (.Y (nx8063), .A (CALCULATOR_Start_dup_1261)) ;
    inv02 ix8064 (.Y (nx8065), .A (CALCULATOR_Start_dup_1261)) ;
    inv02 ix8066 (.Y (nx8067), .A (CALCULATOR_Start_dup_1261)) ;
    inv02 ix8068 (.Y (nx8069), .A (CALCULATOR_Start_dup_1261)) ;
    inv02 ix8070 (.Y (nx8071), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix8072 (.Y (nx8073), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix8074 (.Y (nx8075), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv01 ix8076 (.Y (nx8077), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_AddPToBoothOperand)) ;
    inv02 ix8078 (.Y (nx8079), .A (nx8077)) ;
    inv02 ix8080 (.Y (nx8081), .A (nx8077)) ;
    inv02 ix8082 (.Y (nx8083), .A (nx8077)) ;
    inv02 ix8084 (.Y (nx8085), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix8086 (.Y (nx8087), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix8088 (.Y (nx8089), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv01 ix8090 (.Y (nx8091), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx80)) ;
    inv02 ix8092 (.Y (nx8093), .A (nx8091)) ;
    inv02 ix8094 (.Y (nx8095), .A (nx8091)) ;
    inv02 ix8096 (.Y (nx8097), .A (nx8091)) ;
    inv02 ix8098 (.Y (nx8099), .A (CALCULATOR_Start_dup_1274)) ;
    inv02 ix8100 (.Y (nx8101), .A (CALCULATOR_Start_dup_1274)) ;
    inv02 ix8102 (.Y (nx8103), .A (CALCULATOR_Start_dup_1274)) ;
    inv02 ix8104 (.Y (nx8105), .A (CALCULATOR_Start_dup_1274)) ;
    inv02 ix8106 (.Y (nx8107), .A (CALCULATOR_Start_dup_1274)) ;
    inv02 ix8108 (.Y (nx8109), .A (CALCULATOR_Start_dup_1274)) ;
    inv02 ix8110 (.Y (nx8111), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix8112 (.Y (nx8113), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix8114 (.Y (nx8115), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv01 ix8116 (.Y (nx8117), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_AddPToBoothOperand)) ;
    inv02 ix8118 (.Y (nx8119), .A (nx8117)) ;
    inv02 ix8120 (.Y (nx8121), .A (nx8117)) ;
    inv02 ix8122 (.Y (nx8123), .A (nx8117)) ;
    inv02 ix8124 (.Y (nx8125), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix8126 (.Y (nx8127), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix8128 (.Y (nx8129), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv01 ix8130 (.Y (nx8131), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_nx80)) ;
    inv02 ix8132 (.Y (nx8133), .A (nx8131)) ;
    inv02 ix8134 (.Y (nx8135), .A (nx8131)) ;
    inv02 ix8136 (.Y (nx8137), .A (nx8131)) ;
    inv02 ix8138 (.Y (nx8139), .A (CALCULATOR_Start_dup_1287)) ;
    inv02 ix8140 (.Y (nx8141), .A (CALCULATOR_Start_dup_1287)) ;
    inv02 ix8142 (.Y (nx8143), .A (CALCULATOR_Start_dup_1287)) ;
    inv02 ix8144 (.Y (nx8145), .A (CALCULATOR_Start_dup_1287)) ;
    inv02 ix8146 (.Y (nx8147), .A (CALCULATOR_Start_dup_1287)) ;
    inv02 ix8148 (.Y (nx8149), .A (CALCULATOR_Start_dup_1287)) ;
    inv02 ix8150 (.Y (nx8151), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix8152 (.Y (nx8153), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix8154 (.Y (nx8155), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv01 ix8156 (.Y (nx8157), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_AddPToBoothOperand)) ;
    inv02 ix8158 (.Y (nx8159), .A (nx8157)) ;
    inv02 ix8160 (.Y (nx8161), .A (nx8157)) ;
    inv02 ix8162 (.Y (nx8163), .A (nx8157)) ;
    inv02 ix8164 (.Y (nx8165), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix8166 (.Y (nx8167), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix8168 (.Y (nx8169), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv01 ix8170 (.Y (nx8171), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_nx80)) ;
    inv02 ix8172 (.Y (nx8173), .A (nx8171)) ;
    inv02 ix8174 (.Y (nx8175), .A (nx8171)) ;
    inv02 ix8176 (.Y (nx8177), .A (nx8171)) ;
    inv02 ix8178 (.Y (nx8179), .A (CALCULATOR_Start_dup_1300)) ;
    inv02 ix8180 (.Y (nx8181), .A (CALCULATOR_Start_dup_1300)) ;
    inv02 ix8182 (.Y (nx8183), .A (CALCULATOR_Start_dup_1300)) ;
    inv02 ix8184 (.Y (nx8185), .A (CALCULATOR_Start_dup_1300)) ;
    inv02 ix8186 (.Y (nx8187), .A (CALCULATOR_Start_dup_1300)) ;
    inv02 ix8188 (.Y (nx8189), .A (CALCULATOR_Start_dup_1300)) ;
    inv02 ix8190 (.Y (nx8191), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix8192 (.Y (nx8193), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix8194 (.Y (nx8195), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv01 ix8196 (.Y (nx8197), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_AddPToBoothOperand)) ;
    inv02 ix8198 (.Y (nx8199), .A (nx8197)) ;
    inv02 ix8200 (.Y (nx8201), .A (nx8197)) ;
    inv02 ix8202 (.Y (nx8203), .A (nx8197)) ;
    inv02 ix8204 (.Y (nx8205), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix8206 (.Y (nx8207), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix8208 (.Y (nx8209), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv01 ix8210 (.Y (nx8211), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_nx80)) ;
    inv02 ix8212 (.Y (nx8213), .A (nx8211)) ;
    inv02 ix8214 (.Y (nx8215), .A (nx8211)) ;
    inv02 ix8216 (.Y (nx8217), .A (nx8211)) ;
    inv02 ix8218 (.Y (nx8219), .A (CALCULATOR_Start_dup_1313)) ;
    inv02 ix8220 (.Y (nx8221), .A (CALCULATOR_Start_dup_1313)) ;
    inv02 ix8222 (.Y (nx8223), .A (CALCULATOR_Start_dup_1313)) ;
    inv02 ix8224 (.Y (nx8225), .A (CALCULATOR_Start_dup_1313)) ;
    inv02 ix8226 (.Y (nx8227), .A (CALCULATOR_Start_dup_1313)) ;
    inv02 ix8228 (.Y (nx8229), .A (CALCULATOR_Start_dup_1313)) ;
    inv02 ix8230 (.Y (nx8231), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix8232 (.Y (nx8233), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix8234 (.Y (nx8235), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv01 ix8236 (.Y (nx8237), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_AddPToBoothOperand)) ;
    inv02 ix8238 (.Y (nx8239), .A (nx8237)) ;
    inv02 ix8240 (.Y (nx8241), .A (nx8237)) ;
    inv02 ix8242 (.Y (nx8243), .A (nx8237)) ;
    inv02 ix8244 (.Y (nx8245), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix8246 (.Y (nx8247), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix8248 (.Y (nx8249), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv01 ix8250 (.Y (nx8251), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_nx80)) ;
    inv02 ix8252 (.Y (nx8253), .A (nx8251)) ;
    inv02 ix8254 (.Y (nx8255), .A (nx8251)) ;
    inv02 ix8256 (.Y (nx8257), .A (nx8251)) ;
    inv02 ix8258 (.Y (nx8259), .A (CALCULATOR_Start_dup_1326)) ;
    inv02 ix8260 (.Y (nx8261), .A (CALCULATOR_Start_dup_1326)) ;
    inv02 ix8262 (.Y (nx8263), .A (CALCULATOR_Start_dup_1326)) ;
    inv02 ix8264 (.Y (nx8265), .A (CALCULATOR_Start_dup_1326)) ;
    inv02 ix8266 (.Y (nx8267), .A (CALCULATOR_Start_dup_1326)) ;
    inv02 ix8268 (.Y (nx8269), .A (CALCULATOR_Start_dup_1326)) ;
    inv02 ix8270 (.Y (nx8271), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix8272 (.Y (nx8273), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix8274 (.Y (nx8275), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv01 ix8276 (.Y (nx8277), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_AddPToBoothOperand)) ;
    inv02 ix8278 (.Y (nx8279), .A (nx8277)) ;
    inv02 ix8280 (.Y (nx8281), .A (nx8277)) ;
    inv02 ix8282 (.Y (nx8283), .A (nx8277)) ;
    inv02 ix8284 (.Y (nx8285), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix8286 (.Y (nx8287), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix8288 (.Y (nx8289), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv01 ix8290 (.Y (nx8291), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_nx80)) ;
    inv02 ix8292 (.Y (nx8293), .A (nx8291)) ;
    inv02 ix8294 (.Y (nx8295), .A (nx8291)) ;
    inv02 ix8296 (.Y (nx8297), .A (nx8291)) ;
    inv02 ix8298 (.Y (nx8299), .A (CALCULATOR_Start_dup_1339)) ;
    inv02 ix8300 (.Y (nx8301), .A (CALCULATOR_Start_dup_1339)) ;
    inv02 ix8302 (.Y (nx8303), .A (CALCULATOR_Start_dup_1339)) ;
    inv02 ix8304 (.Y (nx8305), .A (CALCULATOR_Start_dup_1339)) ;
    inv02 ix8306 (.Y (nx8307), .A (CALCULATOR_Start_dup_1339)) ;
    inv02 ix8308 (.Y (nx8309), .A (CALCULATOR_Start_dup_1339)) ;
    inv02 ix8310 (.Y (nx8311), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix8312 (.Y (nx8313), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix8314 (.Y (nx8315), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv01 ix8316 (.Y (nx8317), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_AddPToBoothOperand)) ;
    inv02 ix8318 (.Y (nx8319), .A (nx8317)) ;
    inv02 ix8320 (.Y (nx8321), .A (nx8317)) ;
    inv02 ix8322 (.Y (nx8323), .A (nx8317)) ;
    inv02 ix8324 (.Y (nx8325), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix8326 (.Y (nx8327), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix8328 (.Y (nx8329), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv01 ix8330 (.Y (nx8331), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_nx80)) ;
    inv02 ix8332 (.Y (nx8333), .A (nx8331)) ;
    inv02 ix8334 (.Y (nx8335), .A (nx8331)) ;
    inv02 ix8336 (.Y (nx8337), .A (nx8331)) ;
    inv02 ix8338 (.Y (nx8339), .A (CALCULATOR_Start_dup_1352)) ;
    inv02 ix8340 (.Y (nx8341), .A (CALCULATOR_Start_dup_1352)) ;
    inv02 ix8342 (.Y (nx8343), .A (CALCULATOR_Start_dup_1352)) ;
    inv02 ix8344 (.Y (nx8345), .A (CALCULATOR_Start_dup_1352)) ;
    inv02 ix8346 (.Y (nx8347), .A (CALCULATOR_Start_dup_1352)) ;
    inv02 ix8348 (.Y (nx8349), .A (CALCULATOR_Start_dup_1352)) ;
    inv02 ix8350 (.Y (nx8351), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix8352 (.Y (nx8353), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix8354 (.Y (nx8355), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 CACHE_ix974_rep_1 (.Y (nx8357), .A (nx8459)) ;
    inv02 CACHE_ix974_rep_2 (.Y (nx8359), .A (nx8459)) ;
    inv02 CACHE_ix976_rep_1 (.Y (nx8361), .A (nx8459)) ;
    inv02 CACHE_ix976_rep_2 (.Y (nx8363), .A (nx8459)) ;
    inv02 CACHE_ix978_rep_1 (.Y (nx8365), .A (nx8459)) ;
    inv02 CACHE_ix978_rep_2 (.Y (nx8367), .A (nx8459)) ;
    inv02 CACHE_ix980_rep_1 (.Y (nx8369), .A (nx8459)) ;
    inv02 CACHE_ix980_rep_2 (.Y (nx8371), .A (nx8841)) ;
    inv02 CACHE_ix982_rep_1 (.Y (nx8373), .A (nx8841)) ;
    inv02 CACHE_ix982_rep_2 (.Y (nx8375), .A (nx8841)) ;
    inv02 CACHE_ix984_rep_1 (.Y (nx8377), .A (nx8841)) ;
    inv02 CACHE_ix984_rep_2 (.Y (nx8379), .A (nx8841)) ;
    inv02 CACHE_ix986_rep_1 (.Y (nx8381), .A (nx8841)) ;
    inv02 CACHE_ix986_rep_2 (.Y (nx8383), .A (nx8841)) ;
    inv02 CACHE_ix988_rep_1 (.Y (nx8385), .A (nx8463)) ;
    inv02 CACHE_ix988_rep_2 (.Y (nx8387), .A (nx8463)) ;
    inv02 CACHE_ix990_rep_1 (.Y (nx8389), .A (nx8463)) ;
    inv02 CACHE_ix990_rep_2 (.Y (nx8391), .A (nx8463)) ;
    inv02 CACHE_ix992_rep_1 (.Y (nx8393), .A (nx8463)) ;
    inv02 CACHE_ix992_rep_2 (.Y (nx8395), .A (nx8463)) ;
    inv02 CACHE_ix994_rep_1 (.Y (nx8397), .A (nx8463)) ;
    inv02 CACHE_ix994_rep_2 (.Y (nx8399), .A (CACHE_nx1043)) ;
    inv02 CACHE_ix996_rep_1 (.Y (nx8401), .A (CACHE_nx1043)) ;
    inv02 CACHE_ix996_rep_2 (.Y (nx8403), .A (CACHE_nx1043)) ;
    inv02 CACHE_ix998_rep_1 (.Y (nx8405), .A (CACHE_nx1043)) ;
    inv02 CACHE_ix998_rep_2 (.Y (nx8407), .A (CACHE_nx1043)) ;
    inv02 CACHE_ix1000_rep_1 (.Y (nx8409), .A (CACHE_nx1043)) ;
    inv02 CACHE_ix1000_rep_2 (.Y (nx8411), .A (CACHE_nx1043)) ;
    inv02 CACHE_ix1002_rep_1 (.Y (nx8413), .A (nx8467)) ;
    inv02 CACHE_ix1002_rep_2 (.Y (nx8415), .A (nx8467)) ;
    inv02 CACHE_ix1004_rep_1 (.Y (nx8417), .A (nx8467)) ;
    inv02 CACHE_ix1004_rep_2 (.Y (nx8419), .A (nx8467)) ;
    inv02 CACHE_ix1006_rep_1 (.Y (nx8421), .A (nx8467)) ;
    inv02 CACHE_ix1006_rep_2 (.Y (nx8423), .A (nx8467)) ;
    inv02 CACHE_ix1008_rep_1 (.Y (nx8425), .A (nx8467)) ;
    inv02 CACHE_ix1008_rep_2 (.Y (nx8427), .A (CACHE_nx1045)) ;
    inv02 CACHE_ix1010_rep_1 (.Y (nx8429), .A (CACHE_nx1045)) ;
    inv02 CACHE_ix1010_rep_2 (.Y (nx8431), .A (CACHE_nx1045)) ;
    inv02 CACHE_ix1012_rep_1 (.Y (nx8433), .A (CACHE_nx1045)) ;
    inv02 CACHE_ix1012_rep_2 (.Y (nx8435), .A (CACHE_nx1045)) ;
    inv02 CACHE_ix1014_rep_1 (.Y (nx8437), .A (CACHE_nx1045)) ;
    inv02 CACHE_ix1014_rep_2 (.Y (nx8439), .A (CACHE_nx1045)) ;
    inv02 CACHE_ix1016_rep_1 (.Y (nx8441), .A (nx8469)) ;
    inv02 CACHE_ix1016_rep_2 (.Y (nx8443), .A (nx8469)) ;
    inv02 CACHE_ix1018_rep_1 (.Y (nx8445), .A (nx8469)) ;
    inv02 CACHE_ix1018_rep_2 (.Y (nx8447), .A (CACHE_nx1047)) ;
    inv02 CACHE_ix1020_rep_1 (.Y (nx8449), .A (CACHE_nx1047)) ;
    inv02 CACHE_ix1020_rep_2 (.Y (nx8451), .A (CACHE_nx1047)) ;
    inv02 CACHE_ix1022_rep_1 (.Y (nx8453), .A (CACHE_nx1047)) ;
    inv02 CACHE_ix1022_rep_2 (.Y (nx8455), .A (CACHE_nx1047)) ;
    inv02 CACHE_ix1040_rep_1 (.Y (nx8457), .A (nx8833)) ;
    inv02 CACHE_ix1040_rep_2 (.Y (nx8459), .A (nx8833)) ;
    inv02 CACHE_ix1042_rep_1 (.Y (nx8461), .A (nx8833)) ;
    inv02 CACHE_ix1042_rep_2 (.Y (nx8463), .A (nx8833)) ;
    inv02 CACHE_ix1044_rep_1 (.Y (nx8465), .A (nx8835)) ;
    inv02 CACHE_ix1044_rep_2 (.Y (nx8467), .A (nx8835)) ;
    inv02 CACHE_ix1046_rep_1 (.Y (nx8469), .A (nx8835)) ;
    inv02 ix8470 (.Y (nx8471), .A (CONTROLLER_ROW_nx296)) ;
    inv02 ix8472 (.Y (nx8473), .A (CONTROLLER_ROW_nx296)) ;
    inv02 ix8474 (.Y (nx8475), .A (CONTROLLER_COL_nx296)) ;
    inv02 ix8476 (.Y (nx8477), .A (CONTROLLER_COL_nx296)) ;
    inv02 ix8478 (.Y (nx8479), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8480 (.Y (nx8481), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8482 (.Y (nx8483), .A (
          CALCULATOR_L1_0_L2_0_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8484 (.Y (nx8485), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8486 (.Y (nx8487), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8488 (.Y (nx8489), .A (
          CALCULATOR_L1_0_L2_1_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8490 (.Y (nx8491), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8492 (.Y (nx8493), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8494 (.Y (nx8495), .A (
          CALCULATOR_L1_0_L2_2_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8496 (.Y (nx8497), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8498 (.Y (nx8499), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8500 (.Y (nx8501), .A (
          CALCULATOR_L1_0_L2_3_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8502 (.Y (nx8503), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8504 (.Y (nx8505), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8506 (.Y (nx8507), .A (
          CALCULATOR_L1_0_L2_4_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8508 (.Y (nx8509), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8510 (.Y (nx8511), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8512 (.Y (nx8513), .A (
          CALCULATOR_L1_1_L2_0_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8514 (.Y (nx8515), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8516 (.Y (nx8517), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8518 (.Y (nx8519), .A (
          CALCULATOR_L1_1_L2_1_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8520 (.Y (nx8521), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8522 (.Y (nx8523), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8524 (.Y (nx8525), .A (
          CALCULATOR_L1_1_L2_2_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8526 (.Y (nx8527), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8528 (.Y (nx8529), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8530 (.Y (nx8531), .A (
          CALCULATOR_L1_1_L2_3_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8532 (.Y (nx8533), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8534 (.Y (nx8535), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8536 (.Y (nx8537), .A (
          CALCULATOR_L1_1_L2_4_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8538 (.Y (nx8539), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8540 (.Y (nx8541), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8542 (.Y (nx8543), .A (
          CALCULATOR_L1_2_L2_0_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8544 (.Y (nx8545), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8546 (.Y (nx8547), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8548 (.Y (nx8549), .A (
          CALCULATOR_L1_2_L2_1_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8550 (.Y (nx8551), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8552 (.Y (nx8553), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8554 (.Y (nx8555), .A (
          CALCULATOR_L1_2_L2_2_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8556 (.Y (nx8557), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8558 (.Y (nx8559), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8560 (.Y (nx8561), .A (
          CALCULATOR_L1_2_L2_3_G2_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8562 (.Y (nx8563), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8564 (.Y (nx8565), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8566 (.Y (nx8567), .A (
          CALCULATOR_L1_2_L2_4_G2_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8568 (.Y (nx8569), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8570 (.Y (nx8571), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8572 (.Y (nx8573), .A (
          CALCULATOR_L1_3_L2_0_G2_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8574 (.Y (nx8575), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8576 (.Y (nx8577), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8578 (.Y (nx8579), .A (
          CALCULATOR_L1_3_L2_1_G2_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8580 (.Y (nx8581), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8582 (.Y (nx8583), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8584 (.Y (nx8585), .A (
          CALCULATOR_L1_3_L2_2_G2_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8586 (.Y (nx8587), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8588 (.Y (nx8589), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8590 (.Y (nx8591), .A (
          CALCULATOR_L1_3_L2_3_G2_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8592 (.Y (nx8593), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8594 (.Y (nx8595), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8596 (.Y (nx8597), .A (
          CALCULATOR_L1_3_L2_4_G3_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8598 (.Y (nx8599), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8600 (.Y (nx8601), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8602 (.Y (nx8603), .A (
          CALCULATOR_L1_4_L2_0_G3_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8604 (.Y (nx8605), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8606 (.Y (nx8607), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8608 (.Y (nx8609), .A (
          CALCULATOR_L1_4_L2_1_G3_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8610 (.Y (nx8611), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8612 (.Y (nx8613), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8614 (.Y (nx8615), .A (
          CALCULATOR_L1_4_L2_2_G4_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8616 (.Y (nx8617), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8618 (.Y (nx8619), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8620 (.Y (nx8621), .A (
          CALCULATOR_L1_4_L2_3_G5_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8622 (.Y (nx8623), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8624 (.Y (nx8625), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8626 (.Y (nx8627), .A (
          CALCULATOR_L1_4_L2_4_G5_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8628 (.Y (nx8629), .A (CACHE_L0_0_L1_0_Fij_nx296)) ;
    inv02 ix8630 (.Y (nx8631), .A (CACHE_L0_0_L1_0_Fij_nx296)) ;
    inv02 ix8632 (.Y (nx8633), .A (CACHE_L0_0_L1_0_Wij_nx296)) ;
    inv02 ix8634 (.Y (nx8635), .A (CACHE_L0_0_L1_0_Wij_nx296)) ;
    inv02 ix8636 (.Y (nx8637), .A (CACHE_L0_0_L1_1_Fij_nx296)) ;
    inv02 ix8638 (.Y (nx8639), .A (CACHE_L0_0_L1_1_Fij_nx296)) ;
    inv02 ix8640 (.Y (nx8641), .A (CACHE_L0_0_L1_1_Wij_nx296)) ;
    inv02 ix8642 (.Y (nx8643), .A (CACHE_L0_0_L1_1_Wij_nx296)) ;
    inv02 ix8644 (.Y (nx8645), .A (CACHE_L0_0_L1_2_Fij_nx296)) ;
    inv02 ix8646 (.Y (nx8647), .A (CACHE_L0_0_L1_2_Fij_nx296)) ;
    inv02 ix8648 (.Y (nx8649), .A (CACHE_L0_0_L1_2_Wij_nx296)) ;
    inv02 ix8650 (.Y (nx8651), .A (CACHE_L0_0_L1_2_Wij_nx296)) ;
    inv02 ix8652 (.Y (nx8653), .A (CACHE_L0_0_L1_3_Fij_nx296)) ;
    inv02 ix8654 (.Y (nx8655), .A (CACHE_L0_0_L1_3_Fij_nx296)) ;
    inv02 ix8656 (.Y (nx8657), .A (CACHE_L0_0_L1_3_Wij_nx296)) ;
    inv02 ix8658 (.Y (nx8659), .A (CACHE_L0_0_L1_3_Wij_nx296)) ;
    inv02 ix8660 (.Y (nx8661), .A (CACHE_L0_0_L1_4_Fij_nx296)) ;
    inv02 ix8662 (.Y (nx8663), .A (CACHE_L0_0_L1_4_Fij_nx296)) ;
    inv02 ix8664 (.Y (nx8665), .A (CACHE_L0_0_L1_4_Wij_nx296)) ;
    inv02 ix8666 (.Y (nx8667), .A (CACHE_L0_0_L1_4_Wij_nx296)) ;
    inv02 ix8668 (.Y (nx8669), .A (CACHE_L0_1_L1_0_Fij_nx296)) ;
    inv02 ix8670 (.Y (nx8671), .A (CACHE_L0_1_L1_0_Fij_nx296)) ;
    inv02 ix8672 (.Y (nx8673), .A (CACHE_L0_1_L1_0_Wij_nx296)) ;
    inv02 ix8674 (.Y (nx8675), .A (CACHE_L0_1_L1_0_Wij_nx296)) ;
    inv02 ix8676 (.Y (nx8677), .A (CACHE_L0_1_L1_1_Fij_nx296)) ;
    inv02 ix8678 (.Y (nx8679), .A (CACHE_L0_1_L1_1_Fij_nx296)) ;
    inv02 ix8680 (.Y (nx8681), .A (CACHE_L0_1_L1_1_Wij_nx296)) ;
    inv02 ix8682 (.Y (nx8683), .A (CACHE_L0_1_L1_1_Wij_nx296)) ;
    inv02 ix8684 (.Y (nx8685), .A (CACHE_L0_1_L1_2_Fij_nx296)) ;
    inv02 ix8686 (.Y (nx8687), .A (CACHE_L0_1_L1_2_Fij_nx296)) ;
    inv02 ix8688 (.Y (nx8689), .A (CACHE_L0_1_L1_2_Wij_nx296)) ;
    inv02 ix8690 (.Y (nx8691), .A (CACHE_L0_1_L1_2_Wij_nx296)) ;
    inv02 ix8692 (.Y (nx8693), .A (CACHE_L0_1_L1_3_Fij_nx296)) ;
    inv02 ix8694 (.Y (nx8695), .A (CACHE_L0_1_L1_3_Fij_nx296)) ;
    inv02 ix8696 (.Y (nx8697), .A (CACHE_L0_1_L1_3_Wij_nx296)) ;
    inv02 ix8698 (.Y (nx8699), .A (CACHE_L0_1_L1_3_Wij_nx296)) ;
    inv02 ix8700 (.Y (nx8701), .A (CACHE_L0_1_L1_4_Fij_nx296)) ;
    inv02 ix8702 (.Y (nx8703), .A (CACHE_L0_1_L1_4_Fij_nx296)) ;
    inv02 ix8704 (.Y (nx8705), .A (CACHE_L0_1_L1_4_Wij_nx296)) ;
    inv02 ix8706 (.Y (nx8707), .A (CACHE_L0_1_L1_4_Wij_nx296)) ;
    inv02 ix8708 (.Y (nx8709), .A (CACHE_L0_2_L1_0_Fij_nx296)) ;
    inv02 ix8710 (.Y (nx8711), .A (CACHE_L0_2_L1_0_Fij_nx296)) ;
    inv02 ix8712 (.Y (nx8713), .A (CACHE_L0_2_L1_0_Wij_nx296)) ;
    inv02 ix8714 (.Y (nx8715), .A (CACHE_L0_2_L1_0_Wij_nx296)) ;
    inv02 ix8716 (.Y (nx8717), .A (CACHE_L0_2_L1_1_Fij_nx296)) ;
    inv02 ix8718 (.Y (nx8719), .A (CACHE_L0_2_L1_1_Fij_nx296)) ;
    inv02 ix8720 (.Y (nx8721), .A (CACHE_L0_2_L1_1_Wij_nx296)) ;
    inv02 ix8722 (.Y (nx8723), .A (CACHE_L0_2_L1_1_Wij_nx296)) ;
    inv02 ix8724 (.Y (nx8725), .A (CACHE_L0_2_L1_2_Fij_nx296)) ;
    inv02 ix8726 (.Y (nx8727), .A (CACHE_L0_2_L1_2_Fij_nx296)) ;
    inv02 ix8728 (.Y (nx8729), .A (CACHE_L0_2_L1_2_Wij_nx296)) ;
    inv02 ix8730 (.Y (nx8731), .A (CACHE_L0_2_L1_2_Wij_nx296)) ;
    inv02 ix8732 (.Y (nx8733), .A (CACHE_L0_2_L1_3_Fij_nx296)) ;
    inv02 ix8734 (.Y (nx8735), .A (CACHE_L0_2_L1_3_Fij_nx296)) ;
    inv02 ix8736 (.Y (nx8737), .A (CACHE_L0_2_L1_3_Wij_nx296)) ;
    inv02 ix8738 (.Y (nx8739), .A (CACHE_L0_2_L1_3_Wij_nx296)) ;
    inv02 ix8740 (.Y (nx8741), .A (CACHE_L0_2_L1_4_Fij_nx296)) ;
    inv02 ix8742 (.Y (nx8743), .A (CACHE_L0_2_L1_4_Fij_nx296)) ;
    inv02 ix8744 (.Y (nx8745), .A (CACHE_L0_2_L1_4_Wij_nx296)) ;
    inv02 ix8746 (.Y (nx8747), .A (CACHE_L0_2_L1_4_Wij_nx296)) ;
    inv02 ix8748 (.Y (nx8749), .A (CACHE_L0_3_L1_0_Fij_nx296)) ;
    inv02 ix8750 (.Y (nx8751), .A (CACHE_L0_3_L1_0_Fij_nx296)) ;
    inv02 ix8752 (.Y (nx8753), .A (CACHE_L0_3_L1_0_Wij_nx296)) ;
    inv02 ix8754 (.Y (nx8755), .A (CACHE_L0_3_L1_0_Wij_nx296)) ;
    inv02 ix8756 (.Y (nx8757), .A (CACHE_L0_3_L1_1_Fij_nx296)) ;
    inv02 ix8758 (.Y (nx8759), .A (CACHE_L0_3_L1_1_Fij_nx296)) ;
    inv02 ix8760 (.Y (nx8761), .A (CACHE_L0_3_L1_1_Wij_nx296)) ;
    inv02 ix8762 (.Y (nx8763), .A (CACHE_L0_3_L1_1_Wij_nx296)) ;
    inv02 ix8764 (.Y (nx8765), .A (CACHE_L0_3_L1_2_Fij_nx296)) ;
    inv02 ix8766 (.Y (nx8767), .A (CACHE_L0_3_L1_2_Fij_nx296)) ;
    inv02 ix8768 (.Y (nx8769), .A (CACHE_L0_3_L1_2_Wij_nx296)) ;
    inv02 ix8770 (.Y (nx8771), .A (CACHE_L0_3_L1_2_Wij_nx296)) ;
    inv02 ix8772 (.Y (nx8773), .A (CACHE_L0_3_L1_3_Fij_nx296)) ;
    inv02 ix8774 (.Y (nx8775), .A (CACHE_L0_3_L1_3_Fij_nx296)) ;
    inv02 ix8776 (.Y (nx8777), .A (CACHE_L0_3_L1_3_Wij_nx296)) ;
    inv02 ix8778 (.Y (nx8779), .A (CACHE_L0_3_L1_3_Wij_nx296)) ;
    inv02 ix8780 (.Y (nx8781), .A (CACHE_L0_3_L1_4_Fij_nx296)) ;
    inv02 ix8782 (.Y (nx8783), .A (CACHE_L0_3_L1_4_Fij_nx296)) ;
    inv02 ix8784 (.Y (nx8785), .A (CACHE_L0_3_L1_4_Wij_nx296)) ;
    inv02 ix8786 (.Y (nx8787), .A (CACHE_L0_3_L1_4_Wij_nx296)) ;
    inv02 ix8788 (.Y (nx8789), .A (CACHE_L0_4_L1_0_Fij_nx296)) ;
    inv02 ix8790 (.Y (nx8791), .A (CACHE_L0_4_L1_0_Fij_nx296)) ;
    inv02 ix8792 (.Y (nx8793), .A (CACHE_L0_4_L1_0_Wij_nx296)) ;
    inv02 ix8794 (.Y (nx8795), .A (CACHE_L0_4_L1_0_Wij_nx296)) ;
    inv02 ix8796 (.Y (nx8797), .A (CACHE_L0_4_L1_1_Fij_nx296)) ;
    inv02 ix8798 (.Y (nx8799), .A (CACHE_L0_4_L1_1_Fij_nx296)) ;
    inv02 ix8800 (.Y (nx8801), .A (CACHE_L0_4_L1_1_Wij_nx296)) ;
    inv02 ix8802 (.Y (nx8803), .A (CACHE_L0_4_L1_1_Wij_nx296)) ;
    inv02 ix8804 (.Y (nx8805), .A (CACHE_L0_4_L1_2_Fij_nx296)) ;
    inv02 ix8806 (.Y (nx8807), .A (CACHE_L0_4_L1_2_Fij_nx296)) ;
    inv02 ix8808 (.Y (nx8809), .A (CACHE_L0_4_L1_2_Wij_nx296)) ;
    inv02 ix8810 (.Y (nx8811), .A (CACHE_L0_4_L1_2_Wij_nx296)) ;
    inv02 ix8812 (.Y (nx8813), .A (CACHE_L0_4_L1_3_Fij_nx296)) ;
    inv02 ix8814 (.Y (nx8815), .A (CACHE_L0_4_L1_3_Fij_nx296)) ;
    inv02 ix8816 (.Y (nx8817), .A (CACHE_L0_4_L1_3_Wij_nx296)) ;
    inv02 ix8818 (.Y (nx8819), .A (CACHE_L0_4_L1_3_Wij_nx296)) ;
    inv02 ix8820 (.Y (nx8821), .A (CACHE_L0_4_L1_4_Fij_nx296)) ;
    inv02 ix8822 (.Y (nx8823), .A (CACHE_L0_4_L1_4_Fij_nx296)) ;
    inv02 ix8824 (.Y (nx8825), .A (CACHE_L0_4_L1_4_Wij_nx296)) ;
    inv02 ix8826 (.Y (nx8827), .A (CACHE_L0_4_L1_4_Wij_nx296)) ;
    inv02 ix8832 (.Y (nx8833), .A (CACHE_nx1041)) ;
    inv02 ix8834 (.Y (nx8835), .A (CACHE_nx1041)) ;
    inv01 ix8836 (.Y (nx8837), .A (CALCULATOR_nx1111)) ;
    inv01 ix8838 (.Y (nx8839), .A (CALCULATOR_nx1111)) ;
    inv02 CACHE_ix1040_rep_3 (.Y (nx8841), .A (CacheRST)) ;
endmodule

