//
// Verilog description for cell cache, 
// Sat May 12 15:09:25 2018
//
// LeonardoSpectrum Level 3, 2017a.2 
//


module cache ( CLK, RST, FilterSize, FilterWR, WindowWR, Din, FilterDout_0__0__7, 
               FilterDout_0__0__6, FilterDout_0__0__5, FilterDout_0__0__4, 
               FilterDout_0__0__3, FilterDout_0__0__2, FilterDout_0__0__1, 
               FilterDout_0__0__0, FilterDout_0__1__7, FilterDout_0__1__6, 
               FilterDout_0__1__5, FilterDout_0__1__4, FilterDout_0__1__3, 
               FilterDout_0__1__2, FilterDout_0__1__1, FilterDout_0__1__0, 
               FilterDout_0__2__7, FilterDout_0__2__6, FilterDout_0__2__5, 
               FilterDout_0__2__4, FilterDout_0__2__3, FilterDout_0__2__2, 
               FilterDout_0__2__1, FilterDout_0__2__0, FilterDout_0__3__7, 
               FilterDout_0__3__6, FilterDout_0__3__5, FilterDout_0__3__4, 
               FilterDout_0__3__3, FilterDout_0__3__2, FilterDout_0__3__1, 
               FilterDout_0__3__0, FilterDout_0__4__7, FilterDout_0__4__6, 
               FilterDout_0__4__5, FilterDout_0__4__4, FilterDout_0__4__3, 
               FilterDout_0__4__2, FilterDout_0__4__1, FilterDout_0__4__0, 
               FilterDout_1__0__7, FilterDout_1__0__6, FilterDout_1__0__5, 
               FilterDout_1__0__4, FilterDout_1__0__3, FilterDout_1__0__2, 
               FilterDout_1__0__1, FilterDout_1__0__0, FilterDout_1__1__7, 
               FilterDout_1__1__6, FilterDout_1__1__5, FilterDout_1__1__4, 
               FilterDout_1__1__3, FilterDout_1__1__2, FilterDout_1__1__1, 
               FilterDout_1__1__0, FilterDout_1__2__7, FilterDout_1__2__6, 
               FilterDout_1__2__5, FilterDout_1__2__4, FilterDout_1__2__3, 
               FilterDout_1__2__2, FilterDout_1__2__1, FilterDout_1__2__0, 
               FilterDout_1__3__7, FilterDout_1__3__6, FilterDout_1__3__5, 
               FilterDout_1__3__4, FilterDout_1__3__3, FilterDout_1__3__2, 
               FilterDout_1__3__1, FilterDout_1__3__0, FilterDout_1__4__7, 
               FilterDout_1__4__6, FilterDout_1__4__5, FilterDout_1__4__4, 
               FilterDout_1__4__3, FilterDout_1__4__2, FilterDout_1__4__1, 
               FilterDout_1__4__0, FilterDout_2__0__7, FilterDout_2__0__6, 
               FilterDout_2__0__5, FilterDout_2__0__4, FilterDout_2__0__3, 
               FilterDout_2__0__2, FilterDout_2__0__1, FilterDout_2__0__0, 
               FilterDout_2__1__7, FilterDout_2__1__6, FilterDout_2__1__5, 
               FilterDout_2__1__4, FilterDout_2__1__3, FilterDout_2__1__2, 
               FilterDout_2__1__1, FilterDout_2__1__0, FilterDout_2__2__7, 
               FilterDout_2__2__6, FilterDout_2__2__5, FilterDout_2__2__4, 
               FilterDout_2__2__3, FilterDout_2__2__2, FilterDout_2__2__1, 
               FilterDout_2__2__0, FilterDout_2__3__7, FilterDout_2__3__6, 
               FilterDout_2__3__5, FilterDout_2__3__4, FilterDout_2__3__3, 
               FilterDout_2__3__2, FilterDout_2__3__1, FilterDout_2__3__0, 
               FilterDout_2__4__7, FilterDout_2__4__6, FilterDout_2__4__5, 
               FilterDout_2__4__4, FilterDout_2__4__3, FilterDout_2__4__2, 
               FilterDout_2__4__1, FilterDout_2__4__0, FilterDout_3__0__7, 
               FilterDout_3__0__6, FilterDout_3__0__5, FilterDout_3__0__4, 
               FilterDout_3__0__3, FilterDout_3__0__2, FilterDout_3__0__1, 
               FilterDout_3__0__0, FilterDout_3__1__7, FilterDout_3__1__6, 
               FilterDout_3__1__5, FilterDout_3__1__4, FilterDout_3__1__3, 
               FilterDout_3__1__2, FilterDout_3__1__1, FilterDout_3__1__0, 
               FilterDout_3__2__7, FilterDout_3__2__6, FilterDout_3__2__5, 
               FilterDout_3__2__4, FilterDout_3__2__3, FilterDout_3__2__2, 
               FilterDout_3__2__1, FilterDout_3__2__0, FilterDout_3__3__7, 
               FilterDout_3__3__6, FilterDout_3__3__5, FilterDout_3__3__4, 
               FilterDout_3__3__3, FilterDout_3__3__2, FilterDout_3__3__1, 
               FilterDout_3__3__0, FilterDout_3__4__7, FilterDout_3__4__6, 
               FilterDout_3__4__5, FilterDout_3__4__4, FilterDout_3__4__3, 
               FilterDout_3__4__2, FilterDout_3__4__1, FilterDout_3__4__0, 
               FilterDout_4__0__7, FilterDout_4__0__6, FilterDout_4__0__5, 
               FilterDout_4__0__4, FilterDout_4__0__3, FilterDout_4__0__2, 
               FilterDout_4__0__1, FilterDout_4__0__0, FilterDout_4__1__7, 
               FilterDout_4__1__6, FilterDout_4__1__5, FilterDout_4__1__4, 
               FilterDout_4__1__3, FilterDout_4__1__2, FilterDout_4__1__1, 
               FilterDout_4__1__0, FilterDout_4__2__7, FilterDout_4__2__6, 
               FilterDout_4__2__5, FilterDout_4__2__4, FilterDout_4__2__3, 
               FilterDout_4__2__2, FilterDout_4__2__1, FilterDout_4__2__0, 
               FilterDout_4__3__7, FilterDout_4__3__6, FilterDout_4__3__5, 
               FilterDout_4__3__4, FilterDout_4__3__3, FilterDout_4__3__2, 
               FilterDout_4__3__1, FilterDout_4__3__0, FilterDout_4__4__7, 
               FilterDout_4__4__6, FilterDout_4__4__5, FilterDout_4__4__4, 
               FilterDout_4__4__3, FilterDout_4__4__2, FilterDout_4__4__1, 
               FilterDout_4__4__0, WindowDout_0__0__7, WindowDout_0__0__6, 
               WindowDout_0__0__5, WindowDout_0__0__4, WindowDout_0__0__3, 
               WindowDout_0__0__2, WindowDout_0__0__1, WindowDout_0__0__0, 
               WindowDout_0__1__7, WindowDout_0__1__6, WindowDout_0__1__5, 
               WindowDout_0__1__4, WindowDout_0__1__3, WindowDout_0__1__2, 
               WindowDout_0__1__1, WindowDout_0__1__0, WindowDout_0__2__7, 
               WindowDout_0__2__6, WindowDout_0__2__5, WindowDout_0__2__4, 
               WindowDout_0__2__3, WindowDout_0__2__2, WindowDout_0__2__1, 
               WindowDout_0__2__0, WindowDout_0__3__7, WindowDout_0__3__6, 
               WindowDout_0__3__5, WindowDout_0__3__4, WindowDout_0__3__3, 
               WindowDout_0__3__2, WindowDout_0__3__1, WindowDout_0__3__0, 
               WindowDout_0__4__7, WindowDout_0__4__6, WindowDout_0__4__5, 
               WindowDout_0__4__4, WindowDout_0__4__3, WindowDout_0__4__2, 
               WindowDout_0__4__1, WindowDout_0__4__0, WindowDout_1__0__7, 
               WindowDout_1__0__6, WindowDout_1__0__5, WindowDout_1__0__4, 
               WindowDout_1__0__3, WindowDout_1__0__2, WindowDout_1__0__1, 
               WindowDout_1__0__0, WindowDout_1__1__7, WindowDout_1__1__6, 
               WindowDout_1__1__5, WindowDout_1__1__4, WindowDout_1__1__3, 
               WindowDout_1__1__2, WindowDout_1__1__1, WindowDout_1__1__0, 
               WindowDout_1__2__7, WindowDout_1__2__6, WindowDout_1__2__5, 
               WindowDout_1__2__4, WindowDout_1__2__3, WindowDout_1__2__2, 
               WindowDout_1__2__1, WindowDout_1__2__0, WindowDout_1__3__7, 
               WindowDout_1__3__6, WindowDout_1__3__5, WindowDout_1__3__4, 
               WindowDout_1__3__3, WindowDout_1__3__2, WindowDout_1__3__1, 
               WindowDout_1__3__0, WindowDout_1__4__7, WindowDout_1__4__6, 
               WindowDout_1__4__5, WindowDout_1__4__4, WindowDout_1__4__3, 
               WindowDout_1__4__2, WindowDout_1__4__1, WindowDout_1__4__0, 
               WindowDout_2__0__7, WindowDout_2__0__6, WindowDout_2__0__5, 
               WindowDout_2__0__4, WindowDout_2__0__3, WindowDout_2__0__2, 
               WindowDout_2__0__1, WindowDout_2__0__0, WindowDout_2__1__7, 
               WindowDout_2__1__6, WindowDout_2__1__5, WindowDout_2__1__4, 
               WindowDout_2__1__3, WindowDout_2__1__2, WindowDout_2__1__1, 
               WindowDout_2__1__0, WindowDout_2__2__7, WindowDout_2__2__6, 
               WindowDout_2__2__5, WindowDout_2__2__4, WindowDout_2__2__3, 
               WindowDout_2__2__2, WindowDout_2__2__1, WindowDout_2__2__0, 
               WindowDout_2__3__7, WindowDout_2__3__6, WindowDout_2__3__5, 
               WindowDout_2__3__4, WindowDout_2__3__3, WindowDout_2__3__2, 
               WindowDout_2__3__1, WindowDout_2__3__0, WindowDout_2__4__7, 
               WindowDout_2__4__6, WindowDout_2__4__5, WindowDout_2__4__4, 
               WindowDout_2__4__3, WindowDout_2__4__2, WindowDout_2__4__1, 
               WindowDout_2__4__0, WindowDout_3__0__7, WindowDout_3__0__6, 
               WindowDout_3__0__5, WindowDout_3__0__4, WindowDout_3__0__3, 
               WindowDout_3__0__2, WindowDout_3__0__1, WindowDout_3__0__0, 
               WindowDout_3__1__7, WindowDout_3__1__6, WindowDout_3__1__5, 
               WindowDout_3__1__4, WindowDout_3__1__3, WindowDout_3__1__2, 
               WindowDout_3__1__1, WindowDout_3__1__0, WindowDout_3__2__7, 
               WindowDout_3__2__6, WindowDout_3__2__5, WindowDout_3__2__4, 
               WindowDout_3__2__3, WindowDout_3__2__2, WindowDout_3__2__1, 
               WindowDout_3__2__0, WindowDout_3__3__7, WindowDout_3__3__6, 
               WindowDout_3__3__5, WindowDout_3__3__4, WindowDout_3__3__3, 
               WindowDout_3__3__2, WindowDout_3__3__1, WindowDout_3__3__0, 
               WindowDout_3__4__7, WindowDout_3__4__6, WindowDout_3__4__5, 
               WindowDout_3__4__4, WindowDout_3__4__3, WindowDout_3__4__2, 
               WindowDout_3__4__1, WindowDout_3__4__0, WindowDout_4__0__7, 
               WindowDout_4__0__6, WindowDout_4__0__5, WindowDout_4__0__4, 
               WindowDout_4__0__3, WindowDout_4__0__2, WindowDout_4__0__1, 
               WindowDout_4__0__0, WindowDout_4__1__7, WindowDout_4__1__6, 
               WindowDout_4__1__5, WindowDout_4__1__4, WindowDout_4__1__3, 
               WindowDout_4__1__2, WindowDout_4__1__1, WindowDout_4__1__0, 
               WindowDout_4__2__7, WindowDout_4__2__6, WindowDout_4__2__5, 
               WindowDout_4__2__4, WindowDout_4__2__3, WindowDout_4__2__2, 
               WindowDout_4__2__1, WindowDout_4__2__0, WindowDout_4__3__7, 
               WindowDout_4__3__6, WindowDout_4__3__5, WindowDout_4__3__4, 
               WindowDout_4__3__3, WindowDout_4__3__2, WindowDout_4__3__1, 
               WindowDout_4__3__0, WindowDout_4__4__7, WindowDout_4__4__6, 
               WindowDout_4__4__5, WindowDout_4__4__4, WindowDout_4__4__3, 
               WindowDout_4__4__2, WindowDout_4__4__1, WindowDout_4__4__0 ) ;

    input CLK ;
    input RST ;
    input FilterSize ;
    input FilterWR ;
    input WindowWR ;
    input [39:0]Din ;
    output FilterDout_0__0__7 ;
    output FilterDout_0__0__6 ;
    output FilterDout_0__0__5 ;
    output FilterDout_0__0__4 ;
    output FilterDout_0__0__3 ;
    output FilterDout_0__0__2 ;
    output FilterDout_0__0__1 ;
    output FilterDout_0__0__0 ;
    output FilterDout_0__1__7 ;
    output FilterDout_0__1__6 ;
    output FilterDout_0__1__5 ;
    output FilterDout_0__1__4 ;
    output FilterDout_0__1__3 ;
    output FilterDout_0__1__2 ;
    output FilterDout_0__1__1 ;
    output FilterDout_0__1__0 ;
    output FilterDout_0__2__7 ;
    output FilterDout_0__2__6 ;
    output FilterDout_0__2__5 ;
    output FilterDout_0__2__4 ;
    output FilterDout_0__2__3 ;
    output FilterDout_0__2__2 ;
    output FilterDout_0__2__1 ;
    output FilterDout_0__2__0 ;
    output FilterDout_0__3__7 ;
    output FilterDout_0__3__6 ;
    output FilterDout_0__3__5 ;
    output FilterDout_0__3__4 ;
    output FilterDout_0__3__3 ;
    output FilterDout_0__3__2 ;
    output FilterDout_0__3__1 ;
    output FilterDout_0__3__0 ;
    output FilterDout_0__4__7 ;
    output FilterDout_0__4__6 ;
    output FilterDout_0__4__5 ;
    output FilterDout_0__4__4 ;
    output FilterDout_0__4__3 ;
    output FilterDout_0__4__2 ;
    output FilterDout_0__4__1 ;
    output FilterDout_0__4__0 ;
    output FilterDout_1__0__7 ;
    output FilterDout_1__0__6 ;
    output FilterDout_1__0__5 ;
    output FilterDout_1__0__4 ;
    output FilterDout_1__0__3 ;
    output FilterDout_1__0__2 ;
    output FilterDout_1__0__1 ;
    output FilterDout_1__0__0 ;
    output FilterDout_1__1__7 ;
    output FilterDout_1__1__6 ;
    output FilterDout_1__1__5 ;
    output FilterDout_1__1__4 ;
    output FilterDout_1__1__3 ;
    output FilterDout_1__1__2 ;
    output FilterDout_1__1__1 ;
    output FilterDout_1__1__0 ;
    output FilterDout_1__2__7 ;
    output FilterDout_1__2__6 ;
    output FilterDout_1__2__5 ;
    output FilterDout_1__2__4 ;
    output FilterDout_1__2__3 ;
    output FilterDout_1__2__2 ;
    output FilterDout_1__2__1 ;
    output FilterDout_1__2__0 ;
    output FilterDout_1__3__7 ;
    output FilterDout_1__3__6 ;
    output FilterDout_1__3__5 ;
    output FilterDout_1__3__4 ;
    output FilterDout_1__3__3 ;
    output FilterDout_1__3__2 ;
    output FilterDout_1__3__1 ;
    output FilterDout_1__3__0 ;
    output FilterDout_1__4__7 ;
    output FilterDout_1__4__6 ;
    output FilterDout_1__4__5 ;
    output FilterDout_1__4__4 ;
    output FilterDout_1__4__3 ;
    output FilterDout_1__4__2 ;
    output FilterDout_1__4__1 ;
    output FilterDout_1__4__0 ;
    output FilterDout_2__0__7 ;
    output FilterDout_2__0__6 ;
    output FilterDout_2__0__5 ;
    output FilterDout_2__0__4 ;
    output FilterDout_2__0__3 ;
    output FilterDout_2__0__2 ;
    output FilterDout_2__0__1 ;
    output FilterDout_2__0__0 ;
    output FilterDout_2__1__7 ;
    output FilterDout_2__1__6 ;
    output FilterDout_2__1__5 ;
    output FilterDout_2__1__4 ;
    output FilterDout_2__1__3 ;
    output FilterDout_2__1__2 ;
    output FilterDout_2__1__1 ;
    output FilterDout_2__1__0 ;
    output FilterDout_2__2__7 ;
    output FilterDout_2__2__6 ;
    output FilterDout_2__2__5 ;
    output FilterDout_2__2__4 ;
    output FilterDout_2__2__3 ;
    output FilterDout_2__2__2 ;
    output FilterDout_2__2__1 ;
    output FilterDout_2__2__0 ;
    output FilterDout_2__3__7 ;
    output FilterDout_2__3__6 ;
    output FilterDout_2__3__5 ;
    output FilterDout_2__3__4 ;
    output FilterDout_2__3__3 ;
    output FilterDout_2__3__2 ;
    output FilterDout_2__3__1 ;
    output FilterDout_2__3__0 ;
    output FilterDout_2__4__7 ;
    output FilterDout_2__4__6 ;
    output FilterDout_2__4__5 ;
    output FilterDout_2__4__4 ;
    output FilterDout_2__4__3 ;
    output FilterDout_2__4__2 ;
    output FilterDout_2__4__1 ;
    output FilterDout_2__4__0 ;
    output FilterDout_3__0__7 ;
    output FilterDout_3__0__6 ;
    output FilterDout_3__0__5 ;
    output FilterDout_3__0__4 ;
    output FilterDout_3__0__3 ;
    output FilterDout_3__0__2 ;
    output FilterDout_3__0__1 ;
    output FilterDout_3__0__0 ;
    output FilterDout_3__1__7 ;
    output FilterDout_3__1__6 ;
    output FilterDout_3__1__5 ;
    output FilterDout_3__1__4 ;
    output FilterDout_3__1__3 ;
    output FilterDout_3__1__2 ;
    output FilterDout_3__1__1 ;
    output FilterDout_3__1__0 ;
    output FilterDout_3__2__7 ;
    output FilterDout_3__2__6 ;
    output FilterDout_3__2__5 ;
    output FilterDout_3__2__4 ;
    output FilterDout_3__2__3 ;
    output FilterDout_3__2__2 ;
    output FilterDout_3__2__1 ;
    output FilterDout_3__2__0 ;
    output FilterDout_3__3__7 ;
    output FilterDout_3__3__6 ;
    output FilterDout_3__3__5 ;
    output FilterDout_3__3__4 ;
    output FilterDout_3__3__3 ;
    output FilterDout_3__3__2 ;
    output FilterDout_3__3__1 ;
    output FilterDout_3__3__0 ;
    output FilterDout_3__4__7 ;
    output FilterDout_3__4__6 ;
    output FilterDout_3__4__5 ;
    output FilterDout_3__4__4 ;
    output FilterDout_3__4__3 ;
    output FilterDout_3__4__2 ;
    output FilterDout_3__4__1 ;
    output FilterDout_3__4__0 ;
    output FilterDout_4__0__7 ;
    output FilterDout_4__0__6 ;
    output FilterDout_4__0__5 ;
    output FilterDout_4__0__4 ;
    output FilterDout_4__0__3 ;
    output FilterDout_4__0__2 ;
    output FilterDout_4__0__1 ;
    output FilterDout_4__0__0 ;
    output FilterDout_4__1__7 ;
    output FilterDout_4__1__6 ;
    output FilterDout_4__1__5 ;
    output FilterDout_4__1__4 ;
    output FilterDout_4__1__3 ;
    output FilterDout_4__1__2 ;
    output FilterDout_4__1__1 ;
    output FilterDout_4__1__0 ;
    output FilterDout_4__2__7 ;
    output FilterDout_4__2__6 ;
    output FilterDout_4__2__5 ;
    output FilterDout_4__2__4 ;
    output FilterDout_4__2__3 ;
    output FilterDout_4__2__2 ;
    output FilterDout_4__2__1 ;
    output FilterDout_4__2__0 ;
    output FilterDout_4__3__7 ;
    output FilterDout_4__3__6 ;
    output FilterDout_4__3__5 ;
    output FilterDout_4__3__4 ;
    output FilterDout_4__3__3 ;
    output FilterDout_4__3__2 ;
    output FilterDout_4__3__1 ;
    output FilterDout_4__3__0 ;
    output FilterDout_4__4__7 ;
    output FilterDout_4__4__6 ;
    output FilterDout_4__4__5 ;
    output FilterDout_4__4__4 ;
    output FilterDout_4__4__3 ;
    output FilterDout_4__4__2 ;
    output FilterDout_4__4__1 ;
    output FilterDout_4__4__0 ;
    output WindowDout_0__0__7 ;
    output WindowDout_0__0__6 ;
    output WindowDout_0__0__5 ;
    output WindowDout_0__0__4 ;
    output WindowDout_0__0__3 ;
    output WindowDout_0__0__2 ;
    output WindowDout_0__0__1 ;
    output WindowDout_0__0__0 ;
    output WindowDout_0__1__7 ;
    output WindowDout_0__1__6 ;
    output WindowDout_0__1__5 ;
    output WindowDout_0__1__4 ;
    output WindowDout_0__1__3 ;
    output WindowDout_0__1__2 ;
    output WindowDout_0__1__1 ;
    output WindowDout_0__1__0 ;
    output WindowDout_0__2__7 ;
    output WindowDout_0__2__6 ;
    output WindowDout_0__2__5 ;
    output WindowDout_0__2__4 ;
    output WindowDout_0__2__3 ;
    output WindowDout_0__2__2 ;
    output WindowDout_0__2__1 ;
    output WindowDout_0__2__0 ;
    output WindowDout_0__3__7 ;
    output WindowDout_0__3__6 ;
    output WindowDout_0__3__5 ;
    output WindowDout_0__3__4 ;
    output WindowDout_0__3__3 ;
    output WindowDout_0__3__2 ;
    output WindowDout_0__3__1 ;
    output WindowDout_0__3__0 ;
    output WindowDout_0__4__7 ;
    output WindowDout_0__4__6 ;
    output WindowDout_0__4__5 ;
    output WindowDout_0__4__4 ;
    output WindowDout_0__4__3 ;
    output WindowDout_0__4__2 ;
    output WindowDout_0__4__1 ;
    output WindowDout_0__4__0 ;
    output WindowDout_1__0__7 ;
    output WindowDout_1__0__6 ;
    output WindowDout_1__0__5 ;
    output WindowDout_1__0__4 ;
    output WindowDout_1__0__3 ;
    output WindowDout_1__0__2 ;
    output WindowDout_1__0__1 ;
    output WindowDout_1__0__0 ;
    output WindowDout_1__1__7 ;
    output WindowDout_1__1__6 ;
    output WindowDout_1__1__5 ;
    output WindowDout_1__1__4 ;
    output WindowDout_1__1__3 ;
    output WindowDout_1__1__2 ;
    output WindowDout_1__1__1 ;
    output WindowDout_1__1__0 ;
    output WindowDout_1__2__7 ;
    output WindowDout_1__2__6 ;
    output WindowDout_1__2__5 ;
    output WindowDout_1__2__4 ;
    output WindowDout_1__2__3 ;
    output WindowDout_1__2__2 ;
    output WindowDout_1__2__1 ;
    output WindowDout_1__2__0 ;
    output WindowDout_1__3__7 ;
    output WindowDout_1__3__6 ;
    output WindowDout_1__3__5 ;
    output WindowDout_1__3__4 ;
    output WindowDout_1__3__3 ;
    output WindowDout_1__3__2 ;
    output WindowDout_1__3__1 ;
    output WindowDout_1__3__0 ;
    output WindowDout_1__4__7 ;
    output WindowDout_1__4__6 ;
    output WindowDout_1__4__5 ;
    output WindowDout_1__4__4 ;
    output WindowDout_1__4__3 ;
    output WindowDout_1__4__2 ;
    output WindowDout_1__4__1 ;
    output WindowDout_1__4__0 ;
    output WindowDout_2__0__7 ;
    output WindowDout_2__0__6 ;
    output WindowDout_2__0__5 ;
    output WindowDout_2__0__4 ;
    output WindowDout_2__0__3 ;
    output WindowDout_2__0__2 ;
    output WindowDout_2__0__1 ;
    output WindowDout_2__0__0 ;
    output WindowDout_2__1__7 ;
    output WindowDout_2__1__6 ;
    output WindowDout_2__1__5 ;
    output WindowDout_2__1__4 ;
    output WindowDout_2__1__3 ;
    output WindowDout_2__1__2 ;
    output WindowDout_2__1__1 ;
    output WindowDout_2__1__0 ;
    output WindowDout_2__2__7 ;
    output WindowDout_2__2__6 ;
    output WindowDout_2__2__5 ;
    output WindowDout_2__2__4 ;
    output WindowDout_2__2__3 ;
    output WindowDout_2__2__2 ;
    output WindowDout_2__2__1 ;
    output WindowDout_2__2__0 ;
    output WindowDout_2__3__7 ;
    output WindowDout_2__3__6 ;
    output WindowDout_2__3__5 ;
    output WindowDout_2__3__4 ;
    output WindowDout_2__3__3 ;
    output WindowDout_2__3__2 ;
    output WindowDout_2__3__1 ;
    output WindowDout_2__3__0 ;
    output WindowDout_2__4__7 ;
    output WindowDout_2__4__6 ;
    output WindowDout_2__4__5 ;
    output WindowDout_2__4__4 ;
    output WindowDout_2__4__3 ;
    output WindowDout_2__4__2 ;
    output WindowDout_2__4__1 ;
    output WindowDout_2__4__0 ;
    output WindowDout_3__0__7 ;
    output WindowDout_3__0__6 ;
    output WindowDout_3__0__5 ;
    output WindowDout_3__0__4 ;
    output WindowDout_3__0__3 ;
    output WindowDout_3__0__2 ;
    output WindowDout_3__0__1 ;
    output WindowDout_3__0__0 ;
    output WindowDout_3__1__7 ;
    output WindowDout_3__1__6 ;
    output WindowDout_3__1__5 ;
    output WindowDout_3__1__4 ;
    output WindowDout_3__1__3 ;
    output WindowDout_3__1__2 ;
    output WindowDout_3__1__1 ;
    output WindowDout_3__1__0 ;
    output WindowDout_3__2__7 ;
    output WindowDout_3__2__6 ;
    output WindowDout_3__2__5 ;
    output WindowDout_3__2__4 ;
    output WindowDout_3__2__3 ;
    output WindowDout_3__2__2 ;
    output WindowDout_3__2__1 ;
    output WindowDout_3__2__0 ;
    output WindowDout_3__3__7 ;
    output WindowDout_3__3__6 ;
    output WindowDout_3__3__5 ;
    output WindowDout_3__3__4 ;
    output WindowDout_3__3__3 ;
    output WindowDout_3__3__2 ;
    output WindowDout_3__3__1 ;
    output WindowDout_3__3__0 ;
    output WindowDout_3__4__7 ;
    output WindowDout_3__4__6 ;
    output WindowDout_3__4__5 ;
    output WindowDout_3__4__4 ;
    output WindowDout_3__4__3 ;
    output WindowDout_3__4__2 ;
    output WindowDout_3__4__1 ;
    output WindowDout_3__4__0 ;
    output WindowDout_4__0__7 ;
    output WindowDout_4__0__6 ;
    output WindowDout_4__0__5 ;
    output WindowDout_4__0__4 ;
    output WindowDout_4__0__3 ;
    output WindowDout_4__0__2 ;
    output WindowDout_4__0__1 ;
    output WindowDout_4__0__0 ;
    output WindowDout_4__1__7 ;
    output WindowDout_4__1__6 ;
    output WindowDout_4__1__5 ;
    output WindowDout_4__1__4 ;
    output WindowDout_4__1__3 ;
    output WindowDout_4__1__2 ;
    output WindowDout_4__1__1 ;
    output WindowDout_4__1__0 ;
    output WindowDout_4__2__7 ;
    output WindowDout_4__2__6 ;
    output WindowDout_4__2__5 ;
    output WindowDout_4__2__4 ;
    output WindowDout_4__2__3 ;
    output WindowDout_4__2__2 ;
    output WindowDout_4__2__1 ;
    output WindowDout_4__2__0 ;
    output WindowDout_4__3__7 ;
    output WindowDout_4__3__6 ;
    output WindowDout_4__3__5 ;
    output WindowDout_4__3__4 ;
    output WindowDout_4__3__3 ;
    output WindowDout_4__3__2 ;
    output WindowDout_4__3__1 ;
    output WindowDout_4__3__0 ;
    output WindowDout_4__4__7 ;
    output WindowDout_4__4__6 ;
    output WindowDout_4__4__5 ;
    output WindowDout_4__4__4 ;
    output WindowDout_4__4__3 ;
    output WindowDout_4__4__2 ;
    output WindowDout_4__4__1 ;
    output WindowDout_4__4__0 ;

    wire FilterEN_4__4, WindowEN_4__4, nx941, EN_dup_1411, EN_dup_1279, 
         EN_dup_1147, EN_dup_1081, EN_dup_1015, EN, nx955, EN_dup_1422, 
         EN_dup_1290, EN_dup_1158, EN_dup_1092, EN_dup_1026, EN_dup_1004, 
         L0_0_L1_0_Fij_nx212, L0_0_L1_0_Fij_nx222, L0_0_L1_0_Fij_nx232, 
         L0_0_L1_0_Fij_nx242, L0_0_L1_0_Fij_nx252, L0_0_L1_0_Fij_nx262, 
         L0_0_L1_0_Fij_nx272, L0_0_L1_0_Fij_nx282, L0_0_L1_0_Fij_nx296, 
         L0_0_L1_0_Fij_nx331, L0_0_L1_0_Fij_nx333, L0_0_L1_0_Wij_nx212, 
         L0_0_L1_0_Wij_nx222, L0_0_L1_0_Wij_nx232, L0_0_L1_0_Wij_nx242, 
         L0_0_L1_0_Wij_nx252, L0_0_L1_0_Wij_nx262, L0_0_L1_0_Wij_nx272, 
         L0_0_L1_0_Wij_nx282, L0_0_L1_0_Wij_nx296, L0_0_L1_0_Wij_nx331, 
         L0_0_L1_0_Wij_nx333, L0_0_L1_1_Fij_nx212, L0_0_L1_1_Fij_nx222, 
         L0_0_L1_1_Fij_nx232, L0_0_L1_1_Fij_nx242, L0_0_L1_1_Fij_nx252, 
         L0_0_L1_1_Fij_nx262, L0_0_L1_1_Fij_nx272, L0_0_L1_1_Fij_nx282, 
         L0_0_L1_1_Fij_nx296, L0_0_L1_1_Fij_nx331, L0_0_L1_1_Fij_nx333, 
         L0_0_L1_1_Wij_nx212, L0_0_L1_1_Wij_nx222, L0_0_L1_1_Wij_nx232, 
         L0_0_L1_1_Wij_nx242, L0_0_L1_1_Wij_nx252, L0_0_L1_1_Wij_nx262, 
         L0_0_L1_1_Wij_nx272, L0_0_L1_1_Wij_nx282, L0_0_L1_1_Wij_nx296, 
         L0_0_L1_1_Wij_nx331, L0_0_L1_1_Wij_nx333, L0_0_L1_2_Fij_nx212, 
         L0_0_L1_2_Fij_nx222, L0_0_L1_2_Fij_nx232, L0_0_L1_2_Fij_nx242, 
         L0_0_L1_2_Fij_nx252, L0_0_L1_2_Fij_nx262, L0_0_L1_2_Fij_nx272, 
         L0_0_L1_2_Fij_nx282, L0_0_L1_2_Fij_nx296, L0_0_L1_2_Fij_nx331, 
         L0_0_L1_2_Fij_nx333, L0_0_L1_2_Wij_nx212, L0_0_L1_2_Wij_nx222, 
         L0_0_L1_2_Wij_nx232, L0_0_L1_2_Wij_nx242, L0_0_L1_2_Wij_nx252, 
         L0_0_L1_2_Wij_nx262, L0_0_L1_2_Wij_nx272, L0_0_L1_2_Wij_nx282, 
         L0_0_L1_2_Wij_nx296, L0_0_L1_2_Wij_nx331, L0_0_L1_2_Wij_nx333, 
         L0_0_L1_3_Fij_nx212, L0_0_L1_3_Fij_nx222, L0_0_L1_3_Fij_nx232, 
         L0_0_L1_3_Fij_nx242, L0_0_L1_3_Fij_nx252, L0_0_L1_3_Fij_nx262, 
         L0_0_L1_3_Fij_nx272, L0_0_L1_3_Fij_nx282, L0_0_L1_3_Fij_nx296, 
         L0_0_L1_3_Fij_nx331, L0_0_L1_3_Fij_nx333, L0_0_L1_3_Wij_nx212, 
         L0_0_L1_3_Wij_nx222, L0_0_L1_3_Wij_nx232, L0_0_L1_3_Wij_nx242, 
         L0_0_L1_3_Wij_nx252, L0_0_L1_3_Wij_nx262, L0_0_L1_3_Wij_nx272, 
         L0_0_L1_3_Wij_nx282, L0_0_L1_3_Wij_nx296, L0_0_L1_3_Wij_nx331, 
         L0_0_L1_3_Wij_nx333, L0_0_L1_4_Fij_nx212, L0_0_L1_4_Fij_nx222, 
         L0_0_L1_4_Fij_nx232, L0_0_L1_4_Fij_nx242, L0_0_L1_4_Fij_nx252, 
         L0_0_L1_4_Fij_nx262, L0_0_L1_4_Fij_nx272, L0_0_L1_4_Fij_nx282, 
         L0_0_L1_4_Fij_nx296, L0_0_L1_4_Fij_nx331, L0_0_L1_4_Fij_nx333, 
         L0_0_L1_4_Wij_nx212, L0_0_L1_4_Wij_nx222, L0_0_L1_4_Wij_nx232, 
         L0_0_L1_4_Wij_nx242, L0_0_L1_4_Wij_nx252, L0_0_L1_4_Wij_nx262, 
         L0_0_L1_4_Wij_nx272, L0_0_L1_4_Wij_nx282, L0_0_L1_4_Wij_nx296, 
         L0_0_L1_4_Wij_nx331, L0_0_L1_4_Wij_nx333, L0_1_L1_0_Fij_nx212, 
         L0_1_L1_0_Fij_nx222, L0_1_L1_0_Fij_nx232, L0_1_L1_0_Fij_nx242, 
         L0_1_L1_0_Fij_nx252, L0_1_L1_0_Fij_nx262, L0_1_L1_0_Fij_nx272, 
         L0_1_L1_0_Fij_nx282, L0_1_L1_0_Fij_nx296, L0_1_L1_0_Fij_nx331, 
         L0_1_L1_0_Fij_nx333, L0_1_L1_0_Wij_nx212, L0_1_L1_0_Wij_nx222, 
         L0_1_L1_0_Wij_nx232, L0_1_L1_0_Wij_nx242, L0_1_L1_0_Wij_nx252, 
         L0_1_L1_0_Wij_nx262, L0_1_L1_0_Wij_nx272, L0_1_L1_0_Wij_nx282, 
         L0_1_L1_0_Wij_nx296, L0_1_L1_0_Wij_nx331, L0_1_L1_0_Wij_nx333, 
         L0_1_L1_1_Fij_nx212, L0_1_L1_1_Fij_nx222, L0_1_L1_1_Fij_nx232, 
         L0_1_L1_1_Fij_nx242, L0_1_L1_1_Fij_nx252, L0_1_L1_1_Fij_nx262, 
         L0_1_L1_1_Fij_nx272, L0_1_L1_1_Fij_nx282, L0_1_L1_1_Fij_nx296, 
         L0_1_L1_1_Fij_nx331, L0_1_L1_1_Fij_nx333, L0_1_L1_1_Wij_nx212, 
         L0_1_L1_1_Wij_nx222, L0_1_L1_1_Wij_nx232, L0_1_L1_1_Wij_nx242, 
         L0_1_L1_1_Wij_nx252, L0_1_L1_1_Wij_nx262, L0_1_L1_1_Wij_nx272, 
         L0_1_L1_1_Wij_nx282, L0_1_L1_1_Wij_nx296, L0_1_L1_1_Wij_nx331, 
         L0_1_L1_1_Wij_nx333, L0_1_L1_2_Fij_nx212, L0_1_L1_2_Fij_nx222, 
         L0_1_L1_2_Fij_nx232, L0_1_L1_2_Fij_nx242, L0_1_L1_2_Fij_nx252, 
         L0_1_L1_2_Fij_nx262, L0_1_L1_2_Fij_nx272, L0_1_L1_2_Fij_nx282, 
         L0_1_L1_2_Fij_nx296, L0_1_L1_2_Fij_nx331, L0_1_L1_2_Fij_nx333, 
         L0_1_L1_2_Wij_nx212, L0_1_L1_2_Wij_nx222, L0_1_L1_2_Wij_nx232, 
         L0_1_L1_2_Wij_nx242, L0_1_L1_2_Wij_nx252, L0_1_L1_2_Wij_nx262, 
         L0_1_L1_2_Wij_nx272, L0_1_L1_2_Wij_nx282, L0_1_L1_2_Wij_nx296, 
         L0_1_L1_2_Wij_nx331, L0_1_L1_2_Wij_nx333, L0_1_L1_3_Fij_nx212, 
         L0_1_L1_3_Fij_nx222, L0_1_L1_3_Fij_nx232, L0_1_L1_3_Fij_nx242, 
         L0_1_L1_3_Fij_nx252, L0_1_L1_3_Fij_nx262, L0_1_L1_3_Fij_nx272, 
         L0_1_L1_3_Fij_nx282, L0_1_L1_3_Fij_nx296, L0_1_L1_3_Fij_nx331, 
         L0_1_L1_3_Fij_nx333, L0_1_L1_3_Wij_nx212, L0_1_L1_3_Wij_nx222, 
         L0_1_L1_3_Wij_nx232, L0_1_L1_3_Wij_nx242, L0_1_L1_3_Wij_nx252, 
         L0_1_L1_3_Wij_nx262, L0_1_L1_3_Wij_nx272, L0_1_L1_3_Wij_nx282, 
         L0_1_L1_3_Wij_nx296, L0_1_L1_3_Wij_nx331, L0_1_L1_3_Wij_nx333, 
         L0_1_L1_4_Fij_nx212, L0_1_L1_4_Fij_nx222, L0_1_L1_4_Fij_nx232, 
         L0_1_L1_4_Fij_nx242, L0_1_L1_4_Fij_nx252, L0_1_L1_4_Fij_nx262, 
         L0_1_L1_4_Fij_nx272, L0_1_L1_4_Fij_nx282, L0_1_L1_4_Fij_nx296, 
         L0_1_L1_4_Fij_nx331, L0_1_L1_4_Fij_nx333, L0_1_L1_4_Wij_nx212, 
         L0_1_L1_4_Wij_nx222, L0_1_L1_4_Wij_nx232, L0_1_L1_4_Wij_nx242, 
         L0_1_L1_4_Wij_nx252, L0_1_L1_4_Wij_nx262, L0_1_L1_4_Wij_nx272, 
         L0_1_L1_4_Wij_nx282, L0_1_L1_4_Wij_nx296, L0_1_L1_4_Wij_nx331, 
         L0_1_L1_4_Wij_nx333, L0_2_L1_0_Fij_nx212, L0_2_L1_0_Fij_nx222, 
         L0_2_L1_0_Fij_nx232, L0_2_L1_0_Fij_nx242, L0_2_L1_0_Fij_nx252, 
         L0_2_L1_0_Fij_nx262, L0_2_L1_0_Fij_nx272, L0_2_L1_0_Fij_nx282, 
         L0_2_L1_0_Fij_nx296, L0_2_L1_0_Fij_nx331, L0_2_L1_0_Fij_nx333, 
         L0_2_L1_0_Wij_nx212, L0_2_L1_0_Wij_nx222, L0_2_L1_0_Wij_nx232, 
         L0_2_L1_0_Wij_nx242, L0_2_L1_0_Wij_nx252, L0_2_L1_0_Wij_nx262, 
         L0_2_L1_0_Wij_nx272, L0_2_L1_0_Wij_nx282, L0_2_L1_0_Wij_nx296, 
         L0_2_L1_0_Wij_nx331, L0_2_L1_0_Wij_nx333, L0_2_L1_1_Fij_nx212, 
         L0_2_L1_1_Fij_nx222, L0_2_L1_1_Fij_nx232, L0_2_L1_1_Fij_nx242, 
         L0_2_L1_1_Fij_nx252, L0_2_L1_1_Fij_nx262, L0_2_L1_1_Fij_nx272, 
         L0_2_L1_1_Fij_nx282, L0_2_L1_1_Fij_nx296, L0_2_L1_1_Fij_nx331, 
         L0_2_L1_1_Fij_nx333, L0_2_L1_1_Wij_nx212, L0_2_L1_1_Wij_nx222, 
         L0_2_L1_1_Wij_nx232, L0_2_L1_1_Wij_nx242, L0_2_L1_1_Wij_nx252, 
         L0_2_L1_1_Wij_nx262, L0_2_L1_1_Wij_nx272, L0_2_L1_1_Wij_nx282, 
         L0_2_L1_1_Wij_nx296, L0_2_L1_1_Wij_nx331, L0_2_L1_1_Wij_nx333, 
         L0_2_L1_2_Fij_nx212, L0_2_L1_2_Fij_nx222, L0_2_L1_2_Fij_nx232, 
         L0_2_L1_2_Fij_nx242, L0_2_L1_2_Fij_nx252, L0_2_L1_2_Fij_nx262, 
         L0_2_L1_2_Fij_nx272, L0_2_L1_2_Fij_nx282, L0_2_L1_2_Fij_nx296, 
         L0_2_L1_2_Fij_nx331, L0_2_L1_2_Fij_nx333, L0_2_L1_2_Wij_nx212, 
         L0_2_L1_2_Wij_nx222, L0_2_L1_2_Wij_nx232, L0_2_L1_2_Wij_nx242, 
         L0_2_L1_2_Wij_nx252, L0_2_L1_2_Wij_nx262, L0_2_L1_2_Wij_nx272, 
         L0_2_L1_2_Wij_nx282, L0_2_L1_2_Wij_nx296, L0_2_L1_2_Wij_nx331, 
         L0_2_L1_2_Wij_nx333, L0_2_L1_3_Fij_nx212, L0_2_L1_3_Fij_nx222, 
         L0_2_L1_3_Fij_nx232, L0_2_L1_3_Fij_nx242, L0_2_L1_3_Fij_nx252, 
         L0_2_L1_3_Fij_nx262, L0_2_L1_3_Fij_nx272, L0_2_L1_3_Fij_nx282, 
         L0_2_L1_3_Fij_nx296, L0_2_L1_3_Fij_nx331, L0_2_L1_3_Fij_nx333, 
         L0_2_L1_3_Wij_nx212, L0_2_L1_3_Wij_nx222, L0_2_L1_3_Wij_nx232, 
         L0_2_L1_3_Wij_nx242, L0_2_L1_3_Wij_nx252, L0_2_L1_3_Wij_nx262, 
         L0_2_L1_3_Wij_nx272, L0_2_L1_3_Wij_nx282, L0_2_L1_3_Wij_nx296, 
         L0_2_L1_3_Wij_nx331, L0_2_L1_3_Wij_nx333, L0_2_L1_4_Fij_nx212, 
         L0_2_L1_4_Fij_nx222, L0_2_L1_4_Fij_nx232, L0_2_L1_4_Fij_nx242, 
         L0_2_L1_4_Fij_nx252, L0_2_L1_4_Fij_nx262, L0_2_L1_4_Fij_nx272, 
         L0_2_L1_4_Fij_nx282, L0_2_L1_4_Fij_nx296, L0_2_L1_4_Fij_nx331, 
         L0_2_L1_4_Fij_nx333, L0_2_L1_4_Wij_nx212, L0_2_L1_4_Wij_nx222, 
         L0_2_L1_4_Wij_nx232, L0_2_L1_4_Wij_nx242, L0_2_L1_4_Wij_nx252, 
         L0_2_L1_4_Wij_nx262, L0_2_L1_4_Wij_nx272, L0_2_L1_4_Wij_nx282, 
         L0_2_L1_4_Wij_nx296, L0_2_L1_4_Wij_nx331, L0_2_L1_4_Wij_nx333, 
         L0_3_L1_0_Fij_nx212, L0_3_L1_0_Fij_nx222, L0_3_L1_0_Fij_nx232, 
         L0_3_L1_0_Fij_nx242, L0_3_L1_0_Fij_nx252, L0_3_L1_0_Fij_nx262, 
         L0_3_L1_0_Fij_nx272, L0_3_L1_0_Fij_nx282, L0_3_L1_0_Fij_nx296, 
         L0_3_L1_0_Fij_nx331, L0_3_L1_0_Fij_nx333, L0_3_L1_0_Wij_nx212, 
         L0_3_L1_0_Wij_nx222, L0_3_L1_0_Wij_nx232, L0_3_L1_0_Wij_nx242, 
         L0_3_L1_0_Wij_nx252, L0_3_L1_0_Wij_nx262, L0_3_L1_0_Wij_nx272, 
         L0_3_L1_0_Wij_nx282, L0_3_L1_0_Wij_nx296, L0_3_L1_0_Wij_nx331, 
         L0_3_L1_0_Wij_nx333, L0_3_L1_1_Fij_nx212, L0_3_L1_1_Fij_nx222, 
         L0_3_L1_1_Fij_nx232, L0_3_L1_1_Fij_nx242, L0_3_L1_1_Fij_nx252, 
         L0_3_L1_1_Fij_nx262, L0_3_L1_1_Fij_nx272, L0_3_L1_1_Fij_nx282, 
         L0_3_L1_1_Fij_nx296, L0_3_L1_1_Fij_nx331, L0_3_L1_1_Fij_nx333, 
         L0_3_L1_1_Wij_nx212, L0_3_L1_1_Wij_nx222, L0_3_L1_1_Wij_nx232, 
         L0_3_L1_1_Wij_nx242, L0_3_L1_1_Wij_nx252, L0_3_L1_1_Wij_nx262, 
         L0_3_L1_1_Wij_nx272, L0_3_L1_1_Wij_nx282, L0_3_L1_1_Wij_nx296, 
         L0_3_L1_1_Wij_nx331, L0_3_L1_1_Wij_nx333, L0_3_L1_2_Fij_nx212, 
         L0_3_L1_2_Fij_nx222, L0_3_L1_2_Fij_nx232, L0_3_L1_2_Fij_nx242, 
         L0_3_L1_2_Fij_nx252, L0_3_L1_2_Fij_nx262, L0_3_L1_2_Fij_nx272, 
         L0_3_L1_2_Fij_nx282, L0_3_L1_2_Fij_nx296, L0_3_L1_2_Fij_nx331, 
         L0_3_L1_2_Fij_nx333, L0_3_L1_2_Wij_nx212, L0_3_L1_2_Wij_nx222, 
         L0_3_L1_2_Wij_nx232, L0_3_L1_2_Wij_nx242, L0_3_L1_2_Wij_nx252, 
         L0_3_L1_2_Wij_nx262, L0_3_L1_2_Wij_nx272, L0_3_L1_2_Wij_nx282, 
         L0_3_L1_2_Wij_nx296, L0_3_L1_2_Wij_nx331, L0_3_L1_2_Wij_nx333, 
         L0_3_L1_3_Fij_nx212, L0_3_L1_3_Fij_nx222, L0_3_L1_3_Fij_nx232, 
         L0_3_L1_3_Fij_nx242, L0_3_L1_3_Fij_nx252, L0_3_L1_3_Fij_nx262, 
         L0_3_L1_3_Fij_nx272, L0_3_L1_3_Fij_nx282, L0_3_L1_3_Fij_nx296, 
         L0_3_L1_3_Fij_nx331, L0_3_L1_3_Fij_nx333, L0_3_L1_3_Wij_nx212, 
         L0_3_L1_3_Wij_nx222, L0_3_L1_3_Wij_nx232, L0_3_L1_3_Wij_nx242, 
         L0_3_L1_3_Wij_nx252, L0_3_L1_3_Wij_nx262, L0_3_L1_3_Wij_nx272, 
         L0_3_L1_3_Wij_nx282, L0_3_L1_3_Wij_nx296, L0_3_L1_3_Wij_nx331, 
         L0_3_L1_3_Wij_nx333, L0_3_L1_4_Fij_nx212, L0_3_L1_4_Fij_nx222, 
         L0_3_L1_4_Fij_nx232, L0_3_L1_4_Fij_nx242, L0_3_L1_4_Fij_nx252, 
         L0_3_L1_4_Fij_nx262, L0_3_L1_4_Fij_nx272, L0_3_L1_4_Fij_nx282, 
         L0_3_L1_4_Fij_nx296, L0_3_L1_4_Fij_nx331, L0_3_L1_4_Fij_nx333, 
         L0_3_L1_4_Wij_nx212, L0_3_L1_4_Wij_nx222, L0_3_L1_4_Wij_nx232, 
         L0_3_L1_4_Wij_nx242, L0_3_L1_4_Wij_nx252, L0_3_L1_4_Wij_nx262, 
         L0_3_L1_4_Wij_nx272, L0_3_L1_4_Wij_nx282, L0_3_L1_4_Wij_nx296, 
         L0_3_L1_4_Wij_nx331, L0_3_L1_4_Wij_nx333, L0_4_L1_0_Fij_nx212, 
         L0_4_L1_0_Fij_nx222, L0_4_L1_0_Fij_nx232, L0_4_L1_0_Fij_nx242, 
         L0_4_L1_0_Fij_nx252, L0_4_L1_0_Fij_nx262, L0_4_L1_0_Fij_nx272, 
         L0_4_L1_0_Fij_nx282, L0_4_L1_0_Fij_nx296, L0_4_L1_0_Fij_nx331, 
         L0_4_L1_0_Fij_nx333, L0_4_L1_0_Wij_nx212, L0_4_L1_0_Wij_nx222, 
         L0_4_L1_0_Wij_nx232, L0_4_L1_0_Wij_nx242, L0_4_L1_0_Wij_nx252, 
         L0_4_L1_0_Wij_nx262, L0_4_L1_0_Wij_nx272, L0_4_L1_0_Wij_nx282, 
         L0_4_L1_0_Wij_nx296, L0_4_L1_0_Wij_nx331, L0_4_L1_0_Wij_nx333, 
         L0_4_L1_1_Fij_nx212, L0_4_L1_1_Fij_nx222, L0_4_L1_1_Fij_nx232, 
         L0_4_L1_1_Fij_nx242, L0_4_L1_1_Fij_nx252, L0_4_L1_1_Fij_nx262, 
         L0_4_L1_1_Fij_nx272, L0_4_L1_1_Fij_nx282, L0_4_L1_1_Fij_nx296, 
         L0_4_L1_1_Fij_nx331, L0_4_L1_1_Fij_nx333, L0_4_L1_1_Wij_nx212, 
         L0_4_L1_1_Wij_nx222, L0_4_L1_1_Wij_nx232, L0_4_L1_1_Wij_nx242, 
         L0_4_L1_1_Wij_nx252, L0_4_L1_1_Wij_nx262, L0_4_L1_1_Wij_nx272, 
         L0_4_L1_1_Wij_nx282, L0_4_L1_1_Wij_nx296, L0_4_L1_1_Wij_nx331, 
         L0_4_L1_1_Wij_nx333, L0_4_L1_2_Fij_nx212, L0_4_L1_2_Fij_nx222, 
         L0_4_L1_2_Fij_nx232, L0_4_L1_2_Fij_nx242, L0_4_L1_2_Fij_nx252, 
         L0_4_L1_2_Fij_nx262, L0_4_L1_2_Fij_nx272, L0_4_L1_2_Fij_nx282, 
         L0_4_L1_2_Fij_nx296, L0_4_L1_2_Fij_nx331, L0_4_L1_2_Fij_nx333, 
         L0_4_L1_2_Wij_nx212, L0_4_L1_2_Wij_nx222, L0_4_L1_2_Wij_nx232, 
         L0_4_L1_2_Wij_nx242, L0_4_L1_2_Wij_nx252, L0_4_L1_2_Wij_nx262, 
         L0_4_L1_2_Wij_nx272, L0_4_L1_2_Wij_nx282, L0_4_L1_2_Wij_nx296, 
         L0_4_L1_2_Wij_nx331, L0_4_L1_2_Wij_nx333, L0_4_L1_3_Fij_nx212, 
         L0_4_L1_3_Fij_nx222, L0_4_L1_3_Fij_nx232, L0_4_L1_3_Fij_nx242, 
         L0_4_L1_3_Fij_nx252, L0_4_L1_3_Fij_nx262, L0_4_L1_3_Fij_nx272, 
         L0_4_L1_3_Fij_nx282, L0_4_L1_3_Fij_nx296, L0_4_L1_3_Fij_nx331, 
         L0_4_L1_3_Fij_nx333, L0_4_L1_3_Wij_nx212, L0_4_L1_3_Wij_nx222, 
         L0_4_L1_3_Wij_nx232, L0_4_L1_3_Wij_nx242, L0_4_L1_3_Wij_nx252, 
         L0_4_L1_3_Wij_nx262, L0_4_L1_3_Wij_nx272, L0_4_L1_3_Wij_nx282, 
         L0_4_L1_3_Wij_nx296, L0_4_L1_3_Wij_nx331, L0_4_L1_3_Wij_nx333, 
         L0_4_L1_4_Fij_nx212, L0_4_L1_4_Fij_nx222, L0_4_L1_4_Fij_nx232, 
         L0_4_L1_4_Fij_nx242, L0_4_L1_4_Fij_nx252, L0_4_L1_4_Fij_nx262, 
         L0_4_L1_4_Fij_nx272, L0_4_L1_4_Fij_nx282, L0_4_L1_4_Fij_nx296, 
         L0_4_L1_4_Fij_nx331, L0_4_L1_4_Fij_nx333, L0_4_L1_4_Wij_nx212, 
         L0_4_L1_4_Wij_nx222, L0_4_L1_4_Wij_nx232, L0_4_L1_4_Wij_nx242, 
         L0_4_L1_4_Wij_nx252, L0_4_L1_4_Wij_nx262, L0_4_L1_4_Wij_nx272, 
         L0_4_L1_4_Wij_nx282, L0_4_L1_4_Wij_nx296, L0_4_L1_4_Wij_nx331, 
         L0_4_L1_4_Wij_nx333, nx1576, nx1578, nx1580, nx1584, nx1586, nx1588, 
         nx1590, nx1592, nx1594, nx1596, nx1598, nx1600, nx1602, nx1604, nx1606, 
         nx1608, nx1610, nx1612, nx1614, nx1616, nx1618, nx1622, nx1624, nx1626, 
         nx1628, nx1630, nx1632, nx1634, nx1636, nx1638, nx1640, nx1642, nx1644, 
         nx1646, nx1648, nx1650, nx1652, nx1654, nx1656, nx1660, nx1662, nx1664, 
         nx1666, nx1668, nx1670, nx1672, nx1674, nx1676, nx1678, nx1680, nx1682, 
         nx1684, nx1686, nx1688, nx1690, nx1692, nx1694, nx1698, nx1700, nx1702, 
         nx1704, nx1706, nx1708, nx1710, nx1712, nx1714, nx1716, nx1718, nx1720, 
         nx1722, nx1724, nx1726, nx1728, nx1730, nx1732, nx1736, nx1738, nx1740, 
         nx1742, nx1744, nx1746, nx1748, nx1750, nx1752, nx1754, nx1756, nx1758, 
         nx1760, nx1762, nx1764, nx1766, nx1768, nx1770, nx1774, nx1776, nx1778, 
         nx1780, nx1782, nx1784, nx1786, nx1788, nx1790, nx1792, nx1794, nx1796, 
         nx1798, nx1800, nx1802, nx1804, nx1806, nx1808, nx1812, nx1814, nx1816, 
         nx1818, nx1820, nx1822, nx1824, nx1826, nx1828, nx1830, nx1832, nx1834, 
         nx1836, nx1838, nx1840, nx1842, nx1844, nx1846, nx1850, nx1852, nx1854, 
         nx1856, nx1858, nx1860, nx1862, nx1864, nx1866, nx1868, nx1870, nx1872, 
         nx1874, nx1876, nx1878, nx1880, nx1882, nx1884, nx1888, nx1890, nx1892, 
         nx1894, nx1896, nx1898, nx1900, nx1902, nx1904, nx1906, nx1908, nx1910, 
         nx1912, nx1914, nx1916, nx1918, nx1920, nx1922, nx1926, nx1928, nx1930, 
         nx1932, nx1934, nx1936, nx1938, nx1940, nx1942, nx1944, nx1946, nx1948, 
         nx1950, nx1952, nx1954, nx1956, nx1958, nx1962, nx1964, nx1966, nx1968, 
         nx1970, nx1972, nx1974, nx1976, nx1978, nx1980, nx1984, nx1986, nx1988, 
         nx1990, nx1992, nx1994, nx1996, nx1998, nx2000, nx2002, nx2006, nx2008, 
         nx2010, nx2012, nx2014, nx2016, nx2018, nx2020, nx2022, nx2024, nx2028, 
         nx2030, nx2032, nx2034, nx2036, nx2038, nx2040, nx2042, nx2044, nx2046, 
         nx2050, nx2052, nx2054, nx2056, nx2058, nx2060, nx2062, nx2064, nx2066, 
         nx2068, nx2072, nx2074, nx2076, nx2078, nx2080, nx2082, nx2084, nx2086, 
         nx2088, nx2090, nx2094, nx2096, nx2098, nx2100, nx2102, nx2104, nx2106, 
         nx2108, nx2110, nx2112, nx2116, nx2118, nx2120, nx2122, nx2124, nx2126, 
         nx2128, nx2130, nx2132, nx2134, nx2138, nx2140, nx2142, nx2144, nx2146, 
         nx2148, nx2150, nx2152, nx2154, nx2156, nx2160, nx2162, nx2164, nx2166, 
         nx2168, nx2170, nx2172, nx2174, nx2176, nx2178, nx2182, nx2184, nx2186, 
         nx2188, nx2190, nx2192, nx2194, nx2196, nx2198, nx2200, nx2204, nx2206, 
         nx2208, nx2210, nx2212, nx2214, nx2216, nx2218, nx2220, nx2222, nx2226, 
         nx2228, nx2230, nx2232, nx2234, nx2236, nx2238, nx2240, nx2242, nx2244, 
         nx2248, nx2250, nx2252, nx2254, nx2256, nx2258, nx2260, nx2262, nx2264, 
         nx2266, nx2270, nx2272, nx2274, nx2276, nx2278, nx2280, nx2282, nx2284, 
         nx2286, nx2288, nx2292, nx2294, nx2296, nx2298, nx2300, nx2302, nx2304, 
         nx2306, nx2308, nx2310, nx2314, nx2316, nx2318, nx2320, nx2322, nx2324, 
         nx2326, nx2328, nx2330, nx2332, nx2336, nx2338, nx2340, nx2342, nx2344, 
         nx2346, nx2348, nx2350, nx2352, nx2354, nx2358, nx2360, nx2362, nx2364, 
         nx2366, nx2368, nx2370, nx2372, nx2374, nx2376, nx2380, nx2382, nx2384, 
         nx2386, nx2388, nx2390, nx2392, nx2394, nx2396, nx2398, nx2402, nx2404, 
         nx2406, nx2408, nx2410, nx2412, nx2414, nx2416, nx2418, nx2420, nx2424, 
         nx2426, nx2428, nx2430, nx2432, nx2434, nx2436, nx2438, nx2440, nx2442, 
         nx2446, nx2448, nx2450, nx2452, nx2454, nx2456, nx2458, nx2460, nx2462, 
         nx2464, nx2468, nx2470, nx2472, nx2474, nx2476, nx2478, nx2480, nx2482, 
         nx2484, nx2486, nx2490, nx2492, nx2494, nx2496, nx2498, nx2500, nx2502, 
         nx2504, nx2506, nx2508, nx2512, nx2514, nx2516, nx2518, nx2520, nx2522, 
         nx2524, nx2526, nx2528, nx2530, nx2534, nx2536, nx2538, nx2540, nx2542, 
         nx2544, nx2546, nx2548, nx2550, nx2552, nx2556, nx2558, nx2560, nx2562, 
         nx2564, nx2566, nx2568, nx2570, nx2572, nx2574, nx2578, nx2580, nx2582, 
         nx2584, nx2586, nx2588, nx2590, nx2592, nx2594, nx2596, nx2600, nx2602, 
         nx2604, nx2606, nx2608, nx2610, nx2612, nx2614, nx2616, nx2618, nx2622, 
         nx2624, nx2626, nx2628, nx2630, nx2632, nx2634, nx2636, nx2638, nx2642, 
         nx2644, nx2646, nx2650, nx2652, nx2654, nx2656, nx2658, nx2660, nx2662, 
         nx2664, nx2666, nx2670, nx2672, nx2674, nx2678, nx2680, nx2682, nx2684, 
         nx2686, nx2688, nx2690, nx2692, nx2694, nx2698, nx2700, nx2702, nx2706, 
         nx2708, nx2710, nx2712, nx2714, nx2716, nx2718, nx2720, nx2722, nx2726, 
         nx2728, nx2730, nx2734, nx2736, nx2738, nx2740, nx2742, nx2744, nx2746, 
         nx2748, nx2750, nx2754, nx2756, nx2758, nx2760, nx2762, nx2764, nx2766, 
         nx2768, nx2770, nx2772, nx2774, nx2776, nx2778, nx2780, nx2782, nx2784, 
         nx2786, nx2788, nx2790, nx2792, nx2794, nx2796, nx2798, nx2800, nx2802, 
         nx2804, nx2806, nx2808, nx2810, nx2812, nx2814, nx2816, nx2818, nx2820, 
         nx2822, nx2824, nx2826, nx2828, nx2830, nx2832, nx2834, nx2836, nx2838, 
         nx2840, nx2842, nx2844, nx2846, nx2848, nx2850, nx2852, nx2854, nx2856, 
         nx2858, nx2860, nx2862, nx2864, nx2866, nx2868, nx2870, nx2872, nx2874, 
         nx2876, nx2878, nx2880, nx2882, nx2884, nx2886, nx2888, nx2890, nx2892, 
         nx2894, nx2896, nx2898, nx2900, nx2902, nx2904, nx2906, nx2908, nx2910, 
         nx2912, nx2914, nx2916, nx2918, nx2920, nx2922, nx2924, nx2926, nx2928, 
         nx2930, nx2932, nx2934, nx2936, nx2938, nx2940, nx2942, nx2944, nx2946, 
         nx2948, nx2950, nx2952, nx2954;
    wire [399:0] \$dummy ;




    and02 ix1 (.Y (WindowEN_4__4), .A0 (WindowWR), .A1 (FilterSize)) ;
    and02 ix3 (.Y (FilterEN_4__4), .A0 (FilterSize), .A1 (FilterWR)) ;
    inv01 ix940 (.Y (nx941), .A (FilterEN_4__4)) ;
    inv01 ix942 (.Y (EN_dup_1411), .A (nx941)) ;
    inv01 ix944 (.Y (EN_dup_1279), .A (nx941)) ;
    inv01 ix946 (.Y (EN_dup_1147), .A (nx941)) ;
    inv01 ix948 (.Y (EN_dup_1081), .A (nx941)) ;
    inv01 ix950 (.Y (EN_dup_1015), .A (nx941)) ;
    inv01 ix952 (.Y (EN), .A (nx941)) ;
    inv01 ix954 (.Y (nx955), .A (WindowEN_4__4)) ;
    inv01 ix956 (.Y (EN_dup_1422), .A (nx955)) ;
    inv01 ix958 (.Y (EN_dup_1290), .A (nx955)) ;
    inv01 ix960 (.Y (EN_dup_1158), .A (nx955)) ;
    inv01 ix962 (.Y (EN_dup_1092), .A (nx955)) ;
    inv01 ix964 (.Y (EN_dup_1026), .A (nx955)) ;
    inv01 ix966 (.Y (EN_dup_1004), .A (nx955)) ;
    dff L0_0_L1_0_Fij_reg_Dout_0 (.Q (FilterDout_0__0__0), .QB (\$dummy [0]), .D (
        L0_0_L1_0_Fij_nx212), .CLK (CLK)) ;
    nor02_2x L0_0_L1_0_Fij_ix297 (.Y (L0_0_L1_0_Fij_nx296), .A0 (RST), .A1 (
             L0_0_L1_0_Fij_nx331)) ;
    dff L0_0_L1_0_Fij_reg_Dout_1 (.Q (FilterDout_0__0__1), .QB (\$dummy [1]), .D (
        L0_0_L1_0_Fij_nx222), .CLK (CLK)) ;
    dff L0_0_L1_0_Fij_reg_Dout_2 (.Q (FilterDout_0__0__2), .QB (\$dummy [2]), .D (
        L0_0_L1_0_Fij_nx232), .CLK (CLK)) ;
    dff L0_0_L1_0_Fij_reg_Dout_3 (.Q (FilterDout_0__0__3), .QB (\$dummy [3]), .D (
        L0_0_L1_0_Fij_nx242), .CLK (CLK)) ;
    dff L0_0_L1_0_Fij_reg_Dout_4 (.Q (FilterDout_0__0__4), .QB (\$dummy [4]), .D (
        L0_0_L1_0_Fij_nx252), .CLK (CLK)) ;
    dff L0_0_L1_0_Fij_reg_Dout_5 (.Q (FilterDout_0__0__5), .QB (\$dummy [5]), .D (
        L0_0_L1_0_Fij_nx262), .CLK (CLK)) ;
    dff L0_0_L1_0_Fij_reg_Dout_6 (.Q (FilterDout_0__0__6), .QB (\$dummy [6]), .D (
        L0_0_L1_0_Fij_nx272), .CLK (CLK)) ;
    dff L0_0_L1_0_Fij_reg_Dout_7 (.Q (FilterDout_0__0__7), .QB (\$dummy [7]), .D (
        L0_0_L1_0_Fij_nx282), .CLK (CLK)) ;
    buf02 L0_0_L1_0_Fij_ix330 (.Y (L0_0_L1_0_Fij_nx331), .A (EN)) ;
    buf02 L0_0_L1_0_Fij_ix332 (.Y (L0_0_L1_0_Fij_nx333), .A (EN)) ;
    dff L0_0_L1_0_Wij_reg_Dout_0 (.Q (WindowDout_0__0__0), .QB (\$dummy [8]), .D (
        L0_0_L1_0_Wij_nx212), .CLK (CLK)) ;
    nor02_2x L0_0_L1_0_Wij_ix297 (.Y (L0_0_L1_0_Wij_nx296), .A0 (RST), .A1 (
             L0_0_L1_0_Wij_nx331)) ;
    dff L0_0_L1_0_Wij_reg_Dout_1 (.Q (WindowDout_0__0__1), .QB (\$dummy [9]), .D (
        L0_0_L1_0_Wij_nx222), .CLK (CLK)) ;
    dff L0_0_L1_0_Wij_reg_Dout_2 (.Q (WindowDout_0__0__2), .QB (\$dummy [10]), .D (
        L0_0_L1_0_Wij_nx232), .CLK (CLK)) ;
    dff L0_0_L1_0_Wij_reg_Dout_3 (.Q (WindowDout_0__0__3), .QB (\$dummy [11]), .D (
        L0_0_L1_0_Wij_nx242), .CLK (CLK)) ;
    dff L0_0_L1_0_Wij_reg_Dout_4 (.Q (WindowDout_0__0__4), .QB (\$dummy [12]), .D (
        L0_0_L1_0_Wij_nx252), .CLK (CLK)) ;
    dff L0_0_L1_0_Wij_reg_Dout_5 (.Q (WindowDout_0__0__5), .QB (\$dummy [13]), .D (
        L0_0_L1_0_Wij_nx262), .CLK (CLK)) ;
    dff L0_0_L1_0_Wij_reg_Dout_6 (.Q (WindowDout_0__0__6), .QB (\$dummy [14]), .D (
        L0_0_L1_0_Wij_nx272), .CLK (CLK)) ;
    dff L0_0_L1_0_Wij_reg_Dout_7 (.Q (WindowDout_0__0__7), .QB (\$dummy [15]), .D (
        L0_0_L1_0_Wij_nx282), .CLK (CLK)) ;
    buf02 L0_0_L1_0_Wij_ix330 (.Y (L0_0_L1_0_Wij_nx331), .A (EN_dup_1004)) ;
    buf02 L0_0_L1_0_Wij_ix332 (.Y (L0_0_L1_0_Wij_nx333), .A (EN_dup_1004)) ;
    dff L0_0_L1_1_Fij_reg_Dout_0 (.Q (FilterDout_0__1__0), .QB (\$dummy [16]), .D (
        L0_0_L1_1_Fij_nx212), .CLK (CLK)) ;
    nor02_2x L0_0_L1_1_Fij_ix297 (.Y (L0_0_L1_1_Fij_nx296), .A0 (RST), .A1 (
             L0_0_L1_1_Fij_nx331)) ;
    dff L0_0_L1_1_Fij_reg_Dout_1 (.Q (FilterDout_0__1__1), .QB (\$dummy [17]), .D (
        L0_0_L1_1_Fij_nx222), .CLK (CLK)) ;
    dff L0_0_L1_1_Fij_reg_Dout_2 (.Q (FilterDout_0__1__2), .QB (\$dummy [18]), .D (
        L0_0_L1_1_Fij_nx232), .CLK (CLK)) ;
    dff L0_0_L1_1_Fij_reg_Dout_3 (.Q (FilterDout_0__1__3), .QB (\$dummy [19]), .D (
        L0_0_L1_1_Fij_nx242), .CLK (CLK)) ;
    dff L0_0_L1_1_Fij_reg_Dout_4 (.Q (FilterDout_0__1__4), .QB (\$dummy [20]), .D (
        L0_0_L1_1_Fij_nx252), .CLK (CLK)) ;
    dff L0_0_L1_1_Fij_reg_Dout_5 (.Q (FilterDout_0__1__5), .QB (\$dummy [21]), .D (
        L0_0_L1_1_Fij_nx262), .CLK (CLK)) ;
    dff L0_0_L1_1_Fij_reg_Dout_6 (.Q (FilterDout_0__1__6), .QB (\$dummy [22]), .D (
        L0_0_L1_1_Fij_nx272), .CLK (CLK)) ;
    dff L0_0_L1_1_Fij_reg_Dout_7 (.Q (FilterDout_0__1__7), .QB (\$dummy [23]), .D (
        L0_0_L1_1_Fij_nx282), .CLK (CLK)) ;
    buf02 L0_0_L1_1_Fij_ix330 (.Y (L0_0_L1_1_Fij_nx331), .A (EN_dup_1015)) ;
    buf02 L0_0_L1_1_Fij_ix332 (.Y (L0_0_L1_1_Fij_nx333), .A (EN_dup_1015)) ;
    dff L0_0_L1_1_Wij_reg_Dout_0 (.Q (WindowDout_0__1__0), .QB (\$dummy [24]), .D (
        L0_0_L1_1_Wij_nx212), .CLK (CLK)) ;
    nor02_2x L0_0_L1_1_Wij_ix297 (.Y (L0_0_L1_1_Wij_nx296), .A0 (RST), .A1 (
             L0_0_L1_1_Wij_nx331)) ;
    dff L0_0_L1_1_Wij_reg_Dout_1 (.Q (WindowDout_0__1__1), .QB (\$dummy [25]), .D (
        L0_0_L1_1_Wij_nx222), .CLK (CLK)) ;
    dff L0_0_L1_1_Wij_reg_Dout_2 (.Q (WindowDout_0__1__2), .QB (\$dummy [26]), .D (
        L0_0_L1_1_Wij_nx232), .CLK (CLK)) ;
    dff L0_0_L1_1_Wij_reg_Dout_3 (.Q (WindowDout_0__1__3), .QB (\$dummy [27]), .D (
        L0_0_L1_1_Wij_nx242), .CLK (CLK)) ;
    dff L0_0_L1_1_Wij_reg_Dout_4 (.Q (WindowDout_0__1__4), .QB (\$dummy [28]), .D (
        L0_0_L1_1_Wij_nx252), .CLK (CLK)) ;
    dff L0_0_L1_1_Wij_reg_Dout_5 (.Q (WindowDout_0__1__5), .QB (\$dummy [29]), .D (
        L0_0_L1_1_Wij_nx262), .CLK (CLK)) ;
    dff L0_0_L1_1_Wij_reg_Dout_6 (.Q (WindowDout_0__1__6), .QB (\$dummy [30]), .D (
        L0_0_L1_1_Wij_nx272), .CLK (CLK)) ;
    dff L0_0_L1_1_Wij_reg_Dout_7 (.Q (WindowDout_0__1__7), .QB (\$dummy [31]), .D (
        L0_0_L1_1_Wij_nx282), .CLK (CLK)) ;
    buf02 L0_0_L1_1_Wij_ix330 (.Y (L0_0_L1_1_Wij_nx331), .A (EN_dup_1026)) ;
    buf02 L0_0_L1_1_Wij_ix332 (.Y (L0_0_L1_1_Wij_nx333), .A (EN_dup_1026)) ;
    dff L0_0_L1_2_Fij_reg_Dout_0 (.Q (FilterDout_0__2__0), .QB (\$dummy [32]), .D (
        L0_0_L1_2_Fij_nx212), .CLK (CLK)) ;
    nor02_2x L0_0_L1_2_Fij_ix297 (.Y (L0_0_L1_2_Fij_nx296), .A0 (RST), .A1 (
             L0_0_L1_2_Fij_nx331)) ;
    dff L0_0_L1_2_Fij_reg_Dout_1 (.Q (FilterDout_0__2__1), .QB (\$dummy [33]), .D (
        L0_0_L1_2_Fij_nx222), .CLK (CLK)) ;
    dff L0_0_L1_2_Fij_reg_Dout_2 (.Q (FilterDout_0__2__2), .QB (\$dummy [34]), .D (
        L0_0_L1_2_Fij_nx232), .CLK (CLK)) ;
    dff L0_0_L1_2_Fij_reg_Dout_3 (.Q (FilterDout_0__2__3), .QB (\$dummy [35]), .D (
        L0_0_L1_2_Fij_nx242), .CLK (CLK)) ;
    dff L0_0_L1_2_Fij_reg_Dout_4 (.Q (FilterDout_0__2__4), .QB (\$dummy [36]), .D (
        L0_0_L1_2_Fij_nx252), .CLK (CLK)) ;
    dff L0_0_L1_2_Fij_reg_Dout_5 (.Q (FilterDout_0__2__5), .QB (\$dummy [37]), .D (
        L0_0_L1_2_Fij_nx262), .CLK (CLK)) ;
    dff L0_0_L1_2_Fij_reg_Dout_6 (.Q (FilterDout_0__2__6), .QB (\$dummy [38]), .D (
        L0_0_L1_2_Fij_nx272), .CLK (CLK)) ;
    dff L0_0_L1_2_Fij_reg_Dout_7 (.Q (FilterDout_0__2__7), .QB (\$dummy [39]), .D (
        L0_0_L1_2_Fij_nx282), .CLK (CLK)) ;
    buf02 L0_0_L1_2_Fij_ix330 (.Y (L0_0_L1_2_Fij_nx331), .A (EN_dup_1015)) ;
    buf02 L0_0_L1_2_Fij_ix332 (.Y (L0_0_L1_2_Fij_nx333), .A (EN_dup_1015)) ;
    dff L0_0_L1_2_Wij_reg_Dout_0 (.Q (WindowDout_0__2__0), .QB (\$dummy [40]), .D (
        L0_0_L1_2_Wij_nx212), .CLK (CLK)) ;
    nor02_2x L0_0_L1_2_Wij_ix297 (.Y (L0_0_L1_2_Wij_nx296), .A0 (RST), .A1 (
             L0_0_L1_2_Wij_nx331)) ;
    dff L0_0_L1_2_Wij_reg_Dout_1 (.Q (WindowDout_0__2__1), .QB (\$dummy [41]), .D (
        L0_0_L1_2_Wij_nx222), .CLK (CLK)) ;
    dff L0_0_L1_2_Wij_reg_Dout_2 (.Q (WindowDout_0__2__2), .QB (\$dummy [42]), .D (
        L0_0_L1_2_Wij_nx232), .CLK (CLK)) ;
    dff L0_0_L1_2_Wij_reg_Dout_3 (.Q (WindowDout_0__2__3), .QB (\$dummy [43]), .D (
        L0_0_L1_2_Wij_nx242), .CLK (CLK)) ;
    dff L0_0_L1_2_Wij_reg_Dout_4 (.Q (WindowDout_0__2__4), .QB (\$dummy [44]), .D (
        L0_0_L1_2_Wij_nx252), .CLK (CLK)) ;
    dff L0_0_L1_2_Wij_reg_Dout_5 (.Q (WindowDout_0__2__5), .QB (\$dummy [45]), .D (
        L0_0_L1_2_Wij_nx262), .CLK (CLK)) ;
    dff L0_0_L1_2_Wij_reg_Dout_6 (.Q (WindowDout_0__2__6), .QB (\$dummy [46]), .D (
        L0_0_L1_2_Wij_nx272), .CLK (CLK)) ;
    dff L0_0_L1_2_Wij_reg_Dout_7 (.Q (WindowDout_0__2__7), .QB (\$dummy [47]), .D (
        L0_0_L1_2_Wij_nx282), .CLK (CLK)) ;
    buf02 L0_0_L1_2_Wij_ix330 (.Y (L0_0_L1_2_Wij_nx331), .A (EN_dup_1026)) ;
    buf02 L0_0_L1_2_Wij_ix332 (.Y (L0_0_L1_2_Wij_nx333), .A (EN_dup_1026)) ;
    dff L0_0_L1_3_Fij_reg_Dout_0 (.Q (FilterDout_0__3__0), .QB (\$dummy [48]), .D (
        L0_0_L1_3_Fij_nx212), .CLK (CLK)) ;
    nor02_2x L0_0_L1_3_Fij_ix297 (.Y (L0_0_L1_3_Fij_nx296), .A0 (RST), .A1 (
             L0_0_L1_3_Fij_nx331)) ;
    dff L0_0_L1_3_Fij_reg_Dout_1 (.Q (FilterDout_0__3__1), .QB (\$dummy [49]), .D (
        L0_0_L1_3_Fij_nx222), .CLK (CLK)) ;
    dff L0_0_L1_3_Fij_reg_Dout_2 (.Q (FilterDout_0__3__2), .QB (\$dummy [50]), .D (
        L0_0_L1_3_Fij_nx232), .CLK (CLK)) ;
    dff L0_0_L1_3_Fij_reg_Dout_3 (.Q (FilterDout_0__3__3), .QB (\$dummy [51]), .D (
        L0_0_L1_3_Fij_nx242), .CLK (CLK)) ;
    dff L0_0_L1_3_Fij_reg_Dout_4 (.Q (FilterDout_0__3__4), .QB (\$dummy [52]), .D (
        L0_0_L1_3_Fij_nx252), .CLK (CLK)) ;
    dff L0_0_L1_3_Fij_reg_Dout_5 (.Q (FilterDout_0__3__5), .QB (\$dummy [53]), .D (
        L0_0_L1_3_Fij_nx262), .CLK (CLK)) ;
    dff L0_0_L1_3_Fij_reg_Dout_6 (.Q (FilterDout_0__3__6), .QB (\$dummy [54]), .D (
        L0_0_L1_3_Fij_nx272), .CLK (CLK)) ;
    dff L0_0_L1_3_Fij_reg_Dout_7 (.Q (FilterDout_0__3__7), .QB (\$dummy [55]), .D (
        L0_0_L1_3_Fij_nx282), .CLK (CLK)) ;
    buf02 L0_0_L1_3_Fij_ix330 (.Y (L0_0_L1_3_Fij_nx331), .A (EN_dup_1015)) ;
    buf02 L0_0_L1_3_Fij_ix332 (.Y (L0_0_L1_3_Fij_nx333), .A (EN_dup_1015)) ;
    dff L0_0_L1_3_Wij_reg_Dout_0 (.Q (WindowDout_0__3__0), .QB (\$dummy [56]), .D (
        L0_0_L1_3_Wij_nx212), .CLK (CLK)) ;
    nor02_2x L0_0_L1_3_Wij_ix297 (.Y (L0_0_L1_3_Wij_nx296), .A0 (RST), .A1 (
             L0_0_L1_3_Wij_nx331)) ;
    dff L0_0_L1_3_Wij_reg_Dout_1 (.Q (WindowDout_0__3__1), .QB (\$dummy [57]), .D (
        L0_0_L1_3_Wij_nx222), .CLK (CLK)) ;
    dff L0_0_L1_3_Wij_reg_Dout_2 (.Q (WindowDout_0__3__2), .QB (\$dummy [58]), .D (
        L0_0_L1_3_Wij_nx232), .CLK (CLK)) ;
    dff L0_0_L1_3_Wij_reg_Dout_3 (.Q (WindowDout_0__3__3), .QB (\$dummy [59]), .D (
        L0_0_L1_3_Wij_nx242), .CLK (CLK)) ;
    dff L0_0_L1_3_Wij_reg_Dout_4 (.Q (WindowDout_0__3__4), .QB (\$dummy [60]), .D (
        L0_0_L1_3_Wij_nx252), .CLK (CLK)) ;
    dff L0_0_L1_3_Wij_reg_Dout_5 (.Q (WindowDout_0__3__5), .QB (\$dummy [61]), .D (
        L0_0_L1_3_Wij_nx262), .CLK (CLK)) ;
    dff L0_0_L1_3_Wij_reg_Dout_6 (.Q (WindowDout_0__3__6), .QB (\$dummy [62]), .D (
        L0_0_L1_3_Wij_nx272), .CLK (CLK)) ;
    dff L0_0_L1_3_Wij_reg_Dout_7 (.Q (WindowDout_0__3__7), .QB (\$dummy [63]), .D (
        L0_0_L1_3_Wij_nx282), .CLK (CLK)) ;
    buf02 L0_0_L1_3_Wij_ix330 (.Y (L0_0_L1_3_Wij_nx331), .A (EN_dup_1026)) ;
    buf02 L0_0_L1_3_Wij_ix332 (.Y (L0_0_L1_3_Wij_nx333), .A (EN_dup_1026)) ;
    dff L0_0_L1_4_Fij_reg_Dout_0 (.Q (FilterDout_0__4__0), .QB (\$dummy [64]), .D (
        L0_0_L1_4_Fij_nx212), .CLK (CLK)) ;
    nor02_2x L0_0_L1_4_Fij_ix297 (.Y (L0_0_L1_4_Fij_nx296), .A0 (RST), .A1 (
             L0_0_L1_4_Fij_nx331)) ;
    dff L0_0_L1_4_Fij_reg_Dout_1 (.Q (FilterDout_0__4__1), .QB (\$dummy [65]), .D (
        L0_0_L1_4_Fij_nx222), .CLK (CLK)) ;
    dff L0_0_L1_4_Fij_reg_Dout_2 (.Q (FilterDout_0__4__2), .QB (\$dummy [66]), .D (
        L0_0_L1_4_Fij_nx232), .CLK (CLK)) ;
    dff L0_0_L1_4_Fij_reg_Dout_3 (.Q (FilterDout_0__4__3), .QB (\$dummy [67]), .D (
        L0_0_L1_4_Fij_nx242), .CLK (CLK)) ;
    dff L0_0_L1_4_Fij_reg_Dout_4 (.Q (FilterDout_0__4__4), .QB (\$dummy [68]), .D (
        L0_0_L1_4_Fij_nx252), .CLK (CLK)) ;
    dff L0_0_L1_4_Fij_reg_Dout_5 (.Q (FilterDout_0__4__5), .QB (\$dummy [69]), .D (
        L0_0_L1_4_Fij_nx262), .CLK (CLK)) ;
    dff L0_0_L1_4_Fij_reg_Dout_6 (.Q (FilterDout_0__4__6), .QB (\$dummy [70]), .D (
        L0_0_L1_4_Fij_nx272), .CLK (CLK)) ;
    dff L0_0_L1_4_Fij_reg_Dout_7 (.Q (FilterDout_0__4__7), .QB (\$dummy [71]), .D (
        L0_0_L1_4_Fij_nx282), .CLK (CLK)) ;
    buf02 L0_0_L1_4_Fij_ix330 (.Y (L0_0_L1_4_Fij_nx331), .A (EN_dup_1081)) ;
    buf02 L0_0_L1_4_Fij_ix332 (.Y (L0_0_L1_4_Fij_nx333), .A (EN_dup_1081)) ;
    dff L0_0_L1_4_Wij_reg_Dout_0 (.Q (WindowDout_0__4__0), .QB (\$dummy [72]), .D (
        L0_0_L1_4_Wij_nx212), .CLK (CLK)) ;
    nor02_2x L0_0_L1_4_Wij_ix297 (.Y (L0_0_L1_4_Wij_nx296), .A0 (RST), .A1 (
             L0_0_L1_4_Wij_nx331)) ;
    dff L0_0_L1_4_Wij_reg_Dout_1 (.Q (WindowDout_0__4__1), .QB (\$dummy [73]), .D (
        L0_0_L1_4_Wij_nx222), .CLK (CLK)) ;
    dff L0_0_L1_4_Wij_reg_Dout_2 (.Q (WindowDout_0__4__2), .QB (\$dummy [74]), .D (
        L0_0_L1_4_Wij_nx232), .CLK (CLK)) ;
    dff L0_0_L1_4_Wij_reg_Dout_3 (.Q (WindowDout_0__4__3), .QB (\$dummy [75]), .D (
        L0_0_L1_4_Wij_nx242), .CLK (CLK)) ;
    dff L0_0_L1_4_Wij_reg_Dout_4 (.Q (WindowDout_0__4__4), .QB (\$dummy [76]), .D (
        L0_0_L1_4_Wij_nx252), .CLK (CLK)) ;
    dff L0_0_L1_4_Wij_reg_Dout_5 (.Q (WindowDout_0__4__5), .QB (\$dummy [77]), .D (
        L0_0_L1_4_Wij_nx262), .CLK (CLK)) ;
    dff L0_0_L1_4_Wij_reg_Dout_6 (.Q (WindowDout_0__4__6), .QB (\$dummy [78]), .D (
        L0_0_L1_4_Wij_nx272), .CLK (CLK)) ;
    dff L0_0_L1_4_Wij_reg_Dout_7 (.Q (WindowDout_0__4__7), .QB (\$dummy [79]), .D (
        L0_0_L1_4_Wij_nx282), .CLK (CLK)) ;
    buf02 L0_0_L1_4_Wij_ix330 (.Y (L0_0_L1_4_Wij_nx331), .A (EN_dup_1092)) ;
    buf02 L0_0_L1_4_Wij_ix332 (.Y (L0_0_L1_4_Wij_nx333), .A (EN_dup_1092)) ;
    dff L0_1_L1_0_Fij_reg_Dout_0 (.Q (FilterDout_1__0__0), .QB (\$dummy [80]), .D (
        L0_1_L1_0_Fij_nx212), .CLK (CLK)) ;
    nor02_2x L0_1_L1_0_Fij_ix297 (.Y (L0_1_L1_0_Fij_nx296), .A0 (RST), .A1 (
             L0_1_L1_0_Fij_nx331)) ;
    dff L0_1_L1_0_Fij_reg_Dout_1 (.Q (FilterDout_1__0__1), .QB (\$dummy [81]), .D (
        L0_1_L1_0_Fij_nx222), .CLK (CLK)) ;
    dff L0_1_L1_0_Fij_reg_Dout_2 (.Q (FilterDout_1__0__2), .QB (\$dummy [82]), .D (
        L0_1_L1_0_Fij_nx232), .CLK (CLK)) ;
    dff L0_1_L1_0_Fij_reg_Dout_3 (.Q (FilterDout_1__0__3), .QB (\$dummy [83]), .D (
        L0_1_L1_0_Fij_nx242), .CLK (CLK)) ;
    dff L0_1_L1_0_Fij_reg_Dout_4 (.Q (FilterDout_1__0__4), .QB (\$dummy [84]), .D (
        L0_1_L1_0_Fij_nx252), .CLK (CLK)) ;
    dff L0_1_L1_0_Fij_reg_Dout_5 (.Q (FilterDout_1__0__5), .QB (\$dummy [85]), .D (
        L0_1_L1_0_Fij_nx262), .CLK (CLK)) ;
    dff L0_1_L1_0_Fij_reg_Dout_6 (.Q (FilterDout_1__0__6), .QB (\$dummy [86]), .D (
        L0_1_L1_0_Fij_nx272), .CLK (CLK)) ;
    dff L0_1_L1_0_Fij_reg_Dout_7 (.Q (FilterDout_1__0__7), .QB (\$dummy [87]), .D (
        L0_1_L1_0_Fij_nx282), .CLK (CLK)) ;
    buf02 L0_1_L1_0_Fij_ix330 (.Y (L0_1_L1_0_Fij_nx331), .A (EN_dup_1081)) ;
    buf02 L0_1_L1_0_Fij_ix332 (.Y (L0_1_L1_0_Fij_nx333), .A (EN_dup_1081)) ;
    dff L0_1_L1_0_Wij_reg_Dout_0 (.Q (WindowDout_1__0__0), .QB (\$dummy [88]), .D (
        L0_1_L1_0_Wij_nx212), .CLK (CLK)) ;
    nor02_2x L0_1_L1_0_Wij_ix297 (.Y (L0_1_L1_0_Wij_nx296), .A0 (RST), .A1 (
             L0_1_L1_0_Wij_nx331)) ;
    dff L0_1_L1_0_Wij_reg_Dout_1 (.Q (WindowDout_1__0__1), .QB (\$dummy [89]), .D (
        L0_1_L1_0_Wij_nx222), .CLK (CLK)) ;
    dff L0_1_L1_0_Wij_reg_Dout_2 (.Q (WindowDout_1__0__2), .QB (\$dummy [90]), .D (
        L0_1_L1_0_Wij_nx232), .CLK (CLK)) ;
    dff L0_1_L1_0_Wij_reg_Dout_3 (.Q (WindowDout_1__0__3), .QB (\$dummy [91]), .D (
        L0_1_L1_0_Wij_nx242), .CLK (CLK)) ;
    dff L0_1_L1_0_Wij_reg_Dout_4 (.Q (WindowDout_1__0__4), .QB (\$dummy [92]), .D (
        L0_1_L1_0_Wij_nx252), .CLK (CLK)) ;
    dff L0_1_L1_0_Wij_reg_Dout_5 (.Q (WindowDout_1__0__5), .QB (\$dummy [93]), .D (
        L0_1_L1_0_Wij_nx262), .CLK (CLK)) ;
    dff L0_1_L1_0_Wij_reg_Dout_6 (.Q (WindowDout_1__0__6), .QB (\$dummy [94]), .D (
        L0_1_L1_0_Wij_nx272), .CLK (CLK)) ;
    dff L0_1_L1_0_Wij_reg_Dout_7 (.Q (WindowDout_1__0__7), .QB (\$dummy [95]), .D (
        L0_1_L1_0_Wij_nx282), .CLK (CLK)) ;
    buf02 L0_1_L1_0_Wij_ix330 (.Y (L0_1_L1_0_Wij_nx331), .A (EN_dup_1092)) ;
    buf02 L0_1_L1_0_Wij_ix332 (.Y (L0_1_L1_0_Wij_nx333), .A (EN_dup_1092)) ;
    dff L0_1_L1_1_Fij_reg_Dout_0 (.Q (FilterDout_1__1__0), .QB (\$dummy [96]), .D (
        L0_1_L1_1_Fij_nx212), .CLK (CLK)) ;
    nor02_2x L0_1_L1_1_Fij_ix297 (.Y (L0_1_L1_1_Fij_nx296), .A0 (RST), .A1 (
             L0_1_L1_1_Fij_nx331)) ;
    dff L0_1_L1_1_Fij_reg_Dout_1 (.Q (FilterDout_1__1__1), .QB (\$dummy [97]), .D (
        L0_1_L1_1_Fij_nx222), .CLK (CLK)) ;
    dff L0_1_L1_1_Fij_reg_Dout_2 (.Q (FilterDout_1__1__2), .QB (\$dummy [98]), .D (
        L0_1_L1_1_Fij_nx232), .CLK (CLK)) ;
    dff L0_1_L1_1_Fij_reg_Dout_3 (.Q (FilterDout_1__1__3), .QB (\$dummy [99]), .D (
        L0_1_L1_1_Fij_nx242), .CLK (CLK)) ;
    dff L0_1_L1_1_Fij_reg_Dout_4 (.Q (FilterDout_1__1__4), .QB (\$dummy [100]), 
        .D (L0_1_L1_1_Fij_nx252), .CLK (CLK)) ;
    dff L0_1_L1_1_Fij_reg_Dout_5 (.Q (FilterDout_1__1__5), .QB (\$dummy [101]), 
        .D (L0_1_L1_1_Fij_nx262), .CLK (CLK)) ;
    dff L0_1_L1_1_Fij_reg_Dout_6 (.Q (FilterDout_1__1__6), .QB (\$dummy [102]), 
        .D (L0_1_L1_1_Fij_nx272), .CLK (CLK)) ;
    dff L0_1_L1_1_Fij_reg_Dout_7 (.Q (FilterDout_1__1__7), .QB (\$dummy [103]), 
        .D (L0_1_L1_1_Fij_nx282), .CLK (CLK)) ;
    buf02 L0_1_L1_1_Fij_ix330 (.Y (L0_1_L1_1_Fij_nx331), .A (EN_dup_1081)) ;
    buf02 L0_1_L1_1_Fij_ix332 (.Y (L0_1_L1_1_Fij_nx333), .A (EN_dup_1081)) ;
    dff L0_1_L1_1_Wij_reg_Dout_0 (.Q (WindowDout_1__1__0), .QB (\$dummy [104]), 
        .D (L0_1_L1_1_Wij_nx212), .CLK (CLK)) ;
    nor02_2x L0_1_L1_1_Wij_ix297 (.Y (L0_1_L1_1_Wij_nx296), .A0 (RST), .A1 (
             L0_1_L1_1_Wij_nx331)) ;
    dff L0_1_L1_1_Wij_reg_Dout_1 (.Q (WindowDout_1__1__1), .QB (\$dummy [105]), 
        .D (L0_1_L1_1_Wij_nx222), .CLK (CLK)) ;
    dff L0_1_L1_1_Wij_reg_Dout_2 (.Q (WindowDout_1__1__2), .QB (\$dummy [106]), 
        .D (L0_1_L1_1_Wij_nx232), .CLK (CLK)) ;
    dff L0_1_L1_1_Wij_reg_Dout_3 (.Q (WindowDout_1__1__3), .QB (\$dummy [107]), 
        .D (L0_1_L1_1_Wij_nx242), .CLK (CLK)) ;
    dff L0_1_L1_1_Wij_reg_Dout_4 (.Q (WindowDout_1__1__4), .QB (\$dummy [108]), 
        .D (L0_1_L1_1_Wij_nx252), .CLK (CLK)) ;
    dff L0_1_L1_1_Wij_reg_Dout_5 (.Q (WindowDout_1__1__5), .QB (\$dummy [109]), 
        .D (L0_1_L1_1_Wij_nx262), .CLK (CLK)) ;
    dff L0_1_L1_1_Wij_reg_Dout_6 (.Q (WindowDout_1__1__6), .QB (\$dummy [110]), 
        .D (L0_1_L1_1_Wij_nx272), .CLK (CLK)) ;
    dff L0_1_L1_1_Wij_reg_Dout_7 (.Q (WindowDout_1__1__7), .QB (\$dummy [111]), 
        .D (L0_1_L1_1_Wij_nx282), .CLK (CLK)) ;
    buf02 L0_1_L1_1_Wij_ix330 (.Y (L0_1_L1_1_Wij_nx331), .A (EN_dup_1092)) ;
    buf02 L0_1_L1_1_Wij_ix332 (.Y (L0_1_L1_1_Wij_nx333), .A (EN_dup_1092)) ;
    dff L0_1_L1_2_Fij_reg_Dout_0 (.Q (FilterDout_1__2__0), .QB (\$dummy [112]), 
        .D (L0_1_L1_2_Fij_nx212), .CLK (CLK)) ;
    nor02_2x L0_1_L1_2_Fij_ix297 (.Y (L0_1_L1_2_Fij_nx296), .A0 (RST), .A1 (
             L0_1_L1_2_Fij_nx331)) ;
    dff L0_1_L1_2_Fij_reg_Dout_1 (.Q (FilterDout_1__2__1), .QB (\$dummy [113]), 
        .D (L0_1_L1_2_Fij_nx222), .CLK (CLK)) ;
    dff L0_1_L1_2_Fij_reg_Dout_2 (.Q (FilterDout_1__2__2), .QB (\$dummy [114]), 
        .D (L0_1_L1_2_Fij_nx232), .CLK (CLK)) ;
    dff L0_1_L1_2_Fij_reg_Dout_3 (.Q (FilterDout_1__2__3), .QB (\$dummy [115]), 
        .D (L0_1_L1_2_Fij_nx242), .CLK (CLK)) ;
    dff L0_1_L1_2_Fij_reg_Dout_4 (.Q (FilterDout_1__2__4), .QB (\$dummy [116]), 
        .D (L0_1_L1_2_Fij_nx252), .CLK (CLK)) ;
    dff L0_1_L1_2_Fij_reg_Dout_5 (.Q (FilterDout_1__2__5), .QB (\$dummy [117]), 
        .D (L0_1_L1_2_Fij_nx262), .CLK (CLK)) ;
    dff L0_1_L1_2_Fij_reg_Dout_6 (.Q (FilterDout_1__2__6), .QB (\$dummy [118]), 
        .D (L0_1_L1_2_Fij_nx272), .CLK (CLK)) ;
    dff L0_1_L1_2_Fij_reg_Dout_7 (.Q (FilterDout_1__2__7), .QB (\$dummy [119]), 
        .D (L0_1_L1_2_Fij_nx282), .CLK (CLK)) ;
    buf02 L0_1_L1_2_Fij_ix330 (.Y (L0_1_L1_2_Fij_nx331), .A (EN_dup_1147)) ;
    buf02 L0_1_L1_2_Fij_ix332 (.Y (L0_1_L1_2_Fij_nx333), .A (EN_dup_1147)) ;
    dff L0_1_L1_2_Wij_reg_Dout_0 (.Q (WindowDout_1__2__0), .QB (\$dummy [120]), 
        .D (L0_1_L1_2_Wij_nx212), .CLK (CLK)) ;
    nor02_2x L0_1_L1_2_Wij_ix297 (.Y (L0_1_L1_2_Wij_nx296), .A0 (RST), .A1 (
             L0_1_L1_2_Wij_nx331)) ;
    dff L0_1_L1_2_Wij_reg_Dout_1 (.Q (WindowDout_1__2__1), .QB (\$dummy [121]), 
        .D (L0_1_L1_2_Wij_nx222), .CLK (CLK)) ;
    dff L0_1_L1_2_Wij_reg_Dout_2 (.Q (WindowDout_1__2__2), .QB (\$dummy [122]), 
        .D (L0_1_L1_2_Wij_nx232), .CLK (CLK)) ;
    dff L0_1_L1_2_Wij_reg_Dout_3 (.Q (WindowDout_1__2__3), .QB (\$dummy [123]), 
        .D (L0_1_L1_2_Wij_nx242), .CLK (CLK)) ;
    dff L0_1_L1_2_Wij_reg_Dout_4 (.Q (WindowDout_1__2__4), .QB (\$dummy [124]), 
        .D (L0_1_L1_2_Wij_nx252), .CLK (CLK)) ;
    dff L0_1_L1_2_Wij_reg_Dout_5 (.Q (WindowDout_1__2__5), .QB (\$dummy [125]), 
        .D (L0_1_L1_2_Wij_nx262), .CLK (CLK)) ;
    dff L0_1_L1_2_Wij_reg_Dout_6 (.Q (WindowDout_1__2__6), .QB (\$dummy [126]), 
        .D (L0_1_L1_2_Wij_nx272), .CLK (CLK)) ;
    dff L0_1_L1_2_Wij_reg_Dout_7 (.Q (WindowDout_1__2__7), .QB (\$dummy [127]), 
        .D (L0_1_L1_2_Wij_nx282), .CLK (CLK)) ;
    buf02 L0_1_L1_2_Wij_ix330 (.Y (L0_1_L1_2_Wij_nx331), .A (EN_dup_1158)) ;
    buf02 L0_1_L1_2_Wij_ix332 (.Y (L0_1_L1_2_Wij_nx333), .A (EN_dup_1158)) ;
    dff L0_1_L1_3_Fij_reg_Dout_0 (.Q (FilterDout_1__3__0), .QB (\$dummy [128]), 
        .D (L0_1_L1_3_Fij_nx212), .CLK (CLK)) ;
    nor02_2x L0_1_L1_3_Fij_ix297 (.Y (L0_1_L1_3_Fij_nx296), .A0 (RST), .A1 (
             L0_1_L1_3_Fij_nx331)) ;
    dff L0_1_L1_3_Fij_reg_Dout_1 (.Q (FilterDout_1__3__1), .QB (\$dummy [129]), 
        .D (L0_1_L1_3_Fij_nx222), .CLK (CLK)) ;
    dff L0_1_L1_3_Fij_reg_Dout_2 (.Q (FilterDout_1__3__2), .QB (\$dummy [130]), 
        .D (L0_1_L1_3_Fij_nx232), .CLK (CLK)) ;
    dff L0_1_L1_3_Fij_reg_Dout_3 (.Q (FilterDout_1__3__3), .QB (\$dummy [131]), 
        .D (L0_1_L1_3_Fij_nx242), .CLK (CLK)) ;
    dff L0_1_L1_3_Fij_reg_Dout_4 (.Q (FilterDout_1__3__4), .QB (\$dummy [132]), 
        .D (L0_1_L1_3_Fij_nx252), .CLK (CLK)) ;
    dff L0_1_L1_3_Fij_reg_Dout_5 (.Q (FilterDout_1__3__5), .QB (\$dummy [133]), 
        .D (L0_1_L1_3_Fij_nx262), .CLK (CLK)) ;
    dff L0_1_L1_3_Fij_reg_Dout_6 (.Q (FilterDout_1__3__6), .QB (\$dummy [134]), 
        .D (L0_1_L1_3_Fij_nx272), .CLK (CLK)) ;
    dff L0_1_L1_3_Fij_reg_Dout_7 (.Q (FilterDout_1__3__7), .QB (\$dummy [135]), 
        .D (L0_1_L1_3_Fij_nx282), .CLK (CLK)) ;
    buf02 L0_1_L1_3_Fij_ix330 (.Y (L0_1_L1_3_Fij_nx331), .A (EN_dup_1147)) ;
    buf02 L0_1_L1_3_Fij_ix332 (.Y (L0_1_L1_3_Fij_nx333), .A (EN_dup_1147)) ;
    dff L0_1_L1_3_Wij_reg_Dout_0 (.Q (WindowDout_1__3__0), .QB (\$dummy [136]), 
        .D (L0_1_L1_3_Wij_nx212), .CLK (CLK)) ;
    nor02_2x L0_1_L1_3_Wij_ix297 (.Y (L0_1_L1_3_Wij_nx296), .A0 (RST), .A1 (
             L0_1_L1_3_Wij_nx331)) ;
    dff L0_1_L1_3_Wij_reg_Dout_1 (.Q (WindowDout_1__3__1), .QB (\$dummy [137]), 
        .D (L0_1_L1_3_Wij_nx222), .CLK (CLK)) ;
    dff L0_1_L1_3_Wij_reg_Dout_2 (.Q (WindowDout_1__3__2), .QB (\$dummy [138]), 
        .D (L0_1_L1_3_Wij_nx232), .CLK (CLK)) ;
    dff L0_1_L1_3_Wij_reg_Dout_3 (.Q (WindowDout_1__3__3), .QB (\$dummy [139]), 
        .D (L0_1_L1_3_Wij_nx242), .CLK (CLK)) ;
    dff L0_1_L1_3_Wij_reg_Dout_4 (.Q (WindowDout_1__3__4), .QB (\$dummy [140]), 
        .D (L0_1_L1_3_Wij_nx252), .CLK (CLK)) ;
    dff L0_1_L1_3_Wij_reg_Dout_5 (.Q (WindowDout_1__3__5), .QB (\$dummy [141]), 
        .D (L0_1_L1_3_Wij_nx262), .CLK (CLK)) ;
    dff L0_1_L1_3_Wij_reg_Dout_6 (.Q (WindowDout_1__3__6), .QB (\$dummy [142]), 
        .D (L0_1_L1_3_Wij_nx272), .CLK (CLK)) ;
    dff L0_1_L1_3_Wij_reg_Dout_7 (.Q (WindowDout_1__3__7), .QB (\$dummy [143]), 
        .D (L0_1_L1_3_Wij_nx282), .CLK (CLK)) ;
    buf02 L0_1_L1_3_Wij_ix330 (.Y (L0_1_L1_3_Wij_nx331), .A (EN_dup_1158)) ;
    buf02 L0_1_L1_3_Wij_ix332 (.Y (L0_1_L1_3_Wij_nx333), .A (EN_dup_1158)) ;
    dff L0_1_L1_4_Fij_reg_Dout_0 (.Q (FilterDout_1__4__0), .QB (\$dummy [144]), 
        .D (L0_1_L1_4_Fij_nx212), .CLK (CLK)) ;
    nor02_2x L0_1_L1_4_Fij_ix297 (.Y (L0_1_L1_4_Fij_nx296), .A0 (RST), .A1 (
             L0_1_L1_4_Fij_nx331)) ;
    dff L0_1_L1_4_Fij_reg_Dout_1 (.Q (FilterDout_1__4__1), .QB (\$dummy [145]), 
        .D (L0_1_L1_4_Fij_nx222), .CLK (CLK)) ;
    dff L0_1_L1_4_Fij_reg_Dout_2 (.Q (FilterDout_1__4__2), .QB (\$dummy [146]), 
        .D (L0_1_L1_4_Fij_nx232), .CLK (CLK)) ;
    dff L0_1_L1_4_Fij_reg_Dout_3 (.Q (FilterDout_1__4__3), .QB (\$dummy [147]), 
        .D (L0_1_L1_4_Fij_nx242), .CLK (CLK)) ;
    dff L0_1_L1_4_Fij_reg_Dout_4 (.Q (FilterDout_1__4__4), .QB (\$dummy [148]), 
        .D (L0_1_L1_4_Fij_nx252), .CLK (CLK)) ;
    dff L0_1_L1_4_Fij_reg_Dout_5 (.Q (FilterDout_1__4__5), .QB (\$dummy [149]), 
        .D (L0_1_L1_4_Fij_nx262), .CLK (CLK)) ;
    dff L0_1_L1_4_Fij_reg_Dout_6 (.Q (FilterDout_1__4__6), .QB (\$dummy [150]), 
        .D (L0_1_L1_4_Fij_nx272), .CLK (CLK)) ;
    dff L0_1_L1_4_Fij_reg_Dout_7 (.Q (FilterDout_1__4__7), .QB (\$dummy [151]), 
        .D (L0_1_L1_4_Fij_nx282), .CLK (CLK)) ;
    buf02 L0_1_L1_4_Fij_ix330 (.Y (L0_1_L1_4_Fij_nx331), .A (EN_dup_1147)) ;
    buf02 L0_1_L1_4_Fij_ix332 (.Y (L0_1_L1_4_Fij_nx333), .A (EN_dup_1147)) ;
    dff L0_1_L1_4_Wij_reg_Dout_0 (.Q (WindowDout_1__4__0), .QB (\$dummy [152]), 
        .D (L0_1_L1_4_Wij_nx212), .CLK (CLK)) ;
    nor02_2x L0_1_L1_4_Wij_ix297 (.Y (L0_1_L1_4_Wij_nx296), .A0 (RST), .A1 (
             L0_1_L1_4_Wij_nx331)) ;
    dff L0_1_L1_4_Wij_reg_Dout_1 (.Q (WindowDout_1__4__1), .QB (\$dummy [153]), 
        .D (L0_1_L1_4_Wij_nx222), .CLK (CLK)) ;
    dff L0_1_L1_4_Wij_reg_Dout_2 (.Q (WindowDout_1__4__2), .QB (\$dummy [154]), 
        .D (L0_1_L1_4_Wij_nx232), .CLK (CLK)) ;
    dff L0_1_L1_4_Wij_reg_Dout_3 (.Q (WindowDout_1__4__3), .QB (\$dummy [155]), 
        .D (L0_1_L1_4_Wij_nx242), .CLK (CLK)) ;
    dff L0_1_L1_4_Wij_reg_Dout_4 (.Q (WindowDout_1__4__4), .QB (\$dummy [156]), 
        .D (L0_1_L1_4_Wij_nx252), .CLK (CLK)) ;
    dff L0_1_L1_4_Wij_reg_Dout_5 (.Q (WindowDout_1__4__5), .QB (\$dummy [157]), 
        .D (L0_1_L1_4_Wij_nx262), .CLK (CLK)) ;
    dff L0_1_L1_4_Wij_reg_Dout_6 (.Q (WindowDout_1__4__6), .QB (\$dummy [158]), 
        .D (L0_1_L1_4_Wij_nx272), .CLK (CLK)) ;
    dff L0_1_L1_4_Wij_reg_Dout_7 (.Q (WindowDout_1__4__7), .QB (\$dummy [159]), 
        .D (L0_1_L1_4_Wij_nx282), .CLK (CLK)) ;
    buf02 L0_1_L1_4_Wij_ix330 (.Y (L0_1_L1_4_Wij_nx331), .A (EN_dup_1158)) ;
    buf02 L0_1_L1_4_Wij_ix332 (.Y (L0_1_L1_4_Wij_nx333), .A (EN_dup_1158)) ;
    dff L0_2_L1_0_Fij_reg_Dout_0 (.Q (FilterDout_2__0__0), .QB (\$dummy [160]), 
        .D (L0_2_L1_0_Fij_nx212), .CLK (CLK)) ;
    nor02_2x L0_2_L1_0_Fij_ix297 (.Y (L0_2_L1_0_Fij_nx296), .A0 (RST), .A1 (
             L0_2_L1_0_Fij_nx331)) ;
    dff L0_2_L1_0_Fij_reg_Dout_1 (.Q (FilterDout_2__0__1), .QB (\$dummy [161]), 
        .D (L0_2_L1_0_Fij_nx222), .CLK (CLK)) ;
    dff L0_2_L1_0_Fij_reg_Dout_2 (.Q (FilterDout_2__0__2), .QB (\$dummy [162]), 
        .D (L0_2_L1_0_Fij_nx232), .CLK (CLK)) ;
    dff L0_2_L1_0_Fij_reg_Dout_3 (.Q (FilterDout_2__0__3), .QB (\$dummy [163]), 
        .D (L0_2_L1_0_Fij_nx242), .CLK (CLK)) ;
    dff L0_2_L1_0_Fij_reg_Dout_4 (.Q (FilterDout_2__0__4), .QB (\$dummy [164]), 
        .D (L0_2_L1_0_Fij_nx252), .CLK (CLK)) ;
    dff L0_2_L1_0_Fij_reg_Dout_5 (.Q (FilterDout_2__0__5), .QB (\$dummy [165]), 
        .D (L0_2_L1_0_Fij_nx262), .CLK (CLK)) ;
    dff L0_2_L1_0_Fij_reg_Dout_6 (.Q (FilterDout_2__0__6), .QB (\$dummy [166]), 
        .D (L0_2_L1_0_Fij_nx272), .CLK (CLK)) ;
    dff L0_2_L1_0_Fij_reg_Dout_7 (.Q (FilterDout_2__0__7), .QB (\$dummy [167]), 
        .D (L0_2_L1_0_Fij_nx282), .CLK (CLK)) ;
    buf02 L0_2_L1_0_Fij_ix330 (.Y (L0_2_L1_0_Fij_nx331), .A (FilterWR)) ;
    buf02 L0_2_L1_0_Fij_ix332 (.Y (L0_2_L1_0_Fij_nx333), .A (FilterWR)) ;
    dff L0_2_L1_0_Wij_reg_Dout_0 (.Q (WindowDout_2__0__0), .QB (\$dummy [168]), 
        .D (L0_2_L1_0_Wij_nx212), .CLK (CLK)) ;
    nor02_2x L0_2_L1_0_Wij_ix297 (.Y (L0_2_L1_0_Wij_nx296), .A0 (RST), .A1 (
             L0_2_L1_0_Wij_nx331)) ;
    dff L0_2_L1_0_Wij_reg_Dout_1 (.Q (WindowDout_2__0__1), .QB (\$dummy [169]), 
        .D (L0_2_L1_0_Wij_nx222), .CLK (CLK)) ;
    dff L0_2_L1_0_Wij_reg_Dout_2 (.Q (WindowDout_2__0__2), .QB (\$dummy [170]), 
        .D (L0_2_L1_0_Wij_nx232), .CLK (CLK)) ;
    dff L0_2_L1_0_Wij_reg_Dout_3 (.Q (WindowDout_2__0__3), .QB (\$dummy [171]), 
        .D (L0_2_L1_0_Wij_nx242), .CLK (CLK)) ;
    dff L0_2_L1_0_Wij_reg_Dout_4 (.Q (WindowDout_2__0__4), .QB (\$dummy [172]), 
        .D (L0_2_L1_0_Wij_nx252), .CLK (CLK)) ;
    dff L0_2_L1_0_Wij_reg_Dout_5 (.Q (WindowDout_2__0__5), .QB (\$dummy [173]), 
        .D (L0_2_L1_0_Wij_nx262), .CLK (CLK)) ;
    dff L0_2_L1_0_Wij_reg_Dout_6 (.Q (WindowDout_2__0__6), .QB (\$dummy [174]), 
        .D (L0_2_L1_0_Wij_nx272), .CLK (CLK)) ;
    dff L0_2_L1_0_Wij_reg_Dout_7 (.Q (WindowDout_2__0__7), .QB (\$dummy [175]), 
        .D (L0_2_L1_0_Wij_nx282), .CLK (CLK)) ;
    buf02 L0_2_L1_0_Wij_ix330 (.Y (L0_2_L1_0_Wij_nx331), .A (WindowWR)) ;
    buf02 L0_2_L1_0_Wij_ix332 (.Y (L0_2_L1_0_Wij_nx333), .A (WindowWR)) ;
    dff L0_2_L1_1_Fij_reg_Dout_0 (.Q (FilterDout_2__1__0), .QB (\$dummy [176]), 
        .D (L0_2_L1_1_Fij_nx212), .CLK (CLK)) ;
    nor02_2x L0_2_L1_1_Fij_ix297 (.Y (L0_2_L1_1_Fij_nx296), .A0 (RST), .A1 (
             L0_2_L1_1_Fij_nx331)) ;
    dff L0_2_L1_1_Fij_reg_Dout_1 (.Q (FilterDout_2__1__1), .QB (\$dummy [177]), 
        .D (L0_2_L1_1_Fij_nx222), .CLK (CLK)) ;
    dff L0_2_L1_1_Fij_reg_Dout_2 (.Q (FilterDout_2__1__2), .QB (\$dummy [178]), 
        .D (L0_2_L1_1_Fij_nx232), .CLK (CLK)) ;
    dff L0_2_L1_1_Fij_reg_Dout_3 (.Q (FilterDout_2__1__3), .QB (\$dummy [179]), 
        .D (L0_2_L1_1_Fij_nx242), .CLK (CLK)) ;
    dff L0_2_L1_1_Fij_reg_Dout_4 (.Q (FilterDout_2__1__4), .QB (\$dummy [180]), 
        .D (L0_2_L1_1_Fij_nx252), .CLK (CLK)) ;
    dff L0_2_L1_1_Fij_reg_Dout_5 (.Q (FilterDout_2__1__5), .QB (\$dummy [181]), 
        .D (L0_2_L1_1_Fij_nx262), .CLK (CLK)) ;
    dff L0_2_L1_1_Fij_reg_Dout_6 (.Q (FilterDout_2__1__6), .QB (\$dummy [182]), 
        .D (L0_2_L1_1_Fij_nx272), .CLK (CLK)) ;
    dff L0_2_L1_1_Fij_reg_Dout_7 (.Q (FilterDout_2__1__7), .QB (\$dummy [183]), 
        .D (L0_2_L1_1_Fij_nx282), .CLK (CLK)) ;
    buf02 L0_2_L1_1_Fij_ix330 (.Y (L0_2_L1_1_Fij_nx331), .A (FilterWR)) ;
    buf02 L0_2_L1_1_Fij_ix332 (.Y (L0_2_L1_1_Fij_nx333), .A (FilterWR)) ;
    dff L0_2_L1_1_Wij_reg_Dout_0 (.Q (WindowDout_2__1__0), .QB (\$dummy [184]), 
        .D (L0_2_L1_1_Wij_nx212), .CLK (CLK)) ;
    nor02_2x L0_2_L1_1_Wij_ix297 (.Y (L0_2_L1_1_Wij_nx296), .A0 (RST), .A1 (
             L0_2_L1_1_Wij_nx331)) ;
    dff L0_2_L1_1_Wij_reg_Dout_1 (.Q (WindowDout_2__1__1), .QB (\$dummy [185]), 
        .D (L0_2_L1_1_Wij_nx222), .CLK (CLK)) ;
    dff L0_2_L1_1_Wij_reg_Dout_2 (.Q (WindowDout_2__1__2), .QB (\$dummy [186]), 
        .D (L0_2_L1_1_Wij_nx232), .CLK (CLK)) ;
    dff L0_2_L1_1_Wij_reg_Dout_3 (.Q (WindowDout_2__1__3), .QB (\$dummy [187]), 
        .D (L0_2_L1_1_Wij_nx242), .CLK (CLK)) ;
    dff L0_2_L1_1_Wij_reg_Dout_4 (.Q (WindowDout_2__1__4), .QB (\$dummy [188]), 
        .D (L0_2_L1_1_Wij_nx252), .CLK (CLK)) ;
    dff L0_2_L1_1_Wij_reg_Dout_5 (.Q (WindowDout_2__1__5), .QB (\$dummy [189]), 
        .D (L0_2_L1_1_Wij_nx262), .CLK (CLK)) ;
    dff L0_2_L1_1_Wij_reg_Dout_6 (.Q (WindowDout_2__1__6), .QB (\$dummy [190]), 
        .D (L0_2_L1_1_Wij_nx272), .CLK (CLK)) ;
    dff L0_2_L1_1_Wij_reg_Dout_7 (.Q (WindowDout_2__1__7), .QB (\$dummy [191]), 
        .D (L0_2_L1_1_Wij_nx282), .CLK (CLK)) ;
    buf02 L0_2_L1_1_Wij_ix330 (.Y (L0_2_L1_1_Wij_nx331), .A (WindowWR)) ;
    buf02 L0_2_L1_1_Wij_ix332 (.Y (L0_2_L1_1_Wij_nx333), .A (WindowWR)) ;
    dff L0_2_L1_2_Fij_reg_Dout_0 (.Q (FilterDout_2__2__0), .QB (\$dummy [192]), 
        .D (L0_2_L1_2_Fij_nx212), .CLK (CLK)) ;
    nor02_2x L0_2_L1_2_Fij_ix297 (.Y (L0_2_L1_2_Fij_nx296), .A0 (RST), .A1 (
             L0_2_L1_2_Fij_nx331)) ;
    dff L0_2_L1_2_Fij_reg_Dout_1 (.Q (FilterDout_2__2__1), .QB (\$dummy [193]), 
        .D (L0_2_L1_2_Fij_nx222), .CLK (CLK)) ;
    dff L0_2_L1_2_Fij_reg_Dout_2 (.Q (FilterDout_2__2__2), .QB (\$dummy [194]), 
        .D (L0_2_L1_2_Fij_nx232), .CLK (CLK)) ;
    dff L0_2_L1_2_Fij_reg_Dout_3 (.Q (FilterDout_2__2__3), .QB (\$dummy [195]), 
        .D (L0_2_L1_2_Fij_nx242), .CLK (CLK)) ;
    dff L0_2_L1_2_Fij_reg_Dout_4 (.Q (FilterDout_2__2__4), .QB (\$dummy [196]), 
        .D (L0_2_L1_2_Fij_nx252), .CLK (CLK)) ;
    dff L0_2_L1_2_Fij_reg_Dout_5 (.Q (FilterDout_2__2__5), .QB (\$dummy [197]), 
        .D (L0_2_L1_2_Fij_nx262), .CLK (CLK)) ;
    dff L0_2_L1_2_Fij_reg_Dout_6 (.Q (FilterDout_2__2__6), .QB (\$dummy [198]), 
        .D (L0_2_L1_2_Fij_nx272), .CLK (CLK)) ;
    dff L0_2_L1_2_Fij_reg_Dout_7 (.Q (FilterDout_2__2__7), .QB (\$dummy [199]), 
        .D (L0_2_L1_2_Fij_nx282), .CLK (CLK)) ;
    buf02 L0_2_L1_2_Fij_ix330 (.Y (L0_2_L1_2_Fij_nx331), .A (FilterWR)) ;
    buf02 L0_2_L1_2_Fij_ix332 (.Y (L0_2_L1_2_Fij_nx333), .A (FilterWR)) ;
    dff L0_2_L1_2_Wij_reg_Dout_0 (.Q (WindowDout_2__2__0), .QB (\$dummy [200]), 
        .D (L0_2_L1_2_Wij_nx212), .CLK (CLK)) ;
    nor02_2x L0_2_L1_2_Wij_ix297 (.Y (L0_2_L1_2_Wij_nx296), .A0 (RST), .A1 (
             L0_2_L1_2_Wij_nx331)) ;
    dff L0_2_L1_2_Wij_reg_Dout_1 (.Q (WindowDout_2__2__1), .QB (\$dummy [201]), 
        .D (L0_2_L1_2_Wij_nx222), .CLK (CLK)) ;
    dff L0_2_L1_2_Wij_reg_Dout_2 (.Q (WindowDout_2__2__2), .QB (\$dummy [202]), 
        .D (L0_2_L1_2_Wij_nx232), .CLK (CLK)) ;
    dff L0_2_L1_2_Wij_reg_Dout_3 (.Q (WindowDout_2__2__3), .QB (\$dummy [203]), 
        .D (L0_2_L1_2_Wij_nx242), .CLK (CLK)) ;
    dff L0_2_L1_2_Wij_reg_Dout_4 (.Q (WindowDout_2__2__4), .QB (\$dummy [204]), 
        .D (L0_2_L1_2_Wij_nx252), .CLK (CLK)) ;
    dff L0_2_L1_2_Wij_reg_Dout_5 (.Q (WindowDout_2__2__5), .QB (\$dummy [205]), 
        .D (L0_2_L1_2_Wij_nx262), .CLK (CLK)) ;
    dff L0_2_L1_2_Wij_reg_Dout_6 (.Q (WindowDout_2__2__6), .QB (\$dummy [206]), 
        .D (L0_2_L1_2_Wij_nx272), .CLK (CLK)) ;
    dff L0_2_L1_2_Wij_reg_Dout_7 (.Q (WindowDout_2__2__7), .QB (\$dummy [207]), 
        .D (L0_2_L1_2_Wij_nx282), .CLK (CLK)) ;
    buf02 L0_2_L1_2_Wij_ix330 (.Y (L0_2_L1_2_Wij_nx331), .A (WindowWR)) ;
    buf02 L0_2_L1_2_Wij_ix332 (.Y (L0_2_L1_2_Wij_nx333), .A (WindowWR)) ;
    dff L0_2_L1_3_Fij_reg_Dout_0 (.Q (FilterDout_2__3__0), .QB (\$dummy [208]), 
        .D (L0_2_L1_3_Fij_nx212), .CLK (CLK)) ;
    nor02_2x L0_2_L1_3_Fij_ix297 (.Y (L0_2_L1_3_Fij_nx296), .A0 (RST), .A1 (
             L0_2_L1_3_Fij_nx331)) ;
    dff L0_2_L1_3_Fij_reg_Dout_1 (.Q (FilterDout_2__3__1), .QB (\$dummy [209]), 
        .D (L0_2_L1_3_Fij_nx222), .CLK (CLK)) ;
    dff L0_2_L1_3_Fij_reg_Dout_2 (.Q (FilterDout_2__3__2), .QB (\$dummy [210]), 
        .D (L0_2_L1_3_Fij_nx232), .CLK (CLK)) ;
    dff L0_2_L1_3_Fij_reg_Dout_3 (.Q (FilterDout_2__3__3), .QB (\$dummy [211]), 
        .D (L0_2_L1_3_Fij_nx242), .CLK (CLK)) ;
    dff L0_2_L1_3_Fij_reg_Dout_4 (.Q (FilterDout_2__3__4), .QB (\$dummy [212]), 
        .D (L0_2_L1_3_Fij_nx252), .CLK (CLK)) ;
    dff L0_2_L1_3_Fij_reg_Dout_5 (.Q (FilterDout_2__3__5), .QB (\$dummy [213]), 
        .D (L0_2_L1_3_Fij_nx262), .CLK (CLK)) ;
    dff L0_2_L1_3_Fij_reg_Dout_6 (.Q (FilterDout_2__3__6), .QB (\$dummy [214]), 
        .D (L0_2_L1_3_Fij_nx272), .CLK (CLK)) ;
    dff L0_2_L1_3_Fij_reg_Dout_7 (.Q (FilterDout_2__3__7), .QB (\$dummy [215]), 
        .D (L0_2_L1_3_Fij_nx282), .CLK (CLK)) ;
    buf02 L0_2_L1_3_Fij_ix330 (.Y (L0_2_L1_3_Fij_nx331), .A (EN_dup_1279)) ;
    buf02 L0_2_L1_3_Fij_ix332 (.Y (L0_2_L1_3_Fij_nx333), .A (EN_dup_1279)) ;
    dff L0_2_L1_3_Wij_reg_Dout_0 (.Q (WindowDout_2__3__0), .QB (\$dummy [216]), 
        .D (L0_2_L1_3_Wij_nx212), .CLK (CLK)) ;
    nor02_2x L0_2_L1_3_Wij_ix297 (.Y (L0_2_L1_3_Wij_nx296), .A0 (RST), .A1 (
             L0_2_L1_3_Wij_nx331)) ;
    dff L0_2_L1_3_Wij_reg_Dout_1 (.Q (WindowDout_2__3__1), .QB (\$dummy [217]), 
        .D (L0_2_L1_3_Wij_nx222), .CLK (CLK)) ;
    dff L0_2_L1_3_Wij_reg_Dout_2 (.Q (WindowDout_2__3__2), .QB (\$dummy [218]), 
        .D (L0_2_L1_3_Wij_nx232), .CLK (CLK)) ;
    dff L0_2_L1_3_Wij_reg_Dout_3 (.Q (WindowDout_2__3__3), .QB (\$dummy [219]), 
        .D (L0_2_L1_3_Wij_nx242), .CLK (CLK)) ;
    dff L0_2_L1_3_Wij_reg_Dout_4 (.Q (WindowDout_2__3__4), .QB (\$dummy [220]), 
        .D (L0_2_L1_3_Wij_nx252), .CLK (CLK)) ;
    dff L0_2_L1_3_Wij_reg_Dout_5 (.Q (WindowDout_2__3__5), .QB (\$dummy [221]), 
        .D (L0_2_L1_3_Wij_nx262), .CLK (CLK)) ;
    dff L0_2_L1_3_Wij_reg_Dout_6 (.Q (WindowDout_2__3__6), .QB (\$dummy [222]), 
        .D (L0_2_L1_3_Wij_nx272), .CLK (CLK)) ;
    dff L0_2_L1_3_Wij_reg_Dout_7 (.Q (WindowDout_2__3__7), .QB (\$dummy [223]), 
        .D (L0_2_L1_3_Wij_nx282), .CLK (CLK)) ;
    buf02 L0_2_L1_3_Wij_ix330 (.Y (L0_2_L1_3_Wij_nx331), .A (EN_dup_1290)) ;
    buf02 L0_2_L1_3_Wij_ix332 (.Y (L0_2_L1_3_Wij_nx333), .A (EN_dup_1290)) ;
    dff L0_2_L1_4_Fij_reg_Dout_0 (.Q (FilterDout_2__4__0), .QB (\$dummy [224]), 
        .D (L0_2_L1_4_Fij_nx212), .CLK (CLK)) ;
    nor02_2x L0_2_L1_4_Fij_ix297 (.Y (L0_2_L1_4_Fij_nx296), .A0 (RST), .A1 (
             L0_2_L1_4_Fij_nx331)) ;
    dff L0_2_L1_4_Fij_reg_Dout_1 (.Q (FilterDout_2__4__1), .QB (\$dummy [225]), 
        .D (L0_2_L1_4_Fij_nx222), .CLK (CLK)) ;
    dff L0_2_L1_4_Fij_reg_Dout_2 (.Q (FilterDout_2__4__2), .QB (\$dummy [226]), 
        .D (L0_2_L1_4_Fij_nx232), .CLK (CLK)) ;
    dff L0_2_L1_4_Fij_reg_Dout_3 (.Q (FilterDout_2__4__3), .QB (\$dummy [227]), 
        .D (L0_2_L1_4_Fij_nx242), .CLK (CLK)) ;
    dff L0_2_L1_4_Fij_reg_Dout_4 (.Q (FilterDout_2__4__4), .QB (\$dummy [228]), 
        .D (L0_2_L1_4_Fij_nx252), .CLK (CLK)) ;
    dff L0_2_L1_4_Fij_reg_Dout_5 (.Q (FilterDout_2__4__5), .QB (\$dummy [229]), 
        .D (L0_2_L1_4_Fij_nx262), .CLK (CLK)) ;
    dff L0_2_L1_4_Fij_reg_Dout_6 (.Q (FilterDout_2__4__6), .QB (\$dummy [230]), 
        .D (L0_2_L1_4_Fij_nx272), .CLK (CLK)) ;
    dff L0_2_L1_4_Fij_reg_Dout_7 (.Q (FilterDout_2__4__7), .QB (\$dummy [231]), 
        .D (L0_2_L1_4_Fij_nx282), .CLK (CLK)) ;
    buf02 L0_2_L1_4_Fij_ix330 (.Y (L0_2_L1_4_Fij_nx331), .A (EN_dup_1279)) ;
    buf02 L0_2_L1_4_Fij_ix332 (.Y (L0_2_L1_4_Fij_nx333), .A (EN_dup_1279)) ;
    dff L0_2_L1_4_Wij_reg_Dout_0 (.Q (WindowDout_2__4__0), .QB (\$dummy [232]), 
        .D (L0_2_L1_4_Wij_nx212), .CLK (CLK)) ;
    nor02_2x L0_2_L1_4_Wij_ix297 (.Y (L0_2_L1_4_Wij_nx296), .A0 (RST), .A1 (
             L0_2_L1_4_Wij_nx331)) ;
    dff L0_2_L1_4_Wij_reg_Dout_1 (.Q (WindowDout_2__4__1), .QB (\$dummy [233]), 
        .D (L0_2_L1_4_Wij_nx222), .CLK (CLK)) ;
    dff L0_2_L1_4_Wij_reg_Dout_2 (.Q (WindowDout_2__4__2), .QB (\$dummy [234]), 
        .D (L0_2_L1_4_Wij_nx232), .CLK (CLK)) ;
    dff L0_2_L1_4_Wij_reg_Dout_3 (.Q (WindowDout_2__4__3), .QB (\$dummy [235]), 
        .D (L0_2_L1_4_Wij_nx242), .CLK (CLK)) ;
    dff L0_2_L1_4_Wij_reg_Dout_4 (.Q (WindowDout_2__4__4), .QB (\$dummy [236]), 
        .D (L0_2_L1_4_Wij_nx252), .CLK (CLK)) ;
    dff L0_2_L1_4_Wij_reg_Dout_5 (.Q (WindowDout_2__4__5), .QB (\$dummy [237]), 
        .D (L0_2_L1_4_Wij_nx262), .CLK (CLK)) ;
    dff L0_2_L1_4_Wij_reg_Dout_6 (.Q (WindowDout_2__4__6), .QB (\$dummy [238]), 
        .D (L0_2_L1_4_Wij_nx272), .CLK (CLK)) ;
    dff L0_2_L1_4_Wij_reg_Dout_7 (.Q (WindowDout_2__4__7), .QB (\$dummy [239]), 
        .D (L0_2_L1_4_Wij_nx282), .CLK (CLK)) ;
    buf02 L0_2_L1_4_Wij_ix330 (.Y (L0_2_L1_4_Wij_nx331), .A (EN_dup_1290)) ;
    buf02 L0_2_L1_4_Wij_ix332 (.Y (L0_2_L1_4_Wij_nx333), .A (EN_dup_1290)) ;
    dff L0_3_L1_0_Fij_reg_Dout_0 (.Q (FilterDout_3__0__0), .QB (\$dummy [240]), 
        .D (L0_3_L1_0_Fij_nx212), .CLK (CLK)) ;
    nor02_2x L0_3_L1_0_Fij_ix297 (.Y (L0_3_L1_0_Fij_nx296), .A0 (RST), .A1 (
             L0_3_L1_0_Fij_nx331)) ;
    dff L0_3_L1_0_Fij_reg_Dout_1 (.Q (FilterDout_3__0__1), .QB (\$dummy [241]), 
        .D (L0_3_L1_0_Fij_nx222), .CLK (CLK)) ;
    dff L0_3_L1_0_Fij_reg_Dout_2 (.Q (FilterDout_3__0__2), .QB (\$dummy [242]), 
        .D (L0_3_L1_0_Fij_nx232), .CLK (CLK)) ;
    dff L0_3_L1_0_Fij_reg_Dout_3 (.Q (FilterDout_3__0__3), .QB (\$dummy [243]), 
        .D (L0_3_L1_0_Fij_nx242), .CLK (CLK)) ;
    dff L0_3_L1_0_Fij_reg_Dout_4 (.Q (FilterDout_3__0__4), .QB (\$dummy [244]), 
        .D (L0_3_L1_0_Fij_nx252), .CLK (CLK)) ;
    dff L0_3_L1_0_Fij_reg_Dout_5 (.Q (FilterDout_3__0__5), .QB (\$dummy [245]), 
        .D (L0_3_L1_0_Fij_nx262), .CLK (CLK)) ;
    dff L0_3_L1_0_Fij_reg_Dout_6 (.Q (FilterDout_3__0__6), .QB (\$dummy [246]), 
        .D (L0_3_L1_0_Fij_nx272), .CLK (CLK)) ;
    dff L0_3_L1_0_Fij_reg_Dout_7 (.Q (FilterDout_3__0__7), .QB (\$dummy [247]), 
        .D (L0_3_L1_0_Fij_nx282), .CLK (CLK)) ;
    buf02 L0_3_L1_0_Fij_ix330 (.Y (L0_3_L1_0_Fij_nx331), .A (FilterWR)) ;
    buf02 L0_3_L1_0_Fij_ix332 (.Y (L0_3_L1_0_Fij_nx333), .A (FilterWR)) ;
    dff L0_3_L1_0_Wij_reg_Dout_0 (.Q (WindowDout_3__0__0), .QB (\$dummy [248]), 
        .D (L0_3_L1_0_Wij_nx212), .CLK (CLK)) ;
    nor02_2x L0_3_L1_0_Wij_ix297 (.Y (L0_3_L1_0_Wij_nx296), .A0 (RST), .A1 (
             L0_3_L1_0_Wij_nx331)) ;
    dff L0_3_L1_0_Wij_reg_Dout_1 (.Q (WindowDout_3__0__1), .QB (\$dummy [249]), 
        .D (L0_3_L1_0_Wij_nx222), .CLK (CLK)) ;
    dff L0_3_L1_0_Wij_reg_Dout_2 (.Q (WindowDout_3__0__2), .QB (\$dummy [250]), 
        .D (L0_3_L1_0_Wij_nx232), .CLK (CLK)) ;
    dff L0_3_L1_0_Wij_reg_Dout_3 (.Q (WindowDout_3__0__3), .QB (\$dummy [251]), 
        .D (L0_3_L1_0_Wij_nx242), .CLK (CLK)) ;
    dff L0_3_L1_0_Wij_reg_Dout_4 (.Q (WindowDout_3__0__4), .QB (\$dummy [252]), 
        .D (L0_3_L1_0_Wij_nx252), .CLK (CLK)) ;
    dff L0_3_L1_0_Wij_reg_Dout_5 (.Q (WindowDout_3__0__5), .QB (\$dummy [253]), 
        .D (L0_3_L1_0_Wij_nx262), .CLK (CLK)) ;
    dff L0_3_L1_0_Wij_reg_Dout_6 (.Q (WindowDout_3__0__6), .QB (\$dummy [254]), 
        .D (L0_3_L1_0_Wij_nx272), .CLK (CLK)) ;
    dff L0_3_L1_0_Wij_reg_Dout_7 (.Q (WindowDout_3__0__7), .QB (\$dummy [255]), 
        .D (L0_3_L1_0_Wij_nx282), .CLK (CLK)) ;
    buf02 L0_3_L1_0_Wij_ix330 (.Y (L0_3_L1_0_Wij_nx331), .A (WindowWR)) ;
    buf02 L0_3_L1_0_Wij_ix332 (.Y (L0_3_L1_0_Wij_nx333), .A (WindowWR)) ;
    dff L0_3_L1_1_Fij_reg_Dout_0 (.Q (FilterDout_3__1__0), .QB (\$dummy [256]), 
        .D (L0_3_L1_1_Fij_nx212), .CLK (CLK)) ;
    nor02_2x L0_3_L1_1_Fij_ix297 (.Y (L0_3_L1_1_Fij_nx296), .A0 (RST), .A1 (
             L0_3_L1_1_Fij_nx331)) ;
    dff L0_3_L1_1_Fij_reg_Dout_1 (.Q (FilterDout_3__1__1), .QB (\$dummy [257]), 
        .D (L0_3_L1_1_Fij_nx222), .CLK (CLK)) ;
    dff L0_3_L1_1_Fij_reg_Dout_2 (.Q (FilterDout_3__1__2), .QB (\$dummy [258]), 
        .D (L0_3_L1_1_Fij_nx232), .CLK (CLK)) ;
    dff L0_3_L1_1_Fij_reg_Dout_3 (.Q (FilterDout_3__1__3), .QB (\$dummy [259]), 
        .D (L0_3_L1_1_Fij_nx242), .CLK (CLK)) ;
    dff L0_3_L1_1_Fij_reg_Dout_4 (.Q (FilterDout_3__1__4), .QB (\$dummy [260]), 
        .D (L0_3_L1_1_Fij_nx252), .CLK (CLK)) ;
    dff L0_3_L1_1_Fij_reg_Dout_5 (.Q (FilterDout_3__1__5), .QB (\$dummy [261]), 
        .D (L0_3_L1_1_Fij_nx262), .CLK (CLK)) ;
    dff L0_3_L1_1_Fij_reg_Dout_6 (.Q (FilterDout_3__1__6), .QB (\$dummy [262]), 
        .D (L0_3_L1_1_Fij_nx272), .CLK (CLK)) ;
    dff L0_3_L1_1_Fij_reg_Dout_7 (.Q (FilterDout_3__1__7), .QB (\$dummy [263]), 
        .D (L0_3_L1_1_Fij_nx282), .CLK (CLK)) ;
    buf02 L0_3_L1_1_Fij_ix330 (.Y (L0_3_L1_1_Fij_nx331), .A (FilterWR)) ;
    buf02 L0_3_L1_1_Fij_ix332 (.Y (L0_3_L1_1_Fij_nx333), .A (FilterWR)) ;
    dff L0_3_L1_1_Wij_reg_Dout_0 (.Q (WindowDout_3__1__0), .QB (\$dummy [264]), 
        .D (L0_3_L1_1_Wij_nx212), .CLK (CLK)) ;
    nor02_2x L0_3_L1_1_Wij_ix297 (.Y (L0_3_L1_1_Wij_nx296), .A0 (RST), .A1 (
             L0_3_L1_1_Wij_nx331)) ;
    dff L0_3_L1_1_Wij_reg_Dout_1 (.Q (WindowDout_3__1__1), .QB (\$dummy [265]), 
        .D (L0_3_L1_1_Wij_nx222), .CLK (CLK)) ;
    dff L0_3_L1_1_Wij_reg_Dout_2 (.Q (WindowDout_3__1__2), .QB (\$dummy [266]), 
        .D (L0_3_L1_1_Wij_nx232), .CLK (CLK)) ;
    dff L0_3_L1_1_Wij_reg_Dout_3 (.Q (WindowDout_3__1__3), .QB (\$dummy [267]), 
        .D (L0_3_L1_1_Wij_nx242), .CLK (CLK)) ;
    dff L0_3_L1_1_Wij_reg_Dout_4 (.Q (WindowDout_3__1__4), .QB (\$dummy [268]), 
        .D (L0_3_L1_1_Wij_nx252), .CLK (CLK)) ;
    dff L0_3_L1_1_Wij_reg_Dout_5 (.Q (WindowDout_3__1__5), .QB (\$dummy [269]), 
        .D (L0_3_L1_1_Wij_nx262), .CLK (CLK)) ;
    dff L0_3_L1_1_Wij_reg_Dout_6 (.Q (WindowDout_3__1__6), .QB (\$dummy [270]), 
        .D (L0_3_L1_1_Wij_nx272), .CLK (CLK)) ;
    dff L0_3_L1_1_Wij_reg_Dout_7 (.Q (WindowDout_3__1__7), .QB (\$dummy [271]), 
        .D (L0_3_L1_1_Wij_nx282), .CLK (CLK)) ;
    buf02 L0_3_L1_1_Wij_ix330 (.Y (L0_3_L1_1_Wij_nx331), .A (WindowWR)) ;
    buf02 L0_3_L1_1_Wij_ix332 (.Y (L0_3_L1_1_Wij_nx333), .A (WindowWR)) ;
    dff L0_3_L1_2_Fij_reg_Dout_0 (.Q (FilterDout_3__2__0), .QB (\$dummy [272]), 
        .D (L0_3_L1_2_Fij_nx212), .CLK (CLK)) ;
    nor02_2x L0_3_L1_2_Fij_ix297 (.Y (L0_3_L1_2_Fij_nx296), .A0 (RST), .A1 (
             L0_3_L1_2_Fij_nx331)) ;
    dff L0_3_L1_2_Fij_reg_Dout_1 (.Q (FilterDout_3__2__1), .QB (\$dummy [273]), 
        .D (L0_3_L1_2_Fij_nx222), .CLK (CLK)) ;
    dff L0_3_L1_2_Fij_reg_Dout_2 (.Q (FilterDout_3__2__2), .QB (\$dummy [274]), 
        .D (L0_3_L1_2_Fij_nx232), .CLK (CLK)) ;
    dff L0_3_L1_2_Fij_reg_Dout_3 (.Q (FilterDout_3__2__3), .QB (\$dummy [275]), 
        .D (L0_3_L1_2_Fij_nx242), .CLK (CLK)) ;
    dff L0_3_L1_2_Fij_reg_Dout_4 (.Q (FilterDout_3__2__4), .QB (\$dummy [276]), 
        .D (L0_3_L1_2_Fij_nx252), .CLK (CLK)) ;
    dff L0_3_L1_2_Fij_reg_Dout_5 (.Q (FilterDout_3__2__5), .QB (\$dummy [277]), 
        .D (L0_3_L1_2_Fij_nx262), .CLK (CLK)) ;
    dff L0_3_L1_2_Fij_reg_Dout_6 (.Q (FilterDout_3__2__6), .QB (\$dummy [278]), 
        .D (L0_3_L1_2_Fij_nx272), .CLK (CLK)) ;
    dff L0_3_L1_2_Fij_reg_Dout_7 (.Q (FilterDout_3__2__7), .QB (\$dummy [279]), 
        .D (L0_3_L1_2_Fij_nx282), .CLK (CLK)) ;
    buf02 L0_3_L1_2_Fij_ix330 (.Y (L0_3_L1_2_Fij_nx331), .A (FilterWR)) ;
    buf02 L0_3_L1_2_Fij_ix332 (.Y (L0_3_L1_2_Fij_nx333), .A (FilterWR)) ;
    dff L0_3_L1_2_Wij_reg_Dout_0 (.Q (WindowDout_3__2__0), .QB (\$dummy [280]), 
        .D (L0_3_L1_2_Wij_nx212), .CLK (CLK)) ;
    nor02_2x L0_3_L1_2_Wij_ix297 (.Y (L0_3_L1_2_Wij_nx296), .A0 (RST), .A1 (
             L0_3_L1_2_Wij_nx331)) ;
    dff L0_3_L1_2_Wij_reg_Dout_1 (.Q (WindowDout_3__2__1), .QB (\$dummy [281]), 
        .D (L0_3_L1_2_Wij_nx222), .CLK (CLK)) ;
    dff L0_3_L1_2_Wij_reg_Dout_2 (.Q (WindowDout_3__2__2), .QB (\$dummy [282]), 
        .D (L0_3_L1_2_Wij_nx232), .CLK (CLK)) ;
    dff L0_3_L1_2_Wij_reg_Dout_3 (.Q (WindowDout_3__2__3), .QB (\$dummy [283]), 
        .D (L0_3_L1_2_Wij_nx242), .CLK (CLK)) ;
    dff L0_3_L1_2_Wij_reg_Dout_4 (.Q (WindowDout_3__2__4), .QB (\$dummy [284]), 
        .D (L0_3_L1_2_Wij_nx252), .CLK (CLK)) ;
    dff L0_3_L1_2_Wij_reg_Dout_5 (.Q (WindowDout_3__2__5), .QB (\$dummy [285]), 
        .D (L0_3_L1_2_Wij_nx262), .CLK (CLK)) ;
    dff L0_3_L1_2_Wij_reg_Dout_6 (.Q (WindowDout_3__2__6), .QB (\$dummy [286]), 
        .D (L0_3_L1_2_Wij_nx272), .CLK (CLK)) ;
    dff L0_3_L1_2_Wij_reg_Dout_7 (.Q (WindowDout_3__2__7), .QB (\$dummy [287]), 
        .D (L0_3_L1_2_Wij_nx282), .CLK (CLK)) ;
    buf02 L0_3_L1_2_Wij_ix330 (.Y (L0_3_L1_2_Wij_nx331), .A (WindowWR)) ;
    buf02 L0_3_L1_2_Wij_ix332 (.Y (L0_3_L1_2_Wij_nx333), .A (WindowWR)) ;
    dff L0_3_L1_3_Fij_reg_Dout_0 (.Q (FilterDout_3__3__0), .QB (\$dummy [288]), 
        .D (L0_3_L1_3_Fij_nx212), .CLK (CLK)) ;
    nor02_2x L0_3_L1_3_Fij_ix297 (.Y (L0_3_L1_3_Fij_nx296), .A0 (RST), .A1 (
             L0_3_L1_3_Fij_nx331)) ;
    dff L0_3_L1_3_Fij_reg_Dout_1 (.Q (FilterDout_3__3__1), .QB (\$dummy [289]), 
        .D (L0_3_L1_3_Fij_nx222), .CLK (CLK)) ;
    dff L0_3_L1_3_Fij_reg_Dout_2 (.Q (FilterDout_3__3__2), .QB (\$dummy [290]), 
        .D (L0_3_L1_3_Fij_nx232), .CLK (CLK)) ;
    dff L0_3_L1_3_Fij_reg_Dout_3 (.Q (FilterDout_3__3__3), .QB (\$dummy [291]), 
        .D (L0_3_L1_3_Fij_nx242), .CLK (CLK)) ;
    dff L0_3_L1_3_Fij_reg_Dout_4 (.Q (FilterDout_3__3__4), .QB (\$dummy [292]), 
        .D (L0_3_L1_3_Fij_nx252), .CLK (CLK)) ;
    dff L0_3_L1_3_Fij_reg_Dout_5 (.Q (FilterDout_3__3__5), .QB (\$dummy [293]), 
        .D (L0_3_L1_3_Fij_nx262), .CLK (CLK)) ;
    dff L0_3_L1_3_Fij_reg_Dout_6 (.Q (FilterDout_3__3__6), .QB (\$dummy [294]), 
        .D (L0_3_L1_3_Fij_nx272), .CLK (CLK)) ;
    dff L0_3_L1_3_Fij_reg_Dout_7 (.Q (FilterDout_3__3__7), .QB (\$dummy [295]), 
        .D (L0_3_L1_3_Fij_nx282), .CLK (CLK)) ;
    buf02 L0_3_L1_3_Fij_ix330 (.Y (L0_3_L1_3_Fij_nx331), .A (EN_dup_1279)) ;
    buf02 L0_3_L1_3_Fij_ix332 (.Y (L0_3_L1_3_Fij_nx333), .A (EN_dup_1279)) ;
    dff L0_3_L1_3_Wij_reg_Dout_0 (.Q (WindowDout_3__3__0), .QB (\$dummy [296]), 
        .D (L0_3_L1_3_Wij_nx212), .CLK (CLK)) ;
    nor02_2x L0_3_L1_3_Wij_ix297 (.Y (L0_3_L1_3_Wij_nx296), .A0 (RST), .A1 (
             L0_3_L1_3_Wij_nx331)) ;
    dff L0_3_L1_3_Wij_reg_Dout_1 (.Q (WindowDout_3__3__1), .QB (\$dummy [297]), 
        .D (L0_3_L1_3_Wij_nx222), .CLK (CLK)) ;
    dff L0_3_L1_3_Wij_reg_Dout_2 (.Q (WindowDout_3__3__2), .QB (\$dummy [298]), 
        .D (L0_3_L1_3_Wij_nx232), .CLK (CLK)) ;
    dff L0_3_L1_3_Wij_reg_Dout_3 (.Q (WindowDout_3__3__3), .QB (\$dummy [299]), 
        .D (L0_3_L1_3_Wij_nx242), .CLK (CLK)) ;
    dff L0_3_L1_3_Wij_reg_Dout_4 (.Q (WindowDout_3__3__4), .QB (\$dummy [300]), 
        .D (L0_3_L1_3_Wij_nx252), .CLK (CLK)) ;
    dff L0_3_L1_3_Wij_reg_Dout_5 (.Q (WindowDout_3__3__5), .QB (\$dummy [301]), 
        .D (L0_3_L1_3_Wij_nx262), .CLK (CLK)) ;
    dff L0_3_L1_3_Wij_reg_Dout_6 (.Q (WindowDout_3__3__6), .QB (\$dummy [302]), 
        .D (L0_3_L1_3_Wij_nx272), .CLK (CLK)) ;
    dff L0_3_L1_3_Wij_reg_Dout_7 (.Q (WindowDout_3__3__7), .QB (\$dummy [303]), 
        .D (L0_3_L1_3_Wij_nx282), .CLK (CLK)) ;
    buf02 L0_3_L1_3_Wij_ix330 (.Y (L0_3_L1_3_Wij_nx331), .A (EN_dup_1290)) ;
    buf02 L0_3_L1_3_Wij_ix332 (.Y (L0_3_L1_3_Wij_nx333), .A (EN_dup_1290)) ;
    dff L0_3_L1_4_Fij_reg_Dout_0 (.Q (FilterDout_3__4__0), .QB (\$dummy [304]), 
        .D (L0_3_L1_4_Fij_nx212), .CLK (CLK)) ;
    nor02_2x L0_3_L1_4_Fij_ix297 (.Y (L0_3_L1_4_Fij_nx296), .A0 (RST), .A1 (
             L0_3_L1_4_Fij_nx331)) ;
    dff L0_3_L1_4_Fij_reg_Dout_1 (.Q (FilterDout_3__4__1), .QB (\$dummy [305]), 
        .D (L0_3_L1_4_Fij_nx222), .CLK (CLK)) ;
    dff L0_3_L1_4_Fij_reg_Dout_2 (.Q (FilterDout_3__4__2), .QB (\$dummy [306]), 
        .D (L0_3_L1_4_Fij_nx232), .CLK (CLK)) ;
    dff L0_3_L1_4_Fij_reg_Dout_3 (.Q (FilterDout_3__4__3), .QB (\$dummy [307]), 
        .D (L0_3_L1_4_Fij_nx242), .CLK (CLK)) ;
    dff L0_3_L1_4_Fij_reg_Dout_4 (.Q (FilterDout_3__4__4), .QB (\$dummy [308]), 
        .D (L0_3_L1_4_Fij_nx252), .CLK (CLK)) ;
    dff L0_3_L1_4_Fij_reg_Dout_5 (.Q (FilterDout_3__4__5), .QB (\$dummy [309]), 
        .D (L0_3_L1_4_Fij_nx262), .CLK (CLK)) ;
    dff L0_3_L1_4_Fij_reg_Dout_6 (.Q (FilterDout_3__4__6), .QB (\$dummy [310]), 
        .D (L0_3_L1_4_Fij_nx272), .CLK (CLK)) ;
    dff L0_3_L1_4_Fij_reg_Dout_7 (.Q (FilterDout_3__4__7), .QB (\$dummy [311]), 
        .D (L0_3_L1_4_Fij_nx282), .CLK (CLK)) ;
    buf02 L0_3_L1_4_Fij_ix330 (.Y (L0_3_L1_4_Fij_nx331), .A (EN_dup_1411)) ;
    buf02 L0_3_L1_4_Fij_ix332 (.Y (L0_3_L1_4_Fij_nx333), .A (EN_dup_1411)) ;
    dff L0_3_L1_4_Wij_reg_Dout_0 (.Q (WindowDout_3__4__0), .QB (\$dummy [312]), 
        .D (L0_3_L1_4_Wij_nx212), .CLK (CLK)) ;
    nor02_2x L0_3_L1_4_Wij_ix297 (.Y (L0_3_L1_4_Wij_nx296), .A0 (RST), .A1 (
             L0_3_L1_4_Wij_nx331)) ;
    dff L0_3_L1_4_Wij_reg_Dout_1 (.Q (WindowDout_3__4__1), .QB (\$dummy [313]), 
        .D (L0_3_L1_4_Wij_nx222), .CLK (CLK)) ;
    dff L0_3_L1_4_Wij_reg_Dout_2 (.Q (WindowDout_3__4__2), .QB (\$dummy [314]), 
        .D (L0_3_L1_4_Wij_nx232), .CLK (CLK)) ;
    dff L0_3_L1_4_Wij_reg_Dout_3 (.Q (WindowDout_3__4__3), .QB (\$dummy [315]), 
        .D (L0_3_L1_4_Wij_nx242), .CLK (CLK)) ;
    dff L0_3_L1_4_Wij_reg_Dout_4 (.Q (WindowDout_3__4__4), .QB (\$dummy [316]), 
        .D (L0_3_L1_4_Wij_nx252), .CLK (CLK)) ;
    dff L0_3_L1_4_Wij_reg_Dout_5 (.Q (WindowDout_3__4__5), .QB (\$dummy [317]), 
        .D (L0_3_L1_4_Wij_nx262), .CLK (CLK)) ;
    dff L0_3_L1_4_Wij_reg_Dout_6 (.Q (WindowDout_3__4__6), .QB (\$dummy [318]), 
        .D (L0_3_L1_4_Wij_nx272), .CLK (CLK)) ;
    dff L0_3_L1_4_Wij_reg_Dout_7 (.Q (WindowDout_3__4__7), .QB (\$dummy [319]), 
        .D (L0_3_L1_4_Wij_nx282), .CLK (CLK)) ;
    buf02 L0_3_L1_4_Wij_ix330 (.Y (L0_3_L1_4_Wij_nx331), .A (EN_dup_1422)) ;
    buf02 L0_3_L1_4_Wij_ix332 (.Y (L0_3_L1_4_Wij_nx333), .A (EN_dup_1422)) ;
    dff L0_4_L1_0_Fij_reg_Dout_0 (.Q (FilterDout_4__0__0), .QB (\$dummy [320]), 
        .D (L0_4_L1_0_Fij_nx212), .CLK (CLK)) ;
    nor02_2x L0_4_L1_0_Fij_ix297 (.Y (L0_4_L1_0_Fij_nx296), .A0 (RST), .A1 (
             L0_4_L1_0_Fij_nx331)) ;
    dff L0_4_L1_0_Fij_reg_Dout_1 (.Q (FilterDout_4__0__1), .QB (\$dummy [321]), 
        .D (L0_4_L1_0_Fij_nx222), .CLK (CLK)) ;
    dff L0_4_L1_0_Fij_reg_Dout_2 (.Q (FilterDout_4__0__2), .QB (\$dummy [322]), 
        .D (L0_4_L1_0_Fij_nx232), .CLK (CLK)) ;
    dff L0_4_L1_0_Fij_reg_Dout_3 (.Q (FilterDout_4__0__3), .QB (\$dummy [323]), 
        .D (L0_4_L1_0_Fij_nx242), .CLK (CLK)) ;
    dff L0_4_L1_0_Fij_reg_Dout_4 (.Q (FilterDout_4__0__4), .QB (\$dummy [324]), 
        .D (L0_4_L1_0_Fij_nx252), .CLK (CLK)) ;
    dff L0_4_L1_0_Fij_reg_Dout_5 (.Q (FilterDout_4__0__5), .QB (\$dummy [325]), 
        .D (L0_4_L1_0_Fij_nx262), .CLK (CLK)) ;
    dff L0_4_L1_0_Fij_reg_Dout_6 (.Q (FilterDout_4__0__6), .QB (\$dummy [326]), 
        .D (L0_4_L1_0_Fij_nx272), .CLK (CLK)) ;
    dff L0_4_L1_0_Fij_reg_Dout_7 (.Q (FilterDout_4__0__7), .QB (\$dummy [327]), 
        .D (L0_4_L1_0_Fij_nx282), .CLK (CLK)) ;
    buf02 L0_4_L1_0_Fij_ix330 (.Y (L0_4_L1_0_Fij_nx331), .A (FilterWR)) ;
    buf02 L0_4_L1_0_Fij_ix332 (.Y (L0_4_L1_0_Fij_nx333), .A (FilterWR)) ;
    dff L0_4_L1_0_Wij_reg_Dout_0 (.Q (WindowDout_4__0__0), .QB (\$dummy [328]), 
        .D (L0_4_L1_0_Wij_nx212), .CLK (CLK)) ;
    nor02_2x L0_4_L1_0_Wij_ix297 (.Y (L0_4_L1_0_Wij_nx296), .A0 (RST), .A1 (
             L0_4_L1_0_Wij_nx331)) ;
    dff L0_4_L1_0_Wij_reg_Dout_1 (.Q (WindowDout_4__0__1), .QB (\$dummy [329]), 
        .D (L0_4_L1_0_Wij_nx222), .CLK (CLK)) ;
    dff L0_4_L1_0_Wij_reg_Dout_2 (.Q (WindowDout_4__0__2), .QB (\$dummy [330]), 
        .D (L0_4_L1_0_Wij_nx232), .CLK (CLK)) ;
    dff L0_4_L1_0_Wij_reg_Dout_3 (.Q (WindowDout_4__0__3), .QB (\$dummy [331]), 
        .D (L0_4_L1_0_Wij_nx242), .CLK (CLK)) ;
    dff L0_4_L1_0_Wij_reg_Dout_4 (.Q (WindowDout_4__0__4), .QB (\$dummy [332]), 
        .D (L0_4_L1_0_Wij_nx252), .CLK (CLK)) ;
    dff L0_4_L1_0_Wij_reg_Dout_5 (.Q (WindowDout_4__0__5), .QB (\$dummy [333]), 
        .D (L0_4_L1_0_Wij_nx262), .CLK (CLK)) ;
    dff L0_4_L1_0_Wij_reg_Dout_6 (.Q (WindowDout_4__0__6), .QB (\$dummy [334]), 
        .D (L0_4_L1_0_Wij_nx272), .CLK (CLK)) ;
    dff L0_4_L1_0_Wij_reg_Dout_7 (.Q (WindowDout_4__0__7), .QB (\$dummy [335]), 
        .D (L0_4_L1_0_Wij_nx282), .CLK (CLK)) ;
    buf02 L0_4_L1_0_Wij_ix330 (.Y (L0_4_L1_0_Wij_nx331), .A (WindowWR)) ;
    buf02 L0_4_L1_0_Wij_ix332 (.Y (L0_4_L1_0_Wij_nx333), .A (WindowWR)) ;
    dff L0_4_L1_1_Fij_reg_Dout_0 (.Q (FilterDout_4__1__0), .QB (\$dummy [336]), 
        .D (L0_4_L1_1_Fij_nx212), .CLK (CLK)) ;
    nor02_2x L0_4_L1_1_Fij_ix297 (.Y (L0_4_L1_1_Fij_nx296), .A0 (RST), .A1 (
             L0_4_L1_1_Fij_nx331)) ;
    dff L0_4_L1_1_Fij_reg_Dout_1 (.Q (FilterDout_4__1__1), .QB (\$dummy [337]), 
        .D (L0_4_L1_1_Fij_nx222), .CLK (CLK)) ;
    dff L0_4_L1_1_Fij_reg_Dout_2 (.Q (FilterDout_4__1__2), .QB (\$dummy [338]), 
        .D (L0_4_L1_1_Fij_nx232), .CLK (CLK)) ;
    dff L0_4_L1_1_Fij_reg_Dout_3 (.Q (FilterDout_4__1__3), .QB (\$dummy [339]), 
        .D (L0_4_L1_1_Fij_nx242), .CLK (CLK)) ;
    dff L0_4_L1_1_Fij_reg_Dout_4 (.Q (FilterDout_4__1__4), .QB (\$dummy [340]), 
        .D (L0_4_L1_1_Fij_nx252), .CLK (CLK)) ;
    dff L0_4_L1_1_Fij_reg_Dout_5 (.Q (FilterDout_4__1__5), .QB (\$dummy [341]), 
        .D (L0_4_L1_1_Fij_nx262), .CLK (CLK)) ;
    dff L0_4_L1_1_Fij_reg_Dout_6 (.Q (FilterDout_4__1__6), .QB (\$dummy [342]), 
        .D (L0_4_L1_1_Fij_nx272), .CLK (CLK)) ;
    dff L0_4_L1_1_Fij_reg_Dout_7 (.Q (FilterDout_4__1__7), .QB (\$dummy [343]), 
        .D (L0_4_L1_1_Fij_nx282), .CLK (CLK)) ;
    buf02 L0_4_L1_1_Fij_ix330 (.Y (L0_4_L1_1_Fij_nx331), .A (FilterWR)) ;
    buf02 L0_4_L1_1_Fij_ix332 (.Y (L0_4_L1_1_Fij_nx333), .A (FilterWR)) ;
    dff L0_4_L1_1_Wij_reg_Dout_0 (.Q (WindowDout_4__1__0), .QB (\$dummy [344]), 
        .D (L0_4_L1_1_Wij_nx212), .CLK (CLK)) ;
    nor02_2x L0_4_L1_1_Wij_ix297 (.Y (L0_4_L1_1_Wij_nx296), .A0 (RST), .A1 (
             L0_4_L1_1_Wij_nx331)) ;
    dff L0_4_L1_1_Wij_reg_Dout_1 (.Q (WindowDout_4__1__1), .QB (\$dummy [345]), 
        .D (L0_4_L1_1_Wij_nx222), .CLK (CLK)) ;
    dff L0_4_L1_1_Wij_reg_Dout_2 (.Q (WindowDout_4__1__2), .QB (\$dummy [346]), 
        .D (L0_4_L1_1_Wij_nx232), .CLK (CLK)) ;
    dff L0_4_L1_1_Wij_reg_Dout_3 (.Q (WindowDout_4__1__3), .QB (\$dummy [347]), 
        .D (L0_4_L1_1_Wij_nx242), .CLK (CLK)) ;
    dff L0_4_L1_1_Wij_reg_Dout_4 (.Q (WindowDout_4__1__4), .QB (\$dummy [348]), 
        .D (L0_4_L1_1_Wij_nx252), .CLK (CLK)) ;
    dff L0_4_L1_1_Wij_reg_Dout_5 (.Q (WindowDout_4__1__5), .QB (\$dummy [349]), 
        .D (L0_4_L1_1_Wij_nx262), .CLK (CLK)) ;
    dff L0_4_L1_1_Wij_reg_Dout_6 (.Q (WindowDout_4__1__6), .QB (\$dummy [350]), 
        .D (L0_4_L1_1_Wij_nx272), .CLK (CLK)) ;
    dff L0_4_L1_1_Wij_reg_Dout_7 (.Q (WindowDout_4__1__7), .QB (\$dummy [351]), 
        .D (L0_4_L1_1_Wij_nx282), .CLK (CLK)) ;
    buf02 L0_4_L1_1_Wij_ix330 (.Y (L0_4_L1_1_Wij_nx331), .A (WindowWR)) ;
    buf02 L0_4_L1_1_Wij_ix332 (.Y (L0_4_L1_1_Wij_nx333), .A (WindowWR)) ;
    dff L0_4_L1_2_Fij_reg_Dout_0 (.Q (FilterDout_4__2__0), .QB (\$dummy [352]), 
        .D (L0_4_L1_2_Fij_nx212), .CLK (CLK)) ;
    nor02_2x L0_4_L1_2_Fij_ix297 (.Y (L0_4_L1_2_Fij_nx296), .A0 (RST), .A1 (
             L0_4_L1_2_Fij_nx331)) ;
    dff L0_4_L1_2_Fij_reg_Dout_1 (.Q (FilterDout_4__2__1), .QB (\$dummy [353]), 
        .D (L0_4_L1_2_Fij_nx222), .CLK (CLK)) ;
    dff L0_4_L1_2_Fij_reg_Dout_2 (.Q (FilterDout_4__2__2), .QB (\$dummy [354]), 
        .D (L0_4_L1_2_Fij_nx232), .CLK (CLK)) ;
    dff L0_4_L1_2_Fij_reg_Dout_3 (.Q (FilterDout_4__2__3), .QB (\$dummy [355]), 
        .D (L0_4_L1_2_Fij_nx242), .CLK (CLK)) ;
    dff L0_4_L1_2_Fij_reg_Dout_4 (.Q (FilterDout_4__2__4), .QB (\$dummy [356]), 
        .D (L0_4_L1_2_Fij_nx252), .CLK (CLK)) ;
    dff L0_4_L1_2_Fij_reg_Dout_5 (.Q (FilterDout_4__2__5), .QB (\$dummy [357]), 
        .D (L0_4_L1_2_Fij_nx262), .CLK (CLK)) ;
    dff L0_4_L1_2_Fij_reg_Dout_6 (.Q (FilterDout_4__2__6), .QB (\$dummy [358]), 
        .D (L0_4_L1_2_Fij_nx272), .CLK (CLK)) ;
    dff L0_4_L1_2_Fij_reg_Dout_7 (.Q (FilterDout_4__2__7), .QB (\$dummy [359]), 
        .D (L0_4_L1_2_Fij_nx282), .CLK (CLK)) ;
    buf02 L0_4_L1_2_Fij_ix330 (.Y (L0_4_L1_2_Fij_nx331), .A (FilterWR)) ;
    buf02 L0_4_L1_2_Fij_ix332 (.Y (L0_4_L1_2_Fij_nx333), .A (FilterWR)) ;
    dff L0_4_L1_2_Wij_reg_Dout_0 (.Q (WindowDout_4__2__0), .QB (\$dummy [360]), 
        .D (L0_4_L1_2_Wij_nx212), .CLK (CLK)) ;
    nor02_2x L0_4_L1_2_Wij_ix297 (.Y (L0_4_L1_2_Wij_nx296), .A0 (RST), .A1 (
             L0_4_L1_2_Wij_nx331)) ;
    dff L0_4_L1_2_Wij_reg_Dout_1 (.Q (WindowDout_4__2__1), .QB (\$dummy [361]), 
        .D (L0_4_L1_2_Wij_nx222), .CLK (CLK)) ;
    dff L0_4_L1_2_Wij_reg_Dout_2 (.Q (WindowDout_4__2__2), .QB (\$dummy [362]), 
        .D (L0_4_L1_2_Wij_nx232), .CLK (CLK)) ;
    dff L0_4_L1_2_Wij_reg_Dout_3 (.Q (WindowDout_4__2__3), .QB (\$dummy [363]), 
        .D (L0_4_L1_2_Wij_nx242), .CLK (CLK)) ;
    dff L0_4_L1_2_Wij_reg_Dout_4 (.Q (WindowDout_4__2__4), .QB (\$dummy [364]), 
        .D (L0_4_L1_2_Wij_nx252), .CLK (CLK)) ;
    dff L0_4_L1_2_Wij_reg_Dout_5 (.Q (WindowDout_4__2__5), .QB (\$dummy [365]), 
        .D (L0_4_L1_2_Wij_nx262), .CLK (CLK)) ;
    dff L0_4_L1_2_Wij_reg_Dout_6 (.Q (WindowDout_4__2__6), .QB (\$dummy [366]), 
        .D (L0_4_L1_2_Wij_nx272), .CLK (CLK)) ;
    dff L0_4_L1_2_Wij_reg_Dout_7 (.Q (WindowDout_4__2__7), .QB (\$dummy [367]), 
        .D (L0_4_L1_2_Wij_nx282), .CLK (CLK)) ;
    buf02 L0_4_L1_2_Wij_ix330 (.Y (L0_4_L1_2_Wij_nx331), .A (WindowWR)) ;
    buf02 L0_4_L1_2_Wij_ix332 (.Y (L0_4_L1_2_Wij_nx333), .A (WindowWR)) ;
    dff L0_4_L1_3_Fij_reg_Dout_0 (.Q (FilterDout_4__3__0), .QB (\$dummy [368]), 
        .D (L0_4_L1_3_Fij_nx212), .CLK (CLK)) ;
    nor02_2x L0_4_L1_3_Fij_ix297 (.Y (L0_4_L1_3_Fij_nx296), .A0 (RST), .A1 (
             L0_4_L1_3_Fij_nx331)) ;
    dff L0_4_L1_3_Fij_reg_Dout_1 (.Q (FilterDout_4__3__1), .QB (\$dummy [369]), 
        .D (L0_4_L1_3_Fij_nx222), .CLK (CLK)) ;
    dff L0_4_L1_3_Fij_reg_Dout_2 (.Q (FilterDout_4__3__2), .QB (\$dummy [370]), 
        .D (L0_4_L1_3_Fij_nx232), .CLK (CLK)) ;
    dff L0_4_L1_3_Fij_reg_Dout_3 (.Q (FilterDout_4__3__3), .QB (\$dummy [371]), 
        .D (L0_4_L1_3_Fij_nx242), .CLK (CLK)) ;
    dff L0_4_L1_3_Fij_reg_Dout_4 (.Q (FilterDout_4__3__4), .QB (\$dummy [372]), 
        .D (L0_4_L1_3_Fij_nx252), .CLK (CLK)) ;
    dff L0_4_L1_3_Fij_reg_Dout_5 (.Q (FilterDout_4__3__5), .QB (\$dummy [373]), 
        .D (L0_4_L1_3_Fij_nx262), .CLK (CLK)) ;
    dff L0_4_L1_3_Fij_reg_Dout_6 (.Q (FilterDout_4__3__6), .QB (\$dummy [374]), 
        .D (L0_4_L1_3_Fij_nx272), .CLK (CLK)) ;
    dff L0_4_L1_3_Fij_reg_Dout_7 (.Q (FilterDout_4__3__7), .QB (\$dummy [375]), 
        .D (L0_4_L1_3_Fij_nx282), .CLK (CLK)) ;
    buf02 L0_4_L1_3_Fij_ix330 (.Y (L0_4_L1_3_Fij_nx331), .A (EN_dup_1411)) ;
    buf02 L0_4_L1_3_Fij_ix332 (.Y (L0_4_L1_3_Fij_nx333), .A (EN_dup_1411)) ;
    dff L0_4_L1_3_Wij_reg_Dout_0 (.Q (WindowDout_4__3__0), .QB (\$dummy [376]), 
        .D (L0_4_L1_3_Wij_nx212), .CLK (CLK)) ;
    nor02_2x L0_4_L1_3_Wij_ix297 (.Y (L0_4_L1_3_Wij_nx296), .A0 (RST), .A1 (
             L0_4_L1_3_Wij_nx331)) ;
    dff L0_4_L1_3_Wij_reg_Dout_1 (.Q (WindowDout_4__3__1), .QB (\$dummy [377]), 
        .D (L0_4_L1_3_Wij_nx222), .CLK (CLK)) ;
    dff L0_4_L1_3_Wij_reg_Dout_2 (.Q (WindowDout_4__3__2), .QB (\$dummy [378]), 
        .D (L0_4_L1_3_Wij_nx232), .CLK (CLK)) ;
    dff L0_4_L1_3_Wij_reg_Dout_3 (.Q (WindowDout_4__3__3), .QB (\$dummy [379]), 
        .D (L0_4_L1_3_Wij_nx242), .CLK (CLK)) ;
    dff L0_4_L1_3_Wij_reg_Dout_4 (.Q (WindowDout_4__3__4), .QB (\$dummy [380]), 
        .D (L0_4_L1_3_Wij_nx252), .CLK (CLK)) ;
    dff L0_4_L1_3_Wij_reg_Dout_5 (.Q (WindowDout_4__3__5), .QB (\$dummy [381]), 
        .D (L0_4_L1_3_Wij_nx262), .CLK (CLK)) ;
    dff L0_4_L1_3_Wij_reg_Dout_6 (.Q (WindowDout_4__3__6), .QB (\$dummy [382]), 
        .D (L0_4_L1_3_Wij_nx272), .CLK (CLK)) ;
    dff L0_4_L1_3_Wij_reg_Dout_7 (.Q (WindowDout_4__3__7), .QB (\$dummy [383]), 
        .D (L0_4_L1_3_Wij_nx282), .CLK (CLK)) ;
    buf02 L0_4_L1_3_Wij_ix330 (.Y (L0_4_L1_3_Wij_nx331), .A (EN_dup_1422)) ;
    buf02 L0_4_L1_3_Wij_ix332 (.Y (L0_4_L1_3_Wij_nx333), .A (EN_dup_1422)) ;
    dff L0_4_L1_4_Fij_reg_Dout_0 (.Q (FilterDout_4__4__0), .QB (\$dummy [384]), 
        .D (L0_4_L1_4_Fij_nx212), .CLK (CLK)) ;
    nor02_2x L0_4_L1_4_Fij_ix297 (.Y (L0_4_L1_4_Fij_nx296), .A0 (RST), .A1 (
             L0_4_L1_4_Fij_nx331)) ;
    dff L0_4_L1_4_Fij_reg_Dout_1 (.Q (FilterDout_4__4__1), .QB (\$dummy [385]), 
        .D (L0_4_L1_4_Fij_nx222), .CLK (CLK)) ;
    dff L0_4_L1_4_Fij_reg_Dout_2 (.Q (FilterDout_4__4__2), .QB (\$dummy [386]), 
        .D (L0_4_L1_4_Fij_nx232), .CLK (CLK)) ;
    dff L0_4_L1_4_Fij_reg_Dout_3 (.Q (FilterDout_4__4__3), .QB (\$dummy [387]), 
        .D (L0_4_L1_4_Fij_nx242), .CLK (CLK)) ;
    dff L0_4_L1_4_Fij_reg_Dout_4 (.Q (FilterDout_4__4__4), .QB (\$dummy [388]), 
        .D (L0_4_L1_4_Fij_nx252), .CLK (CLK)) ;
    dff L0_4_L1_4_Fij_reg_Dout_5 (.Q (FilterDout_4__4__5), .QB (\$dummy [389]), 
        .D (L0_4_L1_4_Fij_nx262), .CLK (CLK)) ;
    dff L0_4_L1_4_Fij_reg_Dout_6 (.Q (FilterDout_4__4__6), .QB (\$dummy [390]), 
        .D (L0_4_L1_4_Fij_nx272), .CLK (CLK)) ;
    dff L0_4_L1_4_Fij_reg_Dout_7 (.Q (FilterDout_4__4__7), .QB (\$dummy [391]), 
        .D (L0_4_L1_4_Fij_nx282), .CLK (CLK)) ;
    buf02 L0_4_L1_4_Fij_ix330 (.Y (L0_4_L1_4_Fij_nx331), .A (EN_dup_1411)) ;
    buf02 L0_4_L1_4_Fij_ix332 (.Y (L0_4_L1_4_Fij_nx333), .A (EN_dup_1411)) ;
    dff L0_4_L1_4_Wij_reg_Dout_0 (.Q (WindowDout_4__4__0), .QB (\$dummy [392]), 
        .D (L0_4_L1_4_Wij_nx212), .CLK (CLK)) ;
    nor02_2x L0_4_L1_4_Wij_ix297 (.Y (L0_4_L1_4_Wij_nx296), .A0 (RST), .A1 (
             L0_4_L1_4_Wij_nx331)) ;
    dff L0_4_L1_4_Wij_reg_Dout_1 (.Q (WindowDout_4__4__1), .QB (\$dummy [393]), 
        .D (L0_4_L1_4_Wij_nx222), .CLK (CLK)) ;
    dff L0_4_L1_4_Wij_reg_Dout_2 (.Q (WindowDout_4__4__2), .QB (\$dummy [394]), 
        .D (L0_4_L1_4_Wij_nx232), .CLK (CLK)) ;
    dff L0_4_L1_4_Wij_reg_Dout_3 (.Q (WindowDout_4__4__3), .QB (\$dummy [395]), 
        .D (L0_4_L1_4_Wij_nx242), .CLK (CLK)) ;
    dff L0_4_L1_4_Wij_reg_Dout_4 (.Q (WindowDout_4__4__4), .QB (\$dummy [396]), 
        .D (L0_4_L1_4_Wij_nx252), .CLK (CLK)) ;
    dff L0_4_L1_4_Wij_reg_Dout_5 (.Q (WindowDout_4__4__5), .QB (\$dummy [397]), 
        .D (L0_4_L1_4_Wij_nx262), .CLK (CLK)) ;
    dff L0_4_L1_4_Wij_reg_Dout_6 (.Q (WindowDout_4__4__6), .QB (\$dummy [398]), 
        .D (L0_4_L1_4_Wij_nx272), .CLK (CLK)) ;
    dff L0_4_L1_4_Wij_reg_Dout_7 (.Q (WindowDout_4__4__7), .QB (\$dummy [399]), 
        .D (L0_4_L1_4_Wij_nx282), .CLK (CLK)) ;
    buf02 L0_4_L1_4_Wij_ix330 (.Y (L0_4_L1_4_Wij_nx331), .A (EN_dup_1422)) ;
    buf02 L0_4_L1_4_Wij_ix332 (.Y (L0_4_L1_4_Wij_nx333), .A (EN_dup_1422)) ;
    oai32 L0_0_L1_0_Fij_ix213 (.Y (L0_0_L1_0_Fij_nx212), .A0 (nx1576), .A1 (RST)
          , .A2 (nx1578), .B0 (nx1580), .B1 (nx2756)) ;
    inv01 ix1575 (.Y (nx1576), .A (FilterDout_1__0__0)) ;
    inv02 ix1577 (.Y (nx1578), .A (L0_0_L1_0_Fij_nx331)) ;
    inv01 ix1579 (.Y (nx1580), .A (FilterDout_0__0__0)) ;
    oai32 L0_0_L1_0_Fij_ix223 (.Y (L0_0_L1_0_Fij_nx222), .A0 (nx1584), .A1 (RST)
          , .A2 (nx1578), .B0 (nx1586), .B1 (nx2756)) ;
    inv01 ix1583 (.Y (nx1584), .A (FilterDout_1__0__1)) ;
    inv01 ix1585 (.Y (nx1586), .A (FilterDout_0__0__1)) ;
    oai32 L0_0_L1_0_Fij_ix233 (.Y (L0_0_L1_0_Fij_nx232), .A0 (nx1588), .A1 (RST)
          , .A2 (nx1578), .B0 (nx1590), .B1 (nx2756)) ;
    inv01 ix1587 (.Y (nx1588), .A (FilterDout_1__0__2)) ;
    inv01 ix1589 (.Y (nx1590), .A (FilterDout_0__0__2)) ;
    oai32 L0_0_L1_0_Fij_ix243 (.Y (L0_0_L1_0_Fij_nx242), .A0 (nx1592), .A1 (RST)
          , .A2 (nx1578), .B0 (nx1594), .B1 (nx2756)) ;
    inv01 ix1591 (.Y (nx1592), .A (FilterDout_1__0__3)) ;
    inv01 ix1593 (.Y (nx1594), .A (FilterDout_0__0__3)) ;
    oai32 L0_0_L1_0_Fij_ix253 (.Y (L0_0_L1_0_Fij_nx252), .A0 (nx1596), .A1 (RST)
          , .A2 (nx1578), .B0 (nx1598), .B1 (nx2756)) ;
    inv01 ix1595 (.Y (nx1596), .A (FilterDout_1__0__4)) ;
    inv01 ix1597 (.Y (nx1598), .A (FilterDout_0__0__4)) ;
    oai32 L0_0_L1_0_Fij_ix263 (.Y (L0_0_L1_0_Fij_nx262), .A0 (nx1600), .A1 (RST)
          , .A2 (nx1578), .B0 (nx1602), .B1 (nx2756)) ;
    inv01 ix1599 (.Y (nx1600), .A (FilterDout_1__0__5)) ;
    inv01 ix1601 (.Y (nx1602), .A (FilterDout_0__0__5)) ;
    oai32 L0_0_L1_0_Fij_ix273 (.Y (L0_0_L1_0_Fij_nx272), .A0 (nx1604), .A1 (RST)
          , .A2 (nx1606), .B0 (nx1608), .B1 (nx2756)) ;
    inv01 ix1603 (.Y (nx1604), .A (FilterDout_1__0__6)) ;
    inv01 ix1605 (.Y (nx1606), .A (L0_0_L1_0_Fij_nx333)) ;
    inv01 ix1607 (.Y (nx1608), .A (FilterDout_0__0__6)) ;
    oai32 L0_0_L1_0_Fij_ix283 (.Y (L0_0_L1_0_Fij_nx282), .A0 (nx1610), .A1 (RST)
          , .A2 (nx1606), .B0 (nx1612), .B1 (nx2758)) ;
    inv01 ix1609 (.Y (nx1610), .A (FilterDout_1__0__7)) ;
    inv01 ix1611 (.Y (nx1612), .A (FilterDout_0__0__7)) ;
    oai32 L0_0_L1_0_Wij_ix213 (.Y (L0_0_L1_0_Wij_nx212), .A0 (nx1614), .A1 (RST)
          , .A2 (nx1616), .B0 (nx1618), .B1 (nx2760)) ;
    inv01 ix1613 (.Y (nx1614), .A (WindowDout_1__0__0)) ;
    inv02 ix1615 (.Y (nx1616), .A (L0_0_L1_0_Wij_nx331)) ;
    inv01 ix1617 (.Y (nx1618), .A (WindowDout_0__0__0)) ;
    oai32 L0_0_L1_0_Wij_ix223 (.Y (L0_0_L1_0_Wij_nx222), .A0 (nx1622), .A1 (RST)
          , .A2 (nx1616), .B0 (nx1624), .B1 (nx2760)) ;
    inv01 ix1621 (.Y (nx1622), .A (WindowDout_1__0__1)) ;
    inv01 ix1623 (.Y (nx1624), .A (WindowDout_0__0__1)) ;
    oai32 L0_0_L1_0_Wij_ix233 (.Y (L0_0_L1_0_Wij_nx232), .A0 (nx1626), .A1 (RST)
          , .A2 (nx1616), .B0 (nx1628), .B1 (nx2760)) ;
    inv01 ix1625 (.Y (nx1626), .A (WindowDout_1__0__2)) ;
    inv01 ix1627 (.Y (nx1628), .A (WindowDout_0__0__2)) ;
    oai32 L0_0_L1_0_Wij_ix243 (.Y (L0_0_L1_0_Wij_nx242), .A0 (nx1630), .A1 (RST)
          , .A2 (nx1616), .B0 (nx1632), .B1 (nx2760)) ;
    inv01 ix1629 (.Y (nx1630), .A (WindowDout_1__0__3)) ;
    inv01 ix1631 (.Y (nx1632), .A (WindowDout_0__0__3)) ;
    oai32 L0_0_L1_0_Wij_ix253 (.Y (L0_0_L1_0_Wij_nx252), .A0 (nx1634), .A1 (RST)
          , .A2 (nx1616), .B0 (nx1636), .B1 (nx2760)) ;
    inv01 ix1633 (.Y (nx1634), .A (WindowDout_1__0__4)) ;
    inv01 ix1635 (.Y (nx1636), .A (WindowDout_0__0__4)) ;
    oai32 L0_0_L1_0_Wij_ix263 (.Y (L0_0_L1_0_Wij_nx262), .A0 (nx1638), .A1 (RST)
          , .A2 (nx1616), .B0 (nx1640), .B1 (nx2760)) ;
    inv01 ix1637 (.Y (nx1638), .A (WindowDout_1__0__5)) ;
    inv01 ix1639 (.Y (nx1640), .A (WindowDout_0__0__5)) ;
    oai32 L0_0_L1_0_Wij_ix273 (.Y (L0_0_L1_0_Wij_nx272), .A0 (nx1642), .A1 (RST)
          , .A2 (nx1644), .B0 (nx1646), .B1 (nx2760)) ;
    inv01 ix1641 (.Y (nx1642), .A (WindowDout_1__0__6)) ;
    inv01 ix1643 (.Y (nx1644), .A (L0_0_L1_0_Wij_nx333)) ;
    inv01 ix1645 (.Y (nx1646), .A (WindowDout_0__0__6)) ;
    oai32 L0_0_L1_0_Wij_ix283 (.Y (L0_0_L1_0_Wij_nx282), .A0 (nx1648), .A1 (RST)
          , .A2 (nx1644), .B0 (nx1650), .B1 (nx2762)) ;
    inv01 ix1647 (.Y (nx1648), .A (WindowDout_1__0__7)) ;
    inv01 ix1649 (.Y (nx1650), .A (WindowDout_0__0__7)) ;
    oai32 L0_0_L1_1_Fij_ix213 (.Y (L0_0_L1_1_Fij_nx212), .A0 (nx1652), .A1 (RST)
          , .A2 (nx1654), .B0 (nx1656), .B1 (nx2764)) ;
    inv01 ix1651 (.Y (nx1652), .A (FilterDout_1__1__0)) ;
    inv02 ix1653 (.Y (nx1654), .A (L0_0_L1_1_Fij_nx331)) ;
    inv01 ix1655 (.Y (nx1656), .A (FilterDout_0__1__0)) ;
    oai32 L0_0_L1_1_Fij_ix223 (.Y (L0_0_L1_1_Fij_nx222), .A0 (nx1660), .A1 (RST)
          , .A2 (nx1654), .B0 (nx1662), .B1 (nx2764)) ;
    inv01 ix1659 (.Y (nx1660), .A (FilterDout_1__1__1)) ;
    inv01 ix1661 (.Y (nx1662), .A (FilterDout_0__1__1)) ;
    oai32 L0_0_L1_1_Fij_ix233 (.Y (L0_0_L1_1_Fij_nx232), .A0 (nx1664), .A1 (RST)
          , .A2 (nx1654), .B0 (nx1666), .B1 (nx2764)) ;
    inv01 ix1663 (.Y (nx1664), .A (FilterDout_1__1__2)) ;
    inv01 ix1665 (.Y (nx1666), .A (FilterDout_0__1__2)) ;
    oai32 L0_0_L1_1_Fij_ix243 (.Y (L0_0_L1_1_Fij_nx242), .A0 (nx1668), .A1 (RST)
          , .A2 (nx1654), .B0 (nx1670), .B1 (nx2764)) ;
    inv01 ix1667 (.Y (nx1668), .A (FilterDout_1__1__3)) ;
    inv01 ix1669 (.Y (nx1670), .A (FilterDout_0__1__3)) ;
    oai32 L0_0_L1_1_Fij_ix253 (.Y (L0_0_L1_1_Fij_nx252), .A0 (nx1672), .A1 (RST)
          , .A2 (nx1654), .B0 (nx1674), .B1 (nx2764)) ;
    inv01 ix1671 (.Y (nx1672), .A (FilterDout_1__1__4)) ;
    inv01 ix1673 (.Y (nx1674), .A (FilterDout_0__1__4)) ;
    oai32 L0_0_L1_1_Fij_ix263 (.Y (L0_0_L1_1_Fij_nx262), .A0 (nx1676), .A1 (RST)
          , .A2 (nx1654), .B0 (nx1678), .B1 (nx2764)) ;
    inv01 ix1675 (.Y (nx1676), .A (FilterDout_1__1__5)) ;
    inv01 ix1677 (.Y (nx1678), .A (FilterDout_0__1__5)) ;
    oai32 L0_0_L1_1_Fij_ix273 (.Y (L0_0_L1_1_Fij_nx272), .A0 (nx1680), .A1 (RST)
          , .A2 (nx1682), .B0 (nx1684), .B1 (nx2764)) ;
    inv01 ix1679 (.Y (nx1680), .A (FilterDout_1__1__6)) ;
    inv01 ix1681 (.Y (nx1682), .A (L0_0_L1_1_Fij_nx333)) ;
    inv01 ix1683 (.Y (nx1684), .A (FilterDout_0__1__6)) ;
    oai32 L0_0_L1_1_Fij_ix283 (.Y (L0_0_L1_1_Fij_nx282), .A0 (nx1686), .A1 (RST)
          , .A2 (nx1682), .B0 (nx1688), .B1 (nx2766)) ;
    inv01 ix1685 (.Y (nx1686), .A (FilterDout_1__1__7)) ;
    inv01 ix1687 (.Y (nx1688), .A (FilterDout_0__1__7)) ;
    oai32 L0_0_L1_1_Wij_ix213 (.Y (L0_0_L1_1_Wij_nx212), .A0 (nx1690), .A1 (RST)
          , .A2 (nx1692), .B0 (nx1694), .B1 (nx2768)) ;
    inv01 ix1689 (.Y (nx1690), .A (WindowDout_1__1__0)) ;
    inv02 ix1691 (.Y (nx1692), .A (L0_0_L1_1_Wij_nx331)) ;
    inv01 ix1693 (.Y (nx1694), .A (WindowDout_0__1__0)) ;
    oai32 L0_0_L1_1_Wij_ix223 (.Y (L0_0_L1_1_Wij_nx222), .A0 (nx1698), .A1 (RST)
          , .A2 (nx1692), .B0 (nx1700), .B1 (nx2768)) ;
    inv01 ix1697 (.Y (nx1698), .A (WindowDout_1__1__1)) ;
    inv01 ix1699 (.Y (nx1700), .A (WindowDout_0__1__1)) ;
    oai32 L0_0_L1_1_Wij_ix233 (.Y (L0_0_L1_1_Wij_nx232), .A0 (nx1702), .A1 (RST)
          , .A2 (nx1692), .B0 (nx1704), .B1 (nx2768)) ;
    inv01 ix1701 (.Y (nx1702), .A (WindowDout_1__1__2)) ;
    inv01 ix1703 (.Y (nx1704), .A (WindowDout_0__1__2)) ;
    oai32 L0_0_L1_1_Wij_ix243 (.Y (L0_0_L1_1_Wij_nx242), .A0 (nx1706), .A1 (RST)
          , .A2 (nx1692), .B0 (nx1708), .B1 (nx2768)) ;
    inv01 ix1705 (.Y (nx1706), .A (WindowDout_1__1__3)) ;
    inv01 ix1707 (.Y (nx1708), .A (WindowDout_0__1__3)) ;
    oai32 L0_0_L1_1_Wij_ix253 (.Y (L0_0_L1_1_Wij_nx252), .A0 (nx1710), .A1 (RST)
          , .A2 (nx1692), .B0 (nx1712), .B1 (nx2768)) ;
    inv01 ix1709 (.Y (nx1710), .A (WindowDout_1__1__4)) ;
    inv01 ix1711 (.Y (nx1712), .A (WindowDout_0__1__4)) ;
    oai32 L0_0_L1_1_Wij_ix263 (.Y (L0_0_L1_1_Wij_nx262), .A0 (nx1714), .A1 (RST)
          , .A2 (nx1692), .B0 (nx1716), .B1 (nx2768)) ;
    inv01 ix1713 (.Y (nx1714), .A (WindowDout_1__1__5)) ;
    inv01 ix1715 (.Y (nx1716), .A (WindowDout_0__1__5)) ;
    oai32 L0_0_L1_1_Wij_ix273 (.Y (L0_0_L1_1_Wij_nx272), .A0 (nx1718), .A1 (RST)
          , .A2 (nx1720), .B0 (nx1722), .B1 (nx2768)) ;
    inv01 ix1717 (.Y (nx1718), .A (WindowDout_1__1__6)) ;
    inv01 ix1719 (.Y (nx1720), .A (L0_0_L1_1_Wij_nx333)) ;
    inv01 ix1721 (.Y (nx1722), .A (WindowDout_0__1__6)) ;
    oai32 L0_0_L1_1_Wij_ix283 (.Y (L0_0_L1_1_Wij_nx282), .A0 (nx1724), .A1 (RST)
          , .A2 (nx1720), .B0 (nx1726), .B1 (nx2770)) ;
    inv01 ix1723 (.Y (nx1724), .A (WindowDout_1__1__7)) ;
    inv01 ix1725 (.Y (nx1726), .A (WindowDout_0__1__7)) ;
    oai32 L0_0_L1_2_Fij_ix213 (.Y (L0_0_L1_2_Fij_nx212), .A0 (nx1728), .A1 (RST)
          , .A2 (nx1730), .B0 (nx1732), .B1 (nx2772)) ;
    inv01 ix1727 (.Y (nx1728), .A (FilterDout_1__2__0)) ;
    inv02 ix1729 (.Y (nx1730), .A (L0_0_L1_2_Fij_nx331)) ;
    inv01 ix1731 (.Y (nx1732), .A (FilterDout_0__2__0)) ;
    oai32 L0_0_L1_2_Fij_ix223 (.Y (L0_0_L1_2_Fij_nx222), .A0 (nx1736), .A1 (RST)
          , .A2 (nx1730), .B0 (nx1738), .B1 (nx2772)) ;
    inv01 ix1735 (.Y (nx1736), .A (FilterDout_1__2__1)) ;
    inv01 ix1737 (.Y (nx1738), .A (FilterDout_0__2__1)) ;
    oai32 L0_0_L1_2_Fij_ix233 (.Y (L0_0_L1_2_Fij_nx232), .A0 (nx1740), .A1 (RST)
          , .A2 (nx1730), .B0 (nx1742), .B1 (nx2772)) ;
    inv01 ix1739 (.Y (nx1740), .A (FilterDout_1__2__2)) ;
    inv01 ix1741 (.Y (nx1742), .A (FilterDout_0__2__2)) ;
    oai32 L0_0_L1_2_Fij_ix243 (.Y (L0_0_L1_2_Fij_nx242), .A0 (nx1744), .A1 (RST)
          , .A2 (nx1730), .B0 (nx1746), .B1 (nx2772)) ;
    inv01 ix1743 (.Y (nx1744), .A (FilterDout_1__2__3)) ;
    inv01 ix1745 (.Y (nx1746), .A (FilterDout_0__2__3)) ;
    oai32 L0_0_L1_2_Fij_ix253 (.Y (L0_0_L1_2_Fij_nx252), .A0 (nx1748), .A1 (RST)
          , .A2 (nx1730), .B0 (nx1750), .B1 (nx2772)) ;
    inv01 ix1747 (.Y (nx1748), .A (FilterDout_1__2__4)) ;
    inv01 ix1749 (.Y (nx1750), .A (FilterDout_0__2__4)) ;
    oai32 L0_0_L1_2_Fij_ix263 (.Y (L0_0_L1_2_Fij_nx262), .A0 (nx1752), .A1 (RST)
          , .A2 (nx1730), .B0 (nx1754), .B1 (nx2772)) ;
    inv01 ix1751 (.Y (nx1752), .A (FilterDout_1__2__5)) ;
    inv01 ix1753 (.Y (nx1754), .A (FilterDout_0__2__5)) ;
    oai32 L0_0_L1_2_Fij_ix273 (.Y (L0_0_L1_2_Fij_nx272), .A0 (nx1756), .A1 (RST)
          , .A2 (nx1758), .B0 (nx1760), .B1 (nx2772)) ;
    inv01 ix1755 (.Y (nx1756), .A (FilterDout_1__2__6)) ;
    inv01 ix1757 (.Y (nx1758), .A (L0_0_L1_2_Fij_nx333)) ;
    inv01 ix1759 (.Y (nx1760), .A (FilterDout_0__2__6)) ;
    oai32 L0_0_L1_2_Fij_ix283 (.Y (L0_0_L1_2_Fij_nx282), .A0 (nx1762), .A1 (RST)
          , .A2 (nx1758), .B0 (nx1764), .B1 (nx2774)) ;
    inv01 ix1761 (.Y (nx1762), .A (FilterDout_1__2__7)) ;
    inv01 ix1763 (.Y (nx1764), .A (FilterDout_0__2__7)) ;
    oai32 L0_0_L1_2_Wij_ix213 (.Y (L0_0_L1_2_Wij_nx212), .A0 (nx1766), .A1 (RST)
          , .A2 (nx1768), .B0 (nx1770), .B1 (nx2776)) ;
    inv01 ix1765 (.Y (nx1766), .A (WindowDout_1__2__0)) ;
    inv02 ix1767 (.Y (nx1768), .A (L0_0_L1_2_Wij_nx331)) ;
    inv01 ix1769 (.Y (nx1770), .A (WindowDout_0__2__0)) ;
    oai32 L0_0_L1_2_Wij_ix223 (.Y (L0_0_L1_2_Wij_nx222), .A0 (nx1774), .A1 (RST)
          , .A2 (nx1768), .B0 (nx1776), .B1 (nx2776)) ;
    inv01 ix1773 (.Y (nx1774), .A (WindowDout_1__2__1)) ;
    inv01 ix1775 (.Y (nx1776), .A (WindowDout_0__2__1)) ;
    oai32 L0_0_L1_2_Wij_ix233 (.Y (L0_0_L1_2_Wij_nx232), .A0 (nx1778), .A1 (RST)
          , .A2 (nx1768), .B0 (nx1780), .B1 (nx2776)) ;
    inv01 ix1777 (.Y (nx1778), .A (WindowDout_1__2__2)) ;
    inv01 ix1779 (.Y (nx1780), .A (WindowDout_0__2__2)) ;
    oai32 L0_0_L1_2_Wij_ix243 (.Y (L0_0_L1_2_Wij_nx242), .A0 (nx1782), .A1 (RST)
          , .A2 (nx1768), .B0 (nx1784), .B1 (nx2776)) ;
    inv01 ix1781 (.Y (nx1782), .A (WindowDout_1__2__3)) ;
    inv01 ix1783 (.Y (nx1784), .A (WindowDout_0__2__3)) ;
    oai32 L0_0_L1_2_Wij_ix253 (.Y (L0_0_L1_2_Wij_nx252), .A0 (nx1786), .A1 (RST)
          , .A2 (nx1768), .B0 (nx1788), .B1 (nx2776)) ;
    inv01 ix1785 (.Y (nx1786), .A (WindowDout_1__2__4)) ;
    inv01 ix1787 (.Y (nx1788), .A (WindowDout_0__2__4)) ;
    oai32 L0_0_L1_2_Wij_ix263 (.Y (L0_0_L1_2_Wij_nx262), .A0 (nx1790), .A1 (RST)
          , .A2 (nx1768), .B0 (nx1792), .B1 (nx2776)) ;
    inv01 ix1789 (.Y (nx1790), .A (WindowDout_1__2__5)) ;
    inv01 ix1791 (.Y (nx1792), .A (WindowDout_0__2__5)) ;
    oai32 L0_0_L1_2_Wij_ix273 (.Y (L0_0_L1_2_Wij_nx272), .A0 (nx1794), .A1 (RST)
          , .A2 (nx1796), .B0 (nx1798), .B1 (nx2776)) ;
    inv01 ix1793 (.Y (nx1794), .A (WindowDout_1__2__6)) ;
    inv01 ix1795 (.Y (nx1796), .A (L0_0_L1_2_Wij_nx333)) ;
    inv01 ix1797 (.Y (nx1798), .A (WindowDout_0__2__6)) ;
    oai32 L0_0_L1_2_Wij_ix283 (.Y (L0_0_L1_2_Wij_nx282), .A0 (nx1800), .A1 (RST)
          , .A2 (nx1796), .B0 (nx1802), .B1 (nx2778)) ;
    inv01 ix1799 (.Y (nx1800), .A (WindowDout_1__2__7)) ;
    inv01 ix1801 (.Y (nx1802), .A (WindowDout_0__2__7)) ;
    oai32 L0_0_L1_3_Fij_ix213 (.Y (L0_0_L1_3_Fij_nx212), .A0 (nx1804), .A1 (RST)
          , .A2 (nx1806), .B0 (nx1808), .B1 (nx2780)) ;
    inv01 ix1803 (.Y (nx1804), .A (FilterDout_1__3__0)) ;
    inv02 ix1805 (.Y (nx1806), .A (L0_0_L1_3_Fij_nx331)) ;
    inv01 ix1807 (.Y (nx1808), .A (FilterDout_0__3__0)) ;
    oai32 L0_0_L1_3_Fij_ix223 (.Y (L0_0_L1_3_Fij_nx222), .A0 (nx1812), .A1 (RST)
          , .A2 (nx1806), .B0 (nx1814), .B1 (nx2780)) ;
    inv01 ix1811 (.Y (nx1812), .A (FilterDout_1__3__1)) ;
    inv01 ix1813 (.Y (nx1814), .A (FilterDout_0__3__1)) ;
    oai32 L0_0_L1_3_Fij_ix233 (.Y (L0_0_L1_3_Fij_nx232), .A0 (nx1816), .A1 (RST)
          , .A2 (nx1806), .B0 (nx1818), .B1 (nx2780)) ;
    inv01 ix1815 (.Y (nx1816), .A (FilterDout_1__3__2)) ;
    inv01 ix1817 (.Y (nx1818), .A (FilterDout_0__3__2)) ;
    oai32 L0_0_L1_3_Fij_ix243 (.Y (L0_0_L1_3_Fij_nx242), .A0 (nx1820), .A1 (RST)
          , .A2 (nx1806), .B0 (nx1822), .B1 (nx2780)) ;
    inv01 ix1819 (.Y (nx1820), .A (FilterDout_1__3__3)) ;
    inv01 ix1821 (.Y (nx1822), .A (FilterDout_0__3__3)) ;
    oai32 L0_0_L1_3_Fij_ix253 (.Y (L0_0_L1_3_Fij_nx252), .A0 (nx1824), .A1 (RST)
          , .A2 (nx1806), .B0 (nx1826), .B1 (nx2780)) ;
    inv01 ix1823 (.Y (nx1824), .A (FilterDout_1__3__4)) ;
    inv01 ix1825 (.Y (nx1826), .A (FilterDout_0__3__4)) ;
    oai32 L0_0_L1_3_Fij_ix263 (.Y (L0_0_L1_3_Fij_nx262), .A0 (nx1828), .A1 (RST)
          , .A2 (nx1806), .B0 (nx1830), .B1 (nx2780)) ;
    inv01 ix1827 (.Y (nx1828), .A (FilterDout_1__3__5)) ;
    inv01 ix1829 (.Y (nx1830), .A (FilterDout_0__3__5)) ;
    oai32 L0_0_L1_3_Fij_ix273 (.Y (L0_0_L1_3_Fij_nx272), .A0 (nx1832), .A1 (RST)
          , .A2 (nx1834), .B0 (nx1836), .B1 (nx2780)) ;
    inv01 ix1831 (.Y (nx1832), .A (FilterDout_1__3__6)) ;
    inv01 ix1833 (.Y (nx1834), .A (L0_0_L1_3_Fij_nx333)) ;
    inv01 ix1835 (.Y (nx1836), .A (FilterDout_0__3__6)) ;
    oai32 L0_0_L1_3_Fij_ix283 (.Y (L0_0_L1_3_Fij_nx282), .A0 (nx1838), .A1 (RST)
          , .A2 (nx1834), .B0 (nx1840), .B1 (nx2782)) ;
    inv01 ix1837 (.Y (nx1838), .A (FilterDout_1__3__7)) ;
    inv01 ix1839 (.Y (nx1840), .A (FilterDout_0__3__7)) ;
    oai32 L0_0_L1_3_Wij_ix213 (.Y (L0_0_L1_3_Wij_nx212), .A0 (nx1842), .A1 (RST)
          , .A2 (nx1844), .B0 (nx1846), .B1 (nx2784)) ;
    inv01 ix1841 (.Y (nx1842), .A (WindowDout_1__3__0)) ;
    inv02 ix1843 (.Y (nx1844), .A (L0_0_L1_3_Wij_nx331)) ;
    inv01 ix1845 (.Y (nx1846), .A (WindowDout_0__3__0)) ;
    oai32 L0_0_L1_3_Wij_ix223 (.Y (L0_0_L1_3_Wij_nx222), .A0 (nx1850), .A1 (RST)
          , .A2 (nx1844), .B0 (nx1852), .B1 (nx2784)) ;
    inv01 ix1849 (.Y (nx1850), .A (WindowDout_1__3__1)) ;
    inv01 ix1851 (.Y (nx1852), .A (WindowDout_0__3__1)) ;
    oai32 L0_0_L1_3_Wij_ix233 (.Y (L0_0_L1_3_Wij_nx232), .A0 (nx1854), .A1 (RST)
          , .A2 (nx1844), .B0 (nx1856), .B1 (nx2784)) ;
    inv01 ix1853 (.Y (nx1854), .A (WindowDout_1__3__2)) ;
    inv01 ix1855 (.Y (nx1856), .A (WindowDout_0__3__2)) ;
    oai32 L0_0_L1_3_Wij_ix243 (.Y (L0_0_L1_3_Wij_nx242), .A0 (nx1858), .A1 (RST)
          , .A2 (nx1844), .B0 (nx1860), .B1 (nx2784)) ;
    inv01 ix1857 (.Y (nx1858), .A (WindowDout_1__3__3)) ;
    inv01 ix1859 (.Y (nx1860), .A (WindowDout_0__3__3)) ;
    oai32 L0_0_L1_3_Wij_ix253 (.Y (L0_0_L1_3_Wij_nx252), .A0 (nx1862), .A1 (RST)
          , .A2 (nx1844), .B0 (nx1864), .B1 (nx2784)) ;
    inv01 ix1861 (.Y (nx1862), .A (WindowDout_1__3__4)) ;
    inv01 ix1863 (.Y (nx1864), .A (WindowDout_0__3__4)) ;
    oai32 L0_0_L1_3_Wij_ix263 (.Y (L0_0_L1_3_Wij_nx262), .A0 (nx1866), .A1 (RST)
          , .A2 (nx1844), .B0 (nx1868), .B1 (nx2784)) ;
    inv01 ix1865 (.Y (nx1866), .A (WindowDout_1__3__5)) ;
    inv01 ix1867 (.Y (nx1868), .A (WindowDout_0__3__5)) ;
    oai32 L0_0_L1_3_Wij_ix273 (.Y (L0_0_L1_3_Wij_nx272), .A0 (nx1870), .A1 (RST)
          , .A2 (nx1872), .B0 (nx1874), .B1 (nx2784)) ;
    inv01 ix1869 (.Y (nx1870), .A (WindowDout_1__3__6)) ;
    inv01 ix1871 (.Y (nx1872), .A (L0_0_L1_3_Wij_nx333)) ;
    inv01 ix1873 (.Y (nx1874), .A (WindowDout_0__3__6)) ;
    oai32 L0_0_L1_3_Wij_ix283 (.Y (L0_0_L1_3_Wij_nx282), .A0 (nx1876), .A1 (RST)
          , .A2 (nx1872), .B0 (nx1878), .B1 (nx2786)) ;
    inv01 ix1875 (.Y (nx1876), .A (WindowDout_1__3__7)) ;
    inv01 ix1877 (.Y (nx1878), .A (WindowDout_0__3__7)) ;
    oai32 L0_0_L1_4_Fij_ix213 (.Y (L0_0_L1_4_Fij_nx212), .A0 (nx1880), .A1 (RST)
          , .A2 (nx1882), .B0 (nx1884), .B1 (nx2788)) ;
    inv01 ix1879 (.Y (nx1880), .A (FilterDout_1__4__0)) ;
    inv02 ix1881 (.Y (nx1882), .A (L0_0_L1_4_Fij_nx331)) ;
    inv01 ix1883 (.Y (nx1884), .A (FilterDout_0__4__0)) ;
    oai32 L0_0_L1_4_Fij_ix223 (.Y (L0_0_L1_4_Fij_nx222), .A0 (nx1888), .A1 (RST)
          , .A2 (nx1882), .B0 (nx1890), .B1 (nx2788)) ;
    inv01 ix1887 (.Y (nx1888), .A (FilterDout_1__4__1)) ;
    inv01 ix1889 (.Y (nx1890), .A (FilterDout_0__4__1)) ;
    oai32 L0_0_L1_4_Fij_ix233 (.Y (L0_0_L1_4_Fij_nx232), .A0 (nx1892), .A1 (RST)
          , .A2 (nx1882), .B0 (nx1894), .B1 (nx2788)) ;
    inv01 ix1891 (.Y (nx1892), .A (FilterDout_1__4__2)) ;
    inv01 ix1893 (.Y (nx1894), .A (FilterDout_0__4__2)) ;
    oai32 L0_0_L1_4_Fij_ix243 (.Y (L0_0_L1_4_Fij_nx242), .A0 (nx1896), .A1 (RST)
          , .A2 (nx1882), .B0 (nx1898), .B1 (nx2788)) ;
    inv01 ix1895 (.Y (nx1896), .A (FilterDout_1__4__3)) ;
    inv01 ix1897 (.Y (nx1898), .A (FilterDout_0__4__3)) ;
    oai32 L0_0_L1_4_Fij_ix253 (.Y (L0_0_L1_4_Fij_nx252), .A0 (nx1900), .A1 (RST)
          , .A2 (nx1882), .B0 (nx1902), .B1 (nx2788)) ;
    inv01 ix1899 (.Y (nx1900), .A (FilterDout_1__4__4)) ;
    inv01 ix1901 (.Y (nx1902), .A (FilterDout_0__4__4)) ;
    oai32 L0_0_L1_4_Fij_ix263 (.Y (L0_0_L1_4_Fij_nx262), .A0 (nx1904), .A1 (RST)
          , .A2 (nx1882), .B0 (nx1906), .B1 (nx2788)) ;
    inv01 ix1903 (.Y (nx1904), .A (FilterDout_1__4__5)) ;
    inv01 ix1905 (.Y (nx1906), .A (FilterDout_0__4__5)) ;
    oai32 L0_0_L1_4_Fij_ix273 (.Y (L0_0_L1_4_Fij_nx272), .A0 (nx1908), .A1 (RST)
          , .A2 (nx1910), .B0 (nx1912), .B1 (nx2788)) ;
    inv01 ix1907 (.Y (nx1908), .A (FilterDout_1__4__6)) ;
    inv01 ix1909 (.Y (nx1910), .A (L0_0_L1_4_Fij_nx333)) ;
    inv01 ix1911 (.Y (nx1912), .A (FilterDout_0__4__6)) ;
    oai32 L0_0_L1_4_Fij_ix283 (.Y (L0_0_L1_4_Fij_nx282), .A0 (nx1914), .A1 (RST)
          , .A2 (nx1910), .B0 (nx1916), .B1 (nx2790)) ;
    inv01 ix1913 (.Y (nx1914), .A (FilterDout_1__4__7)) ;
    inv01 ix1915 (.Y (nx1916), .A (FilterDout_0__4__7)) ;
    oai32 L0_0_L1_4_Wij_ix213 (.Y (L0_0_L1_4_Wij_nx212), .A0 (nx1918), .A1 (RST)
          , .A2 (nx1920), .B0 (nx1922), .B1 (nx2792)) ;
    inv01 ix1917 (.Y (nx1918), .A (WindowDout_1__4__0)) ;
    inv02 ix1919 (.Y (nx1920), .A (L0_0_L1_4_Wij_nx331)) ;
    inv01 ix1921 (.Y (nx1922), .A (WindowDout_0__4__0)) ;
    oai32 L0_0_L1_4_Wij_ix223 (.Y (L0_0_L1_4_Wij_nx222), .A0 (nx1926), .A1 (RST)
          , .A2 (nx1920), .B0 (nx1928), .B1 (nx2792)) ;
    inv01 ix1925 (.Y (nx1926), .A (WindowDout_1__4__1)) ;
    inv01 ix1927 (.Y (nx1928), .A (WindowDout_0__4__1)) ;
    oai32 L0_0_L1_4_Wij_ix233 (.Y (L0_0_L1_4_Wij_nx232), .A0 (nx1930), .A1 (RST)
          , .A2 (nx1920), .B0 (nx1932), .B1 (nx2792)) ;
    inv01 ix1929 (.Y (nx1930), .A (WindowDout_1__4__2)) ;
    inv01 ix1931 (.Y (nx1932), .A (WindowDout_0__4__2)) ;
    oai32 L0_0_L1_4_Wij_ix243 (.Y (L0_0_L1_4_Wij_nx242), .A0 (nx1934), .A1 (RST)
          , .A2 (nx1920), .B0 (nx1936), .B1 (nx2792)) ;
    inv01 ix1933 (.Y (nx1934), .A (WindowDout_1__4__3)) ;
    inv01 ix1935 (.Y (nx1936), .A (WindowDout_0__4__3)) ;
    oai32 L0_0_L1_4_Wij_ix253 (.Y (L0_0_L1_4_Wij_nx252), .A0 (nx1938), .A1 (RST)
          , .A2 (nx1920), .B0 (nx1940), .B1 (nx2792)) ;
    inv01 ix1937 (.Y (nx1938), .A (WindowDout_1__4__4)) ;
    inv01 ix1939 (.Y (nx1940), .A (WindowDout_0__4__4)) ;
    oai32 L0_0_L1_4_Wij_ix263 (.Y (L0_0_L1_4_Wij_nx262), .A0 (nx1942), .A1 (RST)
          , .A2 (nx1920), .B0 (nx1944), .B1 (nx2792)) ;
    inv01 ix1941 (.Y (nx1942), .A (WindowDout_1__4__5)) ;
    inv01 ix1943 (.Y (nx1944), .A (WindowDout_0__4__5)) ;
    oai32 L0_0_L1_4_Wij_ix273 (.Y (L0_0_L1_4_Wij_nx272), .A0 (nx1946), .A1 (RST)
          , .A2 (nx1948), .B0 (nx1950), .B1 (nx2792)) ;
    inv01 ix1945 (.Y (nx1946), .A (WindowDout_1__4__6)) ;
    inv01 ix1947 (.Y (nx1948), .A (L0_0_L1_4_Wij_nx333)) ;
    inv01 ix1949 (.Y (nx1950), .A (WindowDout_0__4__6)) ;
    oai32 L0_0_L1_4_Wij_ix283 (.Y (L0_0_L1_4_Wij_nx282), .A0 (nx1952), .A1 (RST)
          , .A2 (nx1948), .B0 (nx1954), .B1 (nx2794)) ;
    inv01 ix1951 (.Y (nx1952), .A (WindowDout_1__4__7)) ;
    inv01 ix1953 (.Y (nx1954), .A (WindowDout_0__4__7)) ;
    oai32 L0_1_L1_0_Fij_ix213 (.Y (L0_1_L1_0_Fij_nx212), .A0 (nx1956), .A1 (RST)
          , .A2 (nx1958), .B0 (nx1576), .B1 (nx2796)) ;
    inv01 ix1955 (.Y (nx1956), .A (FilterDout_2__0__0)) ;
    inv02 ix1957 (.Y (nx1958), .A (L0_1_L1_0_Fij_nx331)) ;
    oai32 L0_1_L1_0_Fij_ix223 (.Y (L0_1_L1_0_Fij_nx222), .A0 (nx1962), .A1 (RST)
          , .A2 (nx1958), .B0 (nx1584), .B1 (nx2796)) ;
    inv01 ix1961 (.Y (nx1962), .A (FilterDout_2__0__1)) ;
    oai32 L0_1_L1_0_Fij_ix233 (.Y (L0_1_L1_0_Fij_nx232), .A0 (nx1964), .A1 (RST)
          , .A2 (nx1958), .B0 (nx1588), .B1 (nx2796)) ;
    inv01 ix1963 (.Y (nx1964), .A (FilterDout_2__0__2)) ;
    oai32 L0_1_L1_0_Fij_ix243 (.Y (L0_1_L1_0_Fij_nx242), .A0 (nx1966), .A1 (RST)
          , .A2 (nx1958), .B0 (nx1592), .B1 (nx2796)) ;
    inv01 ix1965 (.Y (nx1966), .A (FilterDout_2__0__3)) ;
    oai32 L0_1_L1_0_Fij_ix253 (.Y (L0_1_L1_0_Fij_nx252), .A0 (nx1968), .A1 (RST)
          , .A2 (nx1958), .B0 (nx1596), .B1 (nx2796)) ;
    inv01 ix1967 (.Y (nx1968), .A (FilterDout_2__0__4)) ;
    oai32 L0_1_L1_0_Fij_ix263 (.Y (L0_1_L1_0_Fij_nx262), .A0 (nx1970), .A1 (RST)
          , .A2 (nx1958), .B0 (nx1600), .B1 (nx2796)) ;
    inv01 ix1969 (.Y (nx1970), .A (FilterDout_2__0__5)) ;
    oai32 L0_1_L1_0_Fij_ix273 (.Y (L0_1_L1_0_Fij_nx272), .A0 (nx1972), .A1 (RST)
          , .A2 (nx1974), .B0 (nx1604), .B1 (nx2796)) ;
    inv01 ix1971 (.Y (nx1972), .A (FilterDout_2__0__6)) ;
    inv01 ix1973 (.Y (nx1974), .A (L0_1_L1_0_Fij_nx333)) ;
    oai32 L0_1_L1_0_Fij_ix283 (.Y (L0_1_L1_0_Fij_nx282), .A0 (nx1976), .A1 (RST)
          , .A2 (nx1974), .B0 (nx1610), .B1 (nx2798)) ;
    inv01 ix1975 (.Y (nx1976), .A (FilterDout_2__0__7)) ;
    oai32 L0_1_L1_0_Wij_ix213 (.Y (L0_1_L1_0_Wij_nx212), .A0 (nx1978), .A1 (RST)
          , .A2 (nx1980), .B0 (nx1614), .B1 (nx2800)) ;
    inv01 ix1977 (.Y (nx1978), .A (WindowDout_2__0__0)) ;
    inv02 ix1979 (.Y (nx1980), .A (L0_1_L1_0_Wij_nx331)) ;
    oai32 L0_1_L1_0_Wij_ix223 (.Y (L0_1_L1_0_Wij_nx222), .A0 (nx1984), .A1 (RST)
          , .A2 (nx1980), .B0 (nx1622), .B1 (nx2800)) ;
    inv01 ix1983 (.Y (nx1984), .A (WindowDout_2__0__1)) ;
    oai32 L0_1_L1_0_Wij_ix233 (.Y (L0_1_L1_0_Wij_nx232), .A0 (nx1986), .A1 (RST)
          , .A2 (nx1980), .B0 (nx1626), .B1 (nx2800)) ;
    inv01 ix1985 (.Y (nx1986), .A (WindowDout_2__0__2)) ;
    oai32 L0_1_L1_0_Wij_ix243 (.Y (L0_1_L1_0_Wij_nx242), .A0 (nx1988), .A1 (RST)
          , .A2 (nx1980), .B0 (nx1630), .B1 (nx2800)) ;
    inv01 ix1987 (.Y (nx1988), .A (WindowDout_2__0__3)) ;
    oai32 L0_1_L1_0_Wij_ix253 (.Y (L0_1_L1_0_Wij_nx252), .A0 (nx1990), .A1 (RST)
          , .A2 (nx1980), .B0 (nx1634), .B1 (nx2800)) ;
    inv01 ix1989 (.Y (nx1990), .A (WindowDout_2__0__4)) ;
    oai32 L0_1_L1_0_Wij_ix263 (.Y (L0_1_L1_0_Wij_nx262), .A0 (nx1992), .A1 (RST)
          , .A2 (nx1980), .B0 (nx1638), .B1 (nx2800)) ;
    inv01 ix1991 (.Y (nx1992), .A (WindowDout_2__0__5)) ;
    oai32 L0_1_L1_0_Wij_ix273 (.Y (L0_1_L1_0_Wij_nx272), .A0 (nx1994), .A1 (RST)
          , .A2 (nx1996), .B0 (nx1642), .B1 (nx2800)) ;
    inv01 ix1993 (.Y (nx1994), .A (WindowDout_2__0__6)) ;
    inv01 ix1995 (.Y (nx1996), .A (L0_1_L1_0_Wij_nx333)) ;
    oai32 L0_1_L1_0_Wij_ix283 (.Y (L0_1_L1_0_Wij_nx282), .A0 (nx1998), .A1 (RST)
          , .A2 (nx1996), .B0 (nx1648), .B1 (nx2802)) ;
    inv01 ix1997 (.Y (nx1998), .A (WindowDout_2__0__7)) ;
    oai32 L0_1_L1_1_Fij_ix213 (.Y (L0_1_L1_1_Fij_nx212), .A0 (nx2000), .A1 (RST)
          , .A2 (nx2002), .B0 (nx1652), .B1 (nx2804)) ;
    inv01 ix1999 (.Y (nx2000), .A (FilterDout_2__1__0)) ;
    inv02 ix2001 (.Y (nx2002), .A (L0_1_L1_1_Fij_nx331)) ;
    oai32 L0_1_L1_1_Fij_ix223 (.Y (L0_1_L1_1_Fij_nx222), .A0 (nx2006), .A1 (RST)
          , .A2 (nx2002), .B0 (nx1660), .B1 (nx2804)) ;
    inv01 ix2005 (.Y (nx2006), .A (FilterDout_2__1__1)) ;
    oai32 L0_1_L1_1_Fij_ix233 (.Y (L0_1_L1_1_Fij_nx232), .A0 (nx2008), .A1 (RST)
          , .A2 (nx2002), .B0 (nx1664), .B1 (nx2804)) ;
    inv01 ix2007 (.Y (nx2008), .A (FilterDout_2__1__2)) ;
    oai32 L0_1_L1_1_Fij_ix243 (.Y (L0_1_L1_1_Fij_nx242), .A0 (nx2010), .A1 (RST)
          , .A2 (nx2002), .B0 (nx1668), .B1 (nx2804)) ;
    inv01 ix2009 (.Y (nx2010), .A (FilterDout_2__1__3)) ;
    oai32 L0_1_L1_1_Fij_ix253 (.Y (L0_1_L1_1_Fij_nx252), .A0 (nx2012), .A1 (RST)
          , .A2 (nx2002), .B0 (nx1672), .B1 (nx2804)) ;
    inv01 ix2011 (.Y (nx2012), .A (FilterDout_2__1__4)) ;
    oai32 L0_1_L1_1_Fij_ix263 (.Y (L0_1_L1_1_Fij_nx262), .A0 (nx2014), .A1 (RST)
          , .A2 (nx2002), .B0 (nx1676), .B1 (nx2804)) ;
    inv01 ix2013 (.Y (nx2014), .A (FilterDout_2__1__5)) ;
    oai32 L0_1_L1_1_Fij_ix273 (.Y (L0_1_L1_1_Fij_nx272), .A0 (nx2016), .A1 (RST)
          , .A2 (nx2018), .B0 (nx1680), .B1 (nx2804)) ;
    inv01 ix2015 (.Y (nx2016), .A (FilterDout_2__1__6)) ;
    inv01 ix2017 (.Y (nx2018), .A (L0_1_L1_1_Fij_nx333)) ;
    oai32 L0_1_L1_1_Fij_ix283 (.Y (L0_1_L1_1_Fij_nx282), .A0 (nx2020), .A1 (RST)
          , .A2 (nx2018), .B0 (nx1686), .B1 (nx2806)) ;
    inv01 ix2019 (.Y (nx2020), .A (FilterDout_2__1__7)) ;
    oai32 L0_1_L1_1_Wij_ix213 (.Y (L0_1_L1_1_Wij_nx212), .A0 (nx2022), .A1 (RST)
          , .A2 (nx2024), .B0 (nx1690), .B1 (nx2808)) ;
    inv01 ix2021 (.Y (nx2022), .A (WindowDout_2__1__0)) ;
    inv02 ix2023 (.Y (nx2024), .A (L0_1_L1_1_Wij_nx331)) ;
    oai32 L0_1_L1_1_Wij_ix223 (.Y (L0_1_L1_1_Wij_nx222), .A0 (nx2028), .A1 (RST)
          , .A2 (nx2024), .B0 (nx1698), .B1 (nx2808)) ;
    inv01 ix2027 (.Y (nx2028), .A (WindowDout_2__1__1)) ;
    oai32 L0_1_L1_1_Wij_ix233 (.Y (L0_1_L1_1_Wij_nx232), .A0 (nx2030), .A1 (RST)
          , .A2 (nx2024), .B0 (nx1702), .B1 (nx2808)) ;
    inv01 ix2029 (.Y (nx2030), .A (WindowDout_2__1__2)) ;
    oai32 L0_1_L1_1_Wij_ix243 (.Y (L0_1_L1_1_Wij_nx242), .A0 (nx2032), .A1 (RST)
          , .A2 (nx2024), .B0 (nx1706), .B1 (nx2808)) ;
    inv01 ix2031 (.Y (nx2032), .A (WindowDout_2__1__3)) ;
    oai32 L0_1_L1_1_Wij_ix253 (.Y (L0_1_L1_1_Wij_nx252), .A0 (nx2034), .A1 (RST)
          , .A2 (nx2024), .B0 (nx1710), .B1 (nx2808)) ;
    inv01 ix2033 (.Y (nx2034), .A (WindowDout_2__1__4)) ;
    oai32 L0_1_L1_1_Wij_ix263 (.Y (L0_1_L1_1_Wij_nx262), .A0 (nx2036), .A1 (RST)
          , .A2 (nx2024), .B0 (nx1714), .B1 (nx2808)) ;
    inv01 ix2035 (.Y (nx2036), .A (WindowDout_2__1__5)) ;
    oai32 L0_1_L1_1_Wij_ix273 (.Y (L0_1_L1_1_Wij_nx272), .A0 (nx2038), .A1 (RST)
          , .A2 (nx2040), .B0 (nx1718), .B1 (nx2808)) ;
    inv01 ix2037 (.Y (nx2038), .A (WindowDout_2__1__6)) ;
    inv01 ix2039 (.Y (nx2040), .A (L0_1_L1_1_Wij_nx333)) ;
    oai32 L0_1_L1_1_Wij_ix283 (.Y (L0_1_L1_1_Wij_nx282), .A0 (nx2042), .A1 (RST)
          , .A2 (nx2040), .B0 (nx1724), .B1 (nx2810)) ;
    inv01 ix2041 (.Y (nx2042), .A (WindowDout_2__1__7)) ;
    oai32 L0_1_L1_2_Fij_ix213 (.Y (L0_1_L1_2_Fij_nx212), .A0 (nx2044), .A1 (RST)
          , .A2 (nx2046), .B0 (nx1728), .B1 (nx2812)) ;
    inv01 ix2043 (.Y (nx2044), .A (FilterDout_2__2__0)) ;
    inv02 ix2045 (.Y (nx2046), .A (L0_1_L1_2_Fij_nx331)) ;
    oai32 L0_1_L1_2_Fij_ix223 (.Y (L0_1_L1_2_Fij_nx222), .A0 (nx2050), .A1 (RST)
          , .A2 (nx2046), .B0 (nx1736), .B1 (nx2812)) ;
    inv01 ix2049 (.Y (nx2050), .A (FilterDout_2__2__1)) ;
    oai32 L0_1_L1_2_Fij_ix233 (.Y (L0_1_L1_2_Fij_nx232), .A0 (nx2052), .A1 (RST)
          , .A2 (nx2046), .B0 (nx1740), .B1 (nx2812)) ;
    inv01 ix2051 (.Y (nx2052), .A (FilterDout_2__2__2)) ;
    oai32 L0_1_L1_2_Fij_ix243 (.Y (L0_1_L1_2_Fij_nx242), .A0 (nx2054), .A1 (RST)
          , .A2 (nx2046), .B0 (nx1744), .B1 (nx2812)) ;
    inv01 ix2053 (.Y (nx2054), .A (FilterDout_2__2__3)) ;
    oai32 L0_1_L1_2_Fij_ix253 (.Y (L0_1_L1_2_Fij_nx252), .A0 (nx2056), .A1 (RST)
          , .A2 (nx2046), .B0 (nx1748), .B1 (nx2812)) ;
    inv01 ix2055 (.Y (nx2056), .A (FilterDout_2__2__4)) ;
    oai32 L0_1_L1_2_Fij_ix263 (.Y (L0_1_L1_2_Fij_nx262), .A0 (nx2058), .A1 (RST)
          , .A2 (nx2046), .B0 (nx1752), .B1 (nx2812)) ;
    inv01 ix2057 (.Y (nx2058), .A (FilterDout_2__2__5)) ;
    oai32 L0_1_L1_2_Fij_ix273 (.Y (L0_1_L1_2_Fij_nx272), .A0 (nx2060), .A1 (RST)
          , .A2 (nx2062), .B0 (nx1756), .B1 (nx2812)) ;
    inv01 ix2059 (.Y (nx2060), .A (FilterDout_2__2__6)) ;
    inv01 ix2061 (.Y (nx2062), .A (L0_1_L1_2_Fij_nx333)) ;
    oai32 L0_1_L1_2_Fij_ix283 (.Y (L0_1_L1_2_Fij_nx282), .A0 (nx2064), .A1 (RST)
          , .A2 (nx2062), .B0 (nx1762), .B1 (nx2814)) ;
    inv01 ix2063 (.Y (nx2064), .A (FilterDout_2__2__7)) ;
    oai32 L0_1_L1_2_Wij_ix213 (.Y (L0_1_L1_2_Wij_nx212), .A0 (nx2066), .A1 (RST)
          , .A2 (nx2068), .B0 (nx1766), .B1 (nx2816)) ;
    inv01 ix2065 (.Y (nx2066), .A (WindowDout_2__2__0)) ;
    inv02 ix2067 (.Y (nx2068), .A (L0_1_L1_2_Wij_nx331)) ;
    oai32 L0_1_L1_2_Wij_ix223 (.Y (L0_1_L1_2_Wij_nx222), .A0 (nx2072), .A1 (RST)
          , .A2 (nx2068), .B0 (nx1774), .B1 (nx2816)) ;
    inv01 ix2071 (.Y (nx2072), .A (WindowDout_2__2__1)) ;
    oai32 L0_1_L1_2_Wij_ix233 (.Y (L0_1_L1_2_Wij_nx232), .A0 (nx2074), .A1 (RST)
          , .A2 (nx2068), .B0 (nx1778), .B1 (nx2816)) ;
    inv01 ix2073 (.Y (nx2074), .A (WindowDout_2__2__2)) ;
    oai32 L0_1_L1_2_Wij_ix243 (.Y (L0_1_L1_2_Wij_nx242), .A0 (nx2076), .A1 (RST)
          , .A2 (nx2068), .B0 (nx1782), .B1 (nx2816)) ;
    inv01 ix2075 (.Y (nx2076), .A (WindowDout_2__2__3)) ;
    oai32 L0_1_L1_2_Wij_ix253 (.Y (L0_1_L1_2_Wij_nx252), .A0 (nx2078), .A1 (RST)
          , .A2 (nx2068), .B0 (nx1786), .B1 (nx2816)) ;
    inv01 ix2077 (.Y (nx2078), .A (WindowDout_2__2__4)) ;
    oai32 L0_1_L1_2_Wij_ix263 (.Y (L0_1_L1_2_Wij_nx262), .A0 (nx2080), .A1 (RST)
          , .A2 (nx2068), .B0 (nx1790), .B1 (nx2816)) ;
    inv01 ix2079 (.Y (nx2080), .A (WindowDout_2__2__5)) ;
    oai32 L0_1_L1_2_Wij_ix273 (.Y (L0_1_L1_2_Wij_nx272), .A0 (nx2082), .A1 (RST)
          , .A2 (nx2084), .B0 (nx1794), .B1 (nx2816)) ;
    inv01 ix2081 (.Y (nx2082), .A (WindowDout_2__2__6)) ;
    inv01 ix2083 (.Y (nx2084), .A (L0_1_L1_2_Wij_nx333)) ;
    oai32 L0_1_L1_2_Wij_ix283 (.Y (L0_1_L1_2_Wij_nx282), .A0 (nx2086), .A1 (RST)
          , .A2 (nx2084), .B0 (nx1800), .B1 (nx2818)) ;
    inv01 ix2085 (.Y (nx2086), .A (WindowDout_2__2__7)) ;
    oai32 L0_1_L1_3_Fij_ix213 (.Y (L0_1_L1_3_Fij_nx212), .A0 (nx2088), .A1 (RST)
          , .A2 (nx2090), .B0 (nx1804), .B1 (nx2820)) ;
    inv01 ix2087 (.Y (nx2088), .A (FilterDout_2__3__0)) ;
    inv02 ix2089 (.Y (nx2090), .A (L0_1_L1_3_Fij_nx331)) ;
    oai32 L0_1_L1_3_Fij_ix223 (.Y (L0_1_L1_3_Fij_nx222), .A0 (nx2094), .A1 (RST)
          , .A2 (nx2090), .B0 (nx1812), .B1 (nx2820)) ;
    inv01 ix2093 (.Y (nx2094), .A (FilterDout_2__3__1)) ;
    oai32 L0_1_L1_3_Fij_ix233 (.Y (L0_1_L1_3_Fij_nx232), .A0 (nx2096), .A1 (RST)
          , .A2 (nx2090), .B0 (nx1816), .B1 (nx2820)) ;
    inv01 ix2095 (.Y (nx2096), .A (FilterDout_2__3__2)) ;
    oai32 L0_1_L1_3_Fij_ix243 (.Y (L0_1_L1_3_Fij_nx242), .A0 (nx2098), .A1 (RST)
          , .A2 (nx2090), .B0 (nx1820), .B1 (nx2820)) ;
    inv01 ix2097 (.Y (nx2098), .A (FilterDout_2__3__3)) ;
    oai32 L0_1_L1_3_Fij_ix253 (.Y (L0_1_L1_3_Fij_nx252), .A0 (nx2100), .A1 (RST)
          , .A2 (nx2090), .B0 (nx1824), .B1 (nx2820)) ;
    inv01 ix2099 (.Y (nx2100), .A (FilterDout_2__3__4)) ;
    oai32 L0_1_L1_3_Fij_ix263 (.Y (L0_1_L1_3_Fij_nx262), .A0 (nx2102), .A1 (RST)
          , .A2 (nx2090), .B0 (nx1828), .B1 (nx2820)) ;
    inv01 ix2101 (.Y (nx2102), .A (FilterDout_2__3__5)) ;
    oai32 L0_1_L1_3_Fij_ix273 (.Y (L0_1_L1_3_Fij_nx272), .A0 (nx2104), .A1 (RST)
          , .A2 (nx2106), .B0 (nx1832), .B1 (nx2820)) ;
    inv01 ix2103 (.Y (nx2104), .A (FilterDout_2__3__6)) ;
    inv01 ix2105 (.Y (nx2106), .A (L0_1_L1_3_Fij_nx333)) ;
    oai32 L0_1_L1_3_Fij_ix283 (.Y (L0_1_L1_3_Fij_nx282), .A0 (nx2108), .A1 (RST)
          , .A2 (nx2106), .B0 (nx1838), .B1 (nx2822)) ;
    inv01 ix2107 (.Y (nx2108), .A (FilterDout_2__3__7)) ;
    oai32 L0_1_L1_3_Wij_ix213 (.Y (L0_1_L1_3_Wij_nx212), .A0 (nx2110), .A1 (RST)
          , .A2 (nx2112), .B0 (nx1842), .B1 (nx2824)) ;
    inv01 ix2109 (.Y (nx2110), .A (WindowDout_2__3__0)) ;
    inv02 ix2111 (.Y (nx2112), .A (L0_1_L1_3_Wij_nx331)) ;
    oai32 L0_1_L1_3_Wij_ix223 (.Y (L0_1_L1_3_Wij_nx222), .A0 (nx2116), .A1 (RST)
          , .A2 (nx2112), .B0 (nx1850), .B1 (nx2824)) ;
    inv01 ix2115 (.Y (nx2116), .A (WindowDout_2__3__1)) ;
    oai32 L0_1_L1_3_Wij_ix233 (.Y (L0_1_L1_3_Wij_nx232), .A0 (nx2118), .A1 (RST)
          , .A2 (nx2112), .B0 (nx1854), .B1 (nx2824)) ;
    inv01 ix2117 (.Y (nx2118), .A (WindowDout_2__3__2)) ;
    oai32 L0_1_L1_3_Wij_ix243 (.Y (L0_1_L1_3_Wij_nx242), .A0 (nx2120), .A1 (RST)
          , .A2 (nx2112), .B0 (nx1858), .B1 (nx2824)) ;
    inv01 ix2119 (.Y (nx2120), .A (WindowDout_2__3__3)) ;
    oai32 L0_1_L1_3_Wij_ix253 (.Y (L0_1_L1_3_Wij_nx252), .A0 (nx2122), .A1 (RST)
          , .A2 (nx2112), .B0 (nx1862), .B1 (nx2824)) ;
    inv01 ix2121 (.Y (nx2122), .A (WindowDout_2__3__4)) ;
    oai32 L0_1_L1_3_Wij_ix263 (.Y (L0_1_L1_3_Wij_nx262), .A0 (nx2124), .A1 (RST)
          , .A2 (nx2112), .B0 (nx1866), .B1 (nx2824)) ;
    inv01 ix2123 (.Y (nx2124), .A (WindowDout_2__3__5)) ;
    oai32 L0_1_L1_3_Wij_ix273 (.Y (L0_1_L1_3_Wij_nx272), .A0 (nx2126), .A1 (RST)
          , .A2 (nx2128), .B0 (nx1870), .B1 (nx2824)) ;
    inv01 ix2125 (.Y (nx2126), .A (WindowDout_2__3__6)) ;
    inv01 ix2127 (.Y (nx2128), .A (L0_1_L1_3_Wij_nx333)) ;
    oai32 L0_1_L1_3_Wij_ix283 (.Y (L0_1_L1_3_Wij_nx282), .A0 (nx2130), .A1 (RST)
          , .A2 (nx2128), .B0 (nx1876), .B1 (nx2826)) ;
    inv01 ix2129 (.Y (nx2130), .A (WindowDout_2__3__7)) ;
    oai32 L0_1_L1_4_Fij_ix213 (.Y (L0_1_L1_4_Fij_nx212), .A0 (nx2132), .A1 (RST)
          , .A2 (nx2134), .B0 (nx1880), .B1 (nx2828)) ;
    inv01 ix2131 (.Y (nx2132), .A (FilterDout_2__4__0)) ;
    inv02 ix2133 (.Y (nx2134), .A (L0_1_L1_4_Fij_nx331)) ;
    oai32 L0_1_L1_4_Fij_ix223 (.Y (L0_1_L1_4_Fij_nx222), .A0 (nx2138), .A1 (RST)
          , .A2 (nx2134), .B0 (nx1888), .B1 (nx2828)) ;
    inv01 ix2137 (.Y (nx2138), .A (FilterDout_2__4__1)) ;
    oai32 L0_1_L1_4_Fij_ix233 (.Y (L0_1_L1_4_Fij_nx232), .A0 (nx2140), .A1 (RST)
          , .A2 (nx2134), .B0 (nx1892), .B1 (nx2828)) ;
    inv01 ix2139 (.Y (nx2140), .A (FilterDout_2__4__2)) ;
    oai32 L0_1_L1_4_Fij_ix243 (.Y (L0_1_L1_4_Fij_nx242), .A0 (nx2142), .A1 (RST)
          , .A2 (nx2134), .B0 (nx1896), .B1 (nx2828)) ;
    inv01 ix2141 (.Y (nx2142), .A (FilterDout_2__4__3)) ;
    oai32 L0_1_L1_4_Fij_ix253 (.Y (L0_1_L1_4_Fij_nx252), .A0 (nx2144), .A1 (RST)
          , .A2 (nx2134), .B0 (nx1900), .B1 (nx2828)) ;
    inv01 ix2143 (.Y (nx2144), .A (FilterDout_2__4__4)) ;
    oai32 L0_1_L1_4_Fij_ix263 (.Y (L0_1_L1_4_Fij_nx262), .A0 (nx2146), .A1 (RST)
          , .A2 (nx2134), .B0 (nx1904), .B1 (nx2828)) ;
    inv01 ix2145 (.Y (nx2146), .A (FilterDout_2__4__5)) ;
    oai32 L0_1_L1_4_Fij_ix273 (.Y (L0_1_L1_4_Fij_nx272), .A0 (nx2148), .A1 (RST)
          , .A2 (nx2150), .B0 (nx1908), .B1 (nx2828)) ;
    inv01 ix2147 (.Y (nx2148), .A (FilterDout_2__4__6)) ;
    inv01 ix2149 (.Y (nx2150), .A (L0_1_L1_4_Fij_nx333)) ;
    oai32 L0_1_L1_4_Fij_ix283 (.Y (L0_1_L1_4_Fij_nx282), .A0 (nx2152), .A1 (RST)
          , .A2 (nx2150), .B0 (nx1914), .B1 (nx2830)) ;
    inv01 ix2151 (.Y (nx2152), .A (FilterDout_2__4__7)) ;
    oai32 L0_1_L1_4_Wij_ix213 (.Y (L0_1_L1_4_Wij_nx212), .A0 (nx2154), .A1 (RST)
          , .A2 (nx2156), .B0 (nx1918), .B1 (nx2832)) ;
    inv01 ix2153 (.Y (nx2154), .A (WindowDout_2__4__0)) ;
    inv02 ix2155 (.Y (nx2156), .A (L0_1_L1_4_Wij_nx331)) ;
    oai32 L0_1_L1_4_Wij_ix223 (.Y (L0_1_L1_4_Wij_nx222), .A0 (nx2160), .A1 (RST)
          , .A2 (nx2156), .B0 (nx1926), .B1 (nx2832)) ;
    inv01 ix2159 (.Y (nx2160), .A (WindowDout_2__4__1)) ;
    oai32 L0_1_L1_4_Wij_ix233 (.Y (L0_1_L1_4_Wij_nx232), .A0 (nx2162), .A1 (RST)
          , .A2 (nx2156), .B0 (nx1930), .B1 (nx2832)) ;
    inv01 ix2161 (.Y (nx2162), .A (WindowDout_2__4__2)) ;
    oai32 L0_1_L1_4_Wij_ix243 (.Y (L0_1_L1_4_Wij_nx242), .A0 (nx2164), .A1 (RST)
          , .A2 (nx2156), .B0 (nx1934), .B1 (nx2832)) ;
    inv01 ix2163 (.Y (nx2164), .A (WindowDout_2__4__3)) ;
    oai32 L0_1_L1_4_Wij_ix253 (.Y (L0_1_L1_4_Wij_nx252), .A0 (nx2166), .A1 (RST)
          , .A2 (nx2156), .B0 (nx1938), .B1 (nx2832)) ;
    inv01 ix2165 (.Y (nx2166), .A (WindowDout_2__4__4)) ;
    oai32 L0_1_L1_4_Wij_ix263 (.Y (L0_1_L1_4_Wij_nx262), .A0 (nx2168), .A1 (RST)
          , .A2 (nx2156), .B0 (nx1942), .B1 (nx2832)) ;
    inv01 ix2167 (.Y (nx2168), .A (WindowDout_2__4__5)) ;
    oai32 L0_1_L1_4_Wij_ix273 (.Y (L0_1_L1_4_Wij_nx272), .A0 (nx2170), .A1 (RST)
          , .A2 (nx2172), .B0 (nx1946), .B1 (nx2832)) ;
    inv01 ix2169 (.Y (nx2170), .A (WindowDout_2__4__6)) ;
    inv01 ix2171 (.Y (nx2172), .A (L0_1_L1_4_Wij_nx333)) ;
    oai32 L0_1_L1_4_Wij_ix283 (.Y (L0_1_L1_4_Wij_nx282), .A0 (nx2174), .A1 (RST)
          , .A2 (nx2172), .B0 (nx1952), .B1 (nx2834)) ;
    inv01 ix2173 (.Y (nx2174), .A (WindowDout_2__4__7)) ;
    oai32 L0_2_L1_0_Fij_ix213 (.Y (L0_2_L1_0_Fij_nx212), .A0 (nx2176), .A1 (RST)
          , .A2 (nx2178), .B0 (nx1956), .B1 (nx2836)) ;
    inv01 ix2175 (.Y (nx2176), .A (FilterDout_3__0__0)) ;
    inv02 ix2177 (.Y (nx2178), .A (L0_2_L1_0_Fij_nx331)) ;
    oai32 L0_2_L1_0_Fij_ix223 (.Y (L0_2_L1_0_Fij_nx222), .A0 (nx2182), .A1 (RST)
          , .A2 (nx2178), .B0 (nx1962), .B1 (nx2836)) ;
    inv01 ix2181 (.Y (nx2182), .A (FilterDout_3__0__1)) ;
    oai32 L0_2_L1_0_Fij_ix233 (.Y (L0_2_L1_0_Fij_nx232), .A0 (nx2184), .A1 (RST)
          , .A2 (nx2178), .B0 (nx1964), .B1 (nx2836)) ;
    inv01 ix2183 (.Y (nx2184), .A (FilterDout_3__0__2)) ;
    oai32 L0_2_L1_0_Fij_ix243 (.Y (L0_2_L1_0_Fij_nx242), .A0 (nx2186), .A1 (RST)
          , .A2 (nx2178), .B0 (nx1966), .B1 (nx2836)) ;
    inv01 ix2185 (.Y (nx2186), .A (FilterDout_3__0__3)) ;
    oai32 L0_2_L1_0_Fij_ix253 (.Y (L0_2_L1_0_Fij_nx252), .A0 (nx2188), .A1 (RST)
          , .A2 (nx2178), .B0 (nx1968), .B1 (nx2836)) ;
    inv01 ix2187 (.Y (nx2188), .A (FilterDout_3__0__4)) ;
    oai32 L0_2_L1_0_Fij_ix263 (.Y (L0_2_L1_0_Fij_nx262), .A0 (nx2190), .A1 (RST)
          , .A2 (nx2178), .B0 (nx1970), .B1 (nx2836)) ;
    inv01 ix2189 (.Y (nx2190), .A (FilterDout_3__0__5)) ;
    oai32 L0_2_L1_0_Fij_ix273 (.Y (L0_2_L1_0_Fij_nx272), .A0 (nx2192), .A1 (RST)
          , .A2 (nx2194), .B0 (nx1972), .B1 (nx2836)) ;
    inv01 ix2191 (.Y (nx2192), .A (FilterDout_3__0__6)) ;
    inv01 ix2193 (.Y (nx2194), .A (L0_2_L1_0_Fij_nx333)) ;
    oai32 L0_2_L1_0_Fij_ix283 (.Y (L0_2_L1_0_Fij_nx282), .A0 (nx2196), .A1 (RST)
          , .A2 (nx2194), .B0 (nx1976), .B1 (nx2838)) ;
    inv01 ix2195 (.Y (nx2196), .A (FilterDout_3__0__7)) ;
    oai32 L0_2_L1_0_Wij_ix213 (.Y (L0_2_L1_0_Wij_nx212), .A0 (nx2198), .A1 (RST)
          , .A2 (nx2200), .B0 (nx1978), .B1 (nx2840)) ;
    inv01 ix2197 (.Y (nx2198), .A (WindowDout_3__0__0)) ;
    inv02 ix2199 (.Y (nx2200), .A (L0_2_L1_0_Wij_nx331)) ;
    oai32 L0_2_L1_0_Wij_ix223 (.Y (L0_2_L1_0_Wij_nx222), .A0 (nx2204), .A1 (RST)
          , .A2 (nx2200), .B0 (nx1984), .B1 (nx2840)) ;
    inv01 ix2203 (.Y (nx2204), .A (WindowDout_3__0__1)) ;
    oai32 L0_2_L1_0_Wij_ix233 (.Y (L0_2_L1_0_Wij_nx232), .A0 (nx2206), .A1 (RST)
          , .A2 (nx2200), .B0 (nx1986), .B1 (nx2840)) ;
    inv01 ix2205 (.Y (nx2206), .A (WindowDout_3__0__2)) ;
    oai32 L0_2_L1_0_Wij_ix243 (.Y (L0_2_L1_0_Wij_nx242), .A0 (nx2208), .A1 (RST)
          , .A2 (nx2200), .B0 (nx1988), .B1 (nx2840)) ;
    inv01 ix2207 (.Y (nx2208), .A (WindowDout_3__0__3)) ;
    oai32 L0_2_L1_0_Wij_ix253 (.Y (L0_2_L1_0_Wij_nx252), .A0 (nx2210), .A1 (RST)
          , .A2 (nx2200), .B0 (nx1990), .B1 (nx2840)) ;
    inv01 ix2209 (.Y (nx2210), .A (WindowDout_3__0__4)) ;
    oai32 L0_2_L1_0_Wij_ix263 (.Y (L0_2_L1_0_Wij_nx262), .A0 (nx2212), .A1 (RST)
          , .A2 (nx2200), .B0 (nx1992), .B1 (nx2840)) ;
    inv01 ix2211 (.Y (nx2212), .A (WindowDout_3__0__5)) ;
    oai32 L0_2_L1_0_Wij_ix273 (.Y (L0_2_L1_0_Wij_nx272), .A0 (nx2214), .A1 (RST)
          , .A2 (nx2216), .B0 (nx1994), .B1 (nx2840)) ;
    inv01 ix2213 (.Y (nx2214), .A (WindowDout_3__0__6)) ;
    inv01 ix2215 (.Y (nx2216), .A (L0_2_L1_0_Wij_nx333)) ;
    oai32 L0_2_L1_0_Wij_ix283 (.Y (L0_2_L1_0_Wij_nx282), .A0 (nx2218), .A1 (RST)
          , .A2 (nx2216), .B0 (nx1998), .B1 (nx2842)) ;
    inv01 ix2217 (.Y (nx2218), .A (WindowDout_3__0__7)) ;
    oai32 L0_2_L1_1_Fij_ix213 (.Y (L0_2_L1_1_Fij_nx212), .A0 (nx2220), .A1 (RST)
          , .A2 (nx2222), .B0 (nx2000), .B1 (nx2844)) ;
    inv01 ix2219 (.Y (nx2220), .A (FilterDout_3__1__0)) ;
    inv02 ix2221 (.Y (nx2222), .A (L0_2_L1_1_Fij_nx331)) ;
    oai32 L0_2_L1_1_Fij_ix223 (.Y (L0_2_L1_1_Fij_nx222), .A0 (nx2226), .A1 (RST)
          , .A2 (nx2222), .B0 (nx2006), .B1 (nx2844)) ;
    inv01 ix2225 (.Y (nx2226), .A (FilterDout_3__1__1)) ;
    oai32 L0_2_L1_1_Fij_ix233 (.Y (L0_2_L1_1_Fij_nx232), .A0 (nx2228), .A1 (RST)
          , .A2 (nx2222), .B0 (nx2008), .B1 (nx2844)) ;
    inv01 ix2227 (.Y (nx2228), .A (FilterDout_3__1__2)) ;
    oai32 L0_2_L1_1_Fij_ix243 (.Y (L0_2_L1_1_Fij_nx242), .A0 (nx2230), .A1 (RST)
          , .A2 (nx2222), .B0 (nx2010), .B1 (nx2844)) ;
    inv01 ix2229 (.Y (nx2230), .A (FilterDout_3__1__3)) ;
    oai32 L0_2_L1_1_Fij_ix253 (.Y (L0_2_L1_1_Fij_nx252), .A0 (nx2232), .A1 (RST)
          , .A2 (nx2222), .B0 (nx2012), .B1 (nx2844)) ;
    inv01 ix2231 (.Y (nx2232), .A (FilterDout_3__1__4)) ;
    oai32 L0_2_L1_1_Fij_ix263 (.Y (L0_2_L1_1_Fij_nx262), .A0 (nx2234), .A1 (RST)
          , .A2 (nx2222), .B0 (nx2014), .B1 (nx2844)) ;
    inv01 ix2233 (.Y (nx2234), .A (FilterDout_3__1__5)) ;
    oai32 L0_2_L1_1_Fij_ix273 (.Y (L0_2_L1_1_Fij_nx272), .A0 (nx2236), .A1 (RST)
          , .A2 (nx2238), .B0 (nx2016), .B1 (nx2844)) ;
    inv01 ix2235 (.Y (nx2236), .A (FilterDout_3__1__6)) ;
    inv01 ix2237 (.Y (nx2238), .A (L0_2_L1_1_Fij_nx333)) ;
    oai32 L0_2_L1_1_Fij_ix283 (.Y (L0_2_L1_1_Fij_nx282), .A0 (nx2240), .A1 (RST)
          , .A2 (nx2238), .B0 (nx2020), .B1 (nx2846)) ;
    inv01 ix2239 (.Y (nx2240), .A (FilterDout_3__1__7)) ;
    oai32 L0_2_L1_1_Wij_ix213 (.Y (L0_2_L1_1_Wij_nx212), .A0 (nx2242), .A1 (RST)
          , .A2 (nx2244), .B0 (nx2022), .B1 (nx2848)) ;
    inv01 ix2241 (.Y (nx2242), .A (WindowDout_3__1__0)) ;
    inv02 ix2243 (.Y (nx2244), .A (L0_2_L1_1_Wij_nx331)) ;
    oai32 L0_2_L1_1_Wij_ix223 (.Y (L0_2_L1_1_Wij_nx222), .A0 (nx2248), .A1 (RST)
          , .A2 (nx2244), .B0 (nx2028), .B1 (nx2848)) ;
    inv01 ix2247 (.Y (nx2248), .A (WindowDout_3__1__1)) ;
    oai32 L0_2_L1_1_Wij_ix233 (.Y (L0_2_L1_1_Wij_nx232), .A0 (nx2250), .A1 (RST)
          , .A2 (nx2244), .B0 (nx2030), .B1 (nx2848)) ;
    inv01 ix2249 (.Y (nx2250), .A (WindowDout_3__1__2)) ;
    oai32 L0_2_L1_1_Wij_ix243 (.Y (L0_2_L1_1_Wij_nx242), .A0 (nx2252), .A1 (RST)
          , .A2 (nx2244), .B0 (nx2032), .B1 (nx2848)) ;
    inv01 ix2251 (.Y (nx2252), .A (WindowDout_3__1__3)) ;
    oai32 L0_2_L1_1_Wij_ix253 (.Y (L0_2_L1_1_Wij_nx252), .A0 (nx2254), .A1 (RST)
          , .A2 (nx2244), .B0 (nx2034), .B1 (nx2848)) ;
    inv01 ix2253 (.Y (nx2254), .A (WindowDout_3__1__4)) ;
    oai32 L0_2_L1_1_Wij_ix263 (.Y (L0_2_L1_1_Wij_nx262), .A0 (nx2256), .A1 (RST)
          , .A2 (nx2244), .B0 (nx2036), .B1 (nx2848)) ;
    inv01 ix2255 (.Y (nx2256), .A (WindowDout_3__1__5)) ;
    oai32 L0_2_L1_1_Wij_ix273 (.Y (L0_2_L1_1_Wij_nx272), .A0 (nx2258), .A1 (RST)
          , .A2 (nx2260), .B0 (nx2038), .B1 (nx2848)) ;
    inv01 ix2257 (.Y (nx2258), .A (WindowDout_3__1__6)) ;
    inv01 ix2259 (.Y (nx2260), .A (L0_2_L1_1_Wij_nx333)) ;
    oai32 L0_2_L1_1_Wij_ix283 (.Y (L0_2_L1_1_Wij_nx282), .A0 (nx2262), .A1 (RST)
          , .A2 (nx2260), .B0 (nx2042), .B1 (nx2850)) ;
    inv01 ix2261 (.Y (nx2262), .A (WindowDout_3__1__7)) ;
    oai32 L0_2_L1_2_Fij_ix213 (.Y (L0_2_L1_2_Fij_nx212), .A0 (nx2264), .A1 (RST)
          , .A2 (nx2266), .B0 (nx2044), .B1 (nx2852)) ;
    inv01 ix2263 (.Y (nx2264), .A (FilterDout_3__2__0)) ;
    inv02 ix2265 (.Y (nx2266), .A (L0_2_L1_2_Fij_nx331)) ;
    oai32 L0_2_L1_2_Fij_ix223 (.Y (L0_2_L1_2_Fij_nx222), .A0 (nx2270), .A1 (RST)
          , .A2 (nx2266), .B0 (nx2050), .B1 (nx2852)) ;
    inv01 ix2269 (.Y (nx2270), .A (FilterDout_3__2__1)) ;
    oai32 L0_2_L1_2_Fij_ix233 (.Y (L0_2_L1_2_Fij_nx232), .A0 (nx2272), .A1 (RST)
          , .A2 (nx2266), .B0 (nx2052), .B1 (nx2852)) ;
    inv01 ix2271 (.Y (nx2272), .A (FilterDout_3__2__2)) ;
    oai32 L0_2_L1_2_Fij_ix243 (.Y (L0_2_L1_2_Fij_nx242), .A0 (nx2274), .A1 (RST)
          , .A2 (nx2266), .B0 (nx2054), .B1 (nx2852)) ;
    inv01 ix2273 (.Y (nx2274), .A (FilterDout_3__2__3)) ;
    oai32 L0_2_L1_2_Fij_ix253 (.Y (L0_2_L1_2_Fij_nx252), .A0 (nx2276), .A1 (RST)
          , .A2 (nx2266), .B0 (nx2056), .B1 (nx2852)) ;
    inv01 ix2275 (.Y (nx2276), .A (FilterDout_3__2__4)) ;
    oai32 L0_2_L1_2_Fij_ix263 (.Y (L0_2_L1_2_Fij_nx262), .A0 (nx2278), .A1 (RST)
          , .A2 (nx2266), .B0 (nx2058), .B1 (nx2852)) ;
    inv01 ix2277 (.Y (nx2278), .A (FilterDout_3__2__5)) ;
    oai32 L0_2_L1_2_Fij_ix273 (.Y (L0_2_L1_2_Fij_nx272), .A0 (nx2280), .A1 (RST)
          , .A2 (nx2282), .B0 (nx2060), .B1 (nx2852)) ;
    inv01 ix2279 (.Y (nx2280), .A (FilterDout_3__2__6)) ;
    inv01 ix2281 (.Y (nx2282), .A (L0_2_L1_2_Fij_nx333)) ;
    oai32 L0_2_L1_2_Fij_ix283 (.Y (L0_2_L1_2_Fij_nx282), .A0 (nx2284), .A1 (RST)
          , .A2 (nx2282), .B0 (nx2064), .B1 (nx2854)) ;
    inv01 ix2283 (.Y (nx2284), .A (FilterDout_3__2__7)) ;
    oai32 L0_2_L1_2_Wij_ix213 (.Y (L0_2_L1_2_Wij_nx212), .A0 (nx2286), .A1 (RST)
          , .A2 (nx2288), .B0 (nx2066), .B1 (nx2856)) ;
    inv01 ix2285 (.Y (nx2286), .A (WindowDout_3__2__0)) ;
    inv02 ix2287 (.Y (nx2288), .A (L0_2_L1_2_Wij_nx331)) ;
    oai32 L0_2_L1_2_Wij_ix223 (.Y (L0_2_L1_2_Wij_nx222), .A0 (nx2292), .A1 (RST)
          , .A2 (nx2288), .B0 (nx2072), .B1 (nx2856)) ;
    inv01 ix2291 (.Y (nx2292), .A (WindowDout_3__2__1)) ;
    oai32 L0_2_L1_2_Wij_ix233 (.Y (L0_2_L1_2_Wij_nx232), .A0 (nx2294), .A1 (RST)
          , .A2 (nx2288), .B0 (nx2074), .B1 (nx2856)) ;
    inv01 ix2293 (.Y (nx2294), .A (WindowDout_3__2__2)) ;
    oai32 L0_2_L1_2_Wij_ix243 (.Y (L0_2_L1_2_Wij_nx242), .A0 (nx2296), .A1 (RST)
          , .A2 (nx2288), .B0 (nx2076), .B1 (nx2856)) ;
    inv01 ix2295 (.Y (nx2296), .A (WindowDout_3__2__3)) ;
    oai32 L0_2_L1_2_Wij_ix253 (.Y (L0_2_L1_2_Wij_nx252), .A0 (nx2298), .A1 (RST)
          , .A2 (nx2288), .B0 (nx2078), .B1 (nx2856)) ;
    inv01 ix2297 (.Y (nx2298), .A (WindowDout_3__2__4)) ;
    oai32 L0_2_L1_2_Wij_ix263 (.Y (L0_2_L1_2_Wij_nx262), .A0 (nx2300), .A1 (RST)
          , .A2 (nx2288), .B0 (nx2080), .B1 (nx2856)) ;
    inv01 ix2299 (.Y (nx2300), .A (WindowDout_3__2__5)) ;
    oai32 L0_2_L1_2_Wij_ix273 (.Y (L0_2_L1_2_Wij_nx272), .A0 (nx2302), .A1 (RST)
          , .A2 (nx2304), .B0 (nx2082), .B1 (nx2856)) ;
    inv01 ix2301 (.Y (nx2302), .A (WindowDout_3__2__6)) ;
    inv01 ix2303 (.Y (nx2304), .A (L0_2_L1_2_Wij_nx333)) ;
    oai32 L0_2_L1_2_Wij_ix283 (.Y (L0_2_L1_2_Wij_nx282), .A0 (nx2306), .A1 (RST)
          , .A2 (nx2304), .B0 (nx2086), .B1 (nx2858)) ;
    inv01 ix2305 (.Y (nx2306), .A (WindowDout_3__2__7)) ;
    oai32 L0_2_L1_3_Fij_ix213 (.Y (L0_2_L1_3_Fij_nx212), .A0 (nx2308), .A1 (RST)
          , .A2 (nx2310), .B0 (nx2088), .B1 (nx2860)) ;
    inv01 ix2307 (.Y (nx2308), .A (FilterDout_3__3__0)) ;
    inv02 ix2309 (.Y (nx2310), .A (L0_2_L1_3_Fij_nx331)) ;
    oai32 L0_2_L1_3_Fij_ix223 (.Y (L0_2_L1_3_Fij_nx222), .A0 (nx2314), .A1 (RST)
          , .A2 (nx2310), .B0 (nx2094), .B1 (nx2860)) ;
    inv01 ix2313 (.Y (nx2314), .A (FilterDout_3__3__1)) ;
    oai32 L0_2_L1_3_Fij_ix233 (.Y (L0_2_L1_3_Fij_nx232), .A0 (nx2316), .A1 (RST)
          , .A2 (nx2310), .B0 (nx2096), .B1 (nx2860)) ;
    inv01 ix2315 (.Y (nx2316), .A (FilterDout_3__3__2)) ;
    oai32 L0_2_L1_3_Fij_ix243 (.Y (L0_2_L1_3_Fij_nx242), .A0 (nx2318), .A1 (RST)
          , .A2 (nx2310), .B0 (nx2098), .B1 (nx2860)) ;
    inv01 ix2317 (.Y (nx2318), .A (FilterDout_3__3__3)) ;
    oai32 L0_2_L1_3_Fij_ix253 (.Y (L0_2_L1_3_Fij_nx252), .A0 (nx2320), .A1 (RST)
          , .A2 (nx2310), .B0 (nx2100), .B1 (nx2860)) ;
    inv01 ix2319 (.Y (nx2320), .A (FilterDout_3__3__4)) ;
    oai32 L0_2_L1_3_Fij_ix263 (.Y (L0_2_L1_3_Fij_nx262), .A0 (nx2322), .A1 (RST)
          , .A2 (nx2310), .B0 (nx2102), .B1 (nx2860)) ;
    inv01 ix2321 (.Y (nx2322), .A (FilterDout_3__3__5)) ;
    oai32 L0_2_L1_3_Fij_ix273 (.Y (L0_2_L1_3_Fij_nx272), .A0 (nx2324), .A1 (RST)
          , .A2 (nx2326), .B0 (nx2104), .B1 (nx2860)) ;
    inv01 ix2323 (.Y (nx2324), .A (FilterDout_3__3__6)) ;
    inv01 ix2325 (.Y (nx2326), .A (L0_2_L1_3_Fij_nx333)) ;
    oai32 L0_2_L1_3_Fij_ix283 (.Y (L0_2_L1_3_Fij_nx282), .A0 (nx2328), .A1 (RST)
          , .A2 (nx2326), .B0 (nx2108), .B1 (nx2862)) ;
    inv01 ix2327 (.Y (nx2328), .A (FilterDout_3__3__7)) ;
    oai32 L0_2_L1_3_Wij_ix213 (.Y (L0_2_L1_3_Wij_nx212), .A0 (nx2330), .A1 (RST)
          , .A2 (nx2332), .B0 (nx2110), .B1 (nx2864)) ;
    inv01 ix2329 (.Y (nx2330), .A (WindowDout_3__3__0)) ;
    inv02 ix2331 (.Y (nx2332), .A (L0_2_L1_3_Wij_nx331)) ;
    oai32 L0_2_L1_3_Wij_ix223 (.Y (L0_2_L1_3_Wij_nx222), .A0 (nx2336), .A1 (RST)
          , .A2 (nx2332), .B0 (nx2116), .B1 (nx2864)) ;
    inv01 ix2335 (.Y (nx2336), .A (WindowDout_3__3__1)) ;
    oai32 L0_2_L1_3_Wij_ix233 (.Y (L0_2_L1_3_Wij_nx232), .A0 (nx2338), .A1 (RST)
          , .A2 (nx2332), .B0 (nx2118), .B1 (nx2864)) ;
    inv01 ix2337 (.Y (nx2338), .A (WindowDout_3__3__2)) ;
    oai32 L0_2_L1_3_Wij_ix243 (.Y (L0_2_L1_3_Wij_nx242), .A0 (nx2340), .A1 (RST)
          , .A2 (nx2332), .B0 (nx2120), .B1 (nx2864)) ;
    inv01 ix2339 (.Y (nx2340), .A (WindowDout_3__3__3)) ;
    oai32 L0_2_L1_3_Wij_ix253 (.Y (L0_2_L1_3_Wij_nx252), .A0 (nx2342), .A1 (RST)
          , .A2 (nx2332), .B0 (nx2122), .B1 (nx2864)) ;
    inv01 ix2341 (.Y (nx2342), .A (WindowDout_3__3__4)) ;
    oai32 L0_2_L1_3_Wij_ix263 (.Y (L0_2_L1_3_Wij_nx262), .A0 (nx2344), .A1 (RST)
          , .A2 (nx2332), .B0 (nx2124), .B1 (nx2864)) ;
    inv01 ix2343 (.Y (nx2344), .A (WindowDout_3__3__5)) ;
    oai32 L0_2_L1_3_Wij_ix273 (.Y (L0_2_L1_3_Wij_nx272), .A0 (nx2346), .A1 (RST)
          , .A2 (nx2348), .B0 (nx2126), .B1 (nx2864)) ;
    inv01 ix2345 (.Y (nx2346), .A (WindowDout_3__3__6)) ;
    inv01 ix2347 (.Y (nx2348), .A (L0_2_L1_3_Wij_nx333)) ;
    oai32 L0_2_L1_3_Wij_ix283 (.Y (L0_2_L1_3_Wij_nx282), .A0 (nx2350), .A1 (RST)
          , .A2 (nx2348), .B0 (nx2130), .B1 (nx2866)) ;
    inv01 ix2349 (.Y (nx2350), .A (WindowDout_3__3__7)) ;
    oai32 L0_2_L1_4_Fij_ix213 (.Y (L0_2_L1_4_Fij_nx212), .A0 (nx2352), .A1 (RST)
          , .A2 (nx2354), .B0 (nx2132), .B1 (nx2868)) ;
    inv01 ix2351 (.Y (nx2352), .A (FilterDout_3__4__0)) ;
    inv02 ix2353 (.Y (nx2354), .A (L0_2_L1_4_Fij_nx331)) ;
    oai32 L0_2_L1_4_Fij_ix223 (.Y (L0_2_L1_4_Fij_nx222), .A0 (nx2358), .A1 (RST)
          , .A2 (nx2354), .B0 (nx2138), .B1 (nx2868)) ;
    inv01 ix2357 (.Y (nx2358), .A (FilterDout_3__4__1)) ;
    oai32 L0_2_L1_4_Fij_ix233 (.Y (L0_2_L1_4_Fij_nx232), .A0 (nx2360), .A1 (RST)
          , .A2 (nx2354), .B0 (nx2140), .B1 (nx2868)) ;
    inv01 ix2359 (.Y (nx2360), .A (FilterDout_3__4__2)) ;
    oai32 L0_2_L1_4_Fij_ix243 (.Y (L0_2_L1_4_Fij_nx242), .A0 (nx2362), .A1 (RST)
          , .A2 (nx2354), .B0 (nx2142), .B1 (nx2868)) ;
    inv01 ix2361 (.Y (nx2362), .A (FilterDout_3__4__3)) ;
    oai32 L0_2_L1_4_Fij_ix253 (.Y (L0_2_L1_4_Fij_nx252), .A0 (nx2364), .A1 (RST)
          , .A2 (nx2354), .B0 (nx2144), .B1 (nx2868)) ;
    inv01 ix2363 (.Y (nx2364), .A (FilterDout_3__4__4)) ;
    oai32 L0_2_L1_4_Fij_ix263 (.Y (L0_2_L1_4_Fij_nx262), .A0 (nx2366), .A1 (RST)
          , .A2 (nx2354), .B0 (nx2146), .B1 (nx2868)) ;
    inv01 ix2365 (.Y (nx2366), .A (FilterDout_3__4__5)) ;
    oai32 L0_2_L1_4_Fij_ix273 (.Y (L0_2_L1_4_Fij_nx272), .A0 (nx2368), .A1 (RST)
          , .A2 (nx2370), .B0 (nx2148), .B1 (nx2868)) ;
    inv01 ix2367 (.Y (nx2368), .A (FilterDout_3__4__6)) ;
    inv01 ix2369 (.Y (nx2370), .A (L0_2_L1_4_Fij_nx333)) ;
    oai32 L0_2_L1_4_Fij_ix283 (.Y (L0_2_L1_4_Fij_nx282), .A0 (nx2372), .A1 (RST)
          , .A2 (nx2370), .B0 (nx2152), .B1 (nx2870)) ;
    inv01 ix2371 (.Y (nx2372), .A (FilterDout_3__4__7)) ;
    oai32 L0_2_L1_4_Wij_ix213 (.Y (L0_2_L1_4_Wij_nx212), .A0 (nx2374), .A1 (RST)
          , .A2 (nx2376), .B0 (nx2154), .B1 (nx2872)) ;
    inv01 ix2373 (.Y (nx2374), .A (WindowDout_3__4__0)) ;
    inv02 ix2375 (.Y (nx2376), .A (L0_2_L1_4_Wij_nx331)) ;
    oai32 L0_2_L1_4_Wij_ix223 (.Y (L0_2_L1_4_Wij_nx222), .A0 (nx2380), .A1 (RST)
          , .A2 (nx2376), .B0 (nx2160), .B1 (nx2872)) ;
    inv01 ix2379 (.Y (nx2380), .A (WindowDout_3__4__1)) ;
    oai32 L0_2_L1_4_Wij_ix233 (.Y (L0_2_L1_4_Wij_nx232), .A0 (nx2382), .A1 (RST)
          , .A2 (nx2376), .B0 (nx2162), .B1 (nx2872)) ;
    inv01 ix2381 (.Y (nx2382), .A (WindowDout_3__4__2)) ;
    oai32 L0_2_L1_4_Wij_ix243 (.Y (L0_2_L1_4_Wij_nx242), .A0 (nx2384), .A1 (RST)
          , .A2 (nx2376), .B0 (nx2164), .B1 (nx2872)) ;
    inv01 ix2383 (.Y (nx2384), .A (WindowDout_3__4__3)) ;
    oai32 L0_2_L1_4_Wij_ix253 (.Y (L0_2_L1_4_Wij_nx252), .A0 (nx2386), .A1 (RST)
          , .A2 (nx2376), .B0 (nx2166), .B1 (nx2872)) ;
    inv01 ix2385 (.Y (nx2386), .A (WindowDout_3__4__4)) ;
    oai32 L0_2_L1_4_Wij_ix263 (.Y (L0_2_L1_4_Wij_nx262), .A0 (nx2388), .A1 (RST)
          , .A2 (nx2376), .B0 (nx2168), .B1 (nx2872)) ;
    inv01 ix2387 (.Y (nx2388), .A (WindowDout_3__4__5)) ;
    oai32 L0_2_L1_4_Wij_ix273 (.Y (L0_2_L1_4_Wij_nx272), .A0 (nx2390), .A1 (RST)
          , .A2 (nx2392), .B0 (nx2170), .B1 (nx2872)) ;
    inv01 ix2389 (.Y (nx2390), .A (WindowDout_3__4__6)) ;
    inv01 ix2391 (.Y (nx2392), .A (L0_2_L1_4_Wij_nx333)) ;
    oai32 L0_2_L1_4_Wij_ix283 (.Y (L0_2_L1_4_Wij_nx282), .A0 (nx2394), .A1 (RST)
          , .A2 (nx2392), .B0 (nx2174), .B1 (nx2874)) ;
    inv01 ix2393 (.Y (nx2394), .A (WindowDout_3__4__7)) ;
    oai32 L0_3_L1_0_Fij_ix213 (.Y (L0_3_L1_0_Fij_nx212), .A0 (nx2396), .A1 (RST)
          , .A2 (nx2398), .B0 (nx2176), .B1 (nx2876)) ;
    inv01 ix2395 (.Y (nx2396), .A (FilterDout_4__0__0)) ;
    inv02 ix2397 (.Y (nx2398), .A (L0_3_L1_0_Fij_nx331)) ;
    oai32 L0_3_L1_0_Fij_ix223 (.Y (L0_3_L1_0_Fij_nx222), .A0 (nx2402), .A1 (RST)
          , .A2 (nx2398), .B0 (nx2182), .B1 (nx2876)) ;
    inv01 ix2401 (.Y (nx2402), .A (FilterDout_4__0__1)) ;
    oai32 L0_3_L1_0_Fij_ix233 (.Y (L0_3_L1_0_Fij_nx232), .A0 (nx2404), .A1 (RST)
          , .A2 (nx2398), .B0 (nx2184), .B1 (nx2876)) ;
    inv01 ix2403 (.Y (nx2404), .A (FilterDout_4__0__2)) ;
    oai32 L0_3_L1_0_Fij_ix243 (.Y (L0_3_L1_0_Fij_nx242), .A0 (nx2406), .A1 (RST)
          , .A2 (nx2398), .B0 (nx2186), .B1 (nx2876)) ;
    inv01 ix2405 (.Y (nx2406), .A (FilterDout_4__0__3)) ;
    oai32 L0_3_L1_0_Fij_ix253 (.Y (L0_3_L1_0_Fij_nx252), .A0 (nx2408), .A1 (RST)
          , .A2 (nx2398), .B0 (nx2188), .B1 (nx2876)) ;
    inv01 ix2407 (.Y (nx2408), .A (FilterDout_4__0__4)) ;
    oai32 L0_3_L1_0_Fij_ix263 (.Y (L0_3_L1_0_Fij_nx262), .A0 (nx2410), .A1 (RST)
          , .A2 (nx2398), .B0 (nx2190), .B1 (nx2876)) ;
    inv01 ix2409 (.Y (nx2410), .A (FilterDout_4__0__5)) ;
    oai32 L0_3_L1_0_Fij_ix273 (.Y (L0_3_L1_0_Fij_nx272), .A0 (nx2412), .A1 (RST)
          , .A2 (nx2414), .B0 (nx2192), .B1 (nx2876)) ;
    inv01 ix2411 (.Y (nx2412), .A (FilterDout_4__0__6)) ;
    inv01 ix2413 (.Y (nx2414), .A (L0_3_L1_0_Fij_nx333)) ;
    oai32 L0_3_L1_0_Fij_ix283 (.Y (L0_3_L1_0_Fij_nx282), .A0 (nx2416), .A1 (RST)
          , .A2 (nx2414), .B0 (nx2196), .B1 (nx2878)) ;
    inv01 ix2415 (.Y (nx2416), .A (FilterDout_4__0__7)) ;
    oai32 L0_3_L1_0_Wij_ix213 (.Y (L0_3_L1_0_Wij_nx212), .A0 (nx2418), .A1 (RST)
          , .A2 (nx2420), .B0 (nx2198), .B1 (nx2880)) ;
    inv01 ix2417 (.Y (nx2418), .A (WindowDout_4__0__0)) ;
    inv02 ix2419 (.Y (nx2420), .A (L0_3_L1_0_Wij_nx331)) ;
    oai32 L0_3_L1_0_Wij_ix223 (.Y (L0_3_L1_0_Wij_nx222), .A0 (nx2424), .A1 (RST)
          , .A2 (nx2420), .B0 (nx2204), .B1 (nx2880)) ;
    inv01 ix2423 (.Y (nx2424), .A (WindowDout_4__0__1)) ;
    oai32 L0_3_L1_0_Wij_ix233 (.Y (L0_3_L1_0_Wij_nx232), .A0 (nx2426), .A1 (RST)
          , .A2 (nx2420), .B0 (nx2206), .B1 (nx2880)) ;
    inv01 ix2425 (.Y (nx2426), .A (WindowDout_4__0__2)) ;
    oai32 L0_3_L1_0_Wij_ix243 (.Y (L0_3_L1_0_Wij_nx242), .A0 (nx2428), .A1 (RST)
          , .A2 (nx2420), .B0 (nx2208), .B1 (nx2880)) ;
    inv01 ix2427 (.Y (nx2428), .A (WindowDout_4__0__3)) ;
    oai32 L0_3_L1_0_Wij_ix253 (.Y (L0_3_L1_0_Wij_nx252), .A0 (nx2430), .A1 (RST)
          , .A2 (nx2420), .B0 (nx2210), .B1 (nx2880)) ;
    inv01 ix2429 (.Y (nx2430), .A (WindowDout_4__0__4)) ;
    oai32 L0_3_L1_0_Wij_ix263 (.Y (L0_3_L1_0_Wij_nx262), .A0 (nx2432), .A1 (RST)
          , .A2 (nx2420), .B0 (nx2212), .B1 (nx2880)) ;
    inv01 ix2431 (.Y (nx2432), .A (WindowDout_4__0__5)) ;
    oai32 L0_3_L1_0_Wij_ix273 (.Y (L0_3_L1_0_Wij_nx272), .A0 (nx2434), .A1 (RST)
          , .A2 (nx2436), .B0 (nx2214), .B1 (nx2880)) ;
    inv01 ix2433 (.Y (nx2434), .A (WindowDout_4__0__6)) ;
    inv01 ix2435 (.Y (nx2436), .A (L0_3_L1_0_Wij_nx333)) ;
    oai32 L0_3_L1_0_Wij_ix283 (.Y (L0_3_L1_0_Wij_nx282), .A0 (nx2438), .A1 (RST)
          , .A2 (nx2436), .B0 (nx2218), .B1 (nx2882)) ;
    inv01 ix2437 (.Y (nx2438), .A (WindowDout_4__0__7)) ;
    oai32 L0_3_L1_1_Fij_ix213 (.Y (L0_3_L1_1_Fij_nx212), .A0 (nx2440), .A1 (RST)
          , .A2 (nx2442), .B0 (nx2220), .B1 (nx2884)) ;
    inv01 ix2439 (.Y (nx2440), .A (FilterDout_4__1__0)) ;
    inv02 ix2441 (.Y (nx2442), .A (L0_3_L1_1_Fij_nx331)) ;
    oai32 L0_3_L1_1_Fij_ix223 (.Y (L0_3_L1_1_Fij_nx222), .A0 (nx2446), .A1 (RST)
          , .A2 (nx2442), .B0 (nx2226), .B1 (nx2884)) ;
    inv01 ix2445 (.Y (nx2446), .A (FilterDout_4__1__1)) ;
    oai32 L0_3_L1_1_Fij_ix233 (.Y (L0_3_L1_1_Fij_nx232), .A0 (nx2448), .A1 (RST)
          , .A2 (nx2442), .B0 (nx2228), .B1 (nx2884)) ;
    inv01 ix2447 (.Y (nx2448), .A (FilterDout_4__1__2)) ;
    oai32 L0_3_L1_1_Fij_ix243 (.Y (L0_3_L1_1_Fij_nx242), .A0 (nx2450), .A1 (RST)
          , .A2 (nx2442), .B0 (nx2230), .B1 (nx2884)) ;
    inv01 ix2449 (.Y (nx2450), .A (FilterDout_4__1__3)) ;
    oai32 L0_3_L1_1_Fij_ix253 (.Y (L0_3_L1_1_Fij_nx252), .A0 (nx2452), .A1 (RST)
          , .A2 (nx2442), .B0 (nx2232), .B1 (nx2884)) ;
    inv01 ix2451 (.Y (nx2452), .A (FilterDout_4__1__4)) ;
    oai32 L0_3_L1_1_Fij_ix263 (.Y (L0_3_L1_1_Fij_nx262), .A0 (nx2454), .A1 (RST)
          , .A2 (nx2442), .B0 (nx2234), .B1 (nx2884)) ;
    inv01 ix2453 (.Y (nx2454), .A (FilterDout_4__1__5)) ;
    oai32 L0_3_L1_1_Fij_ix273 (.Y (L0_3_L1_1_Fij_nx272), .A0 (nx2456), .A1 (RST)
          , .A2 (nx2458), .B0 (nx2236), .B1 (nx2884)) ;
    inv01 ix2455 (.Y (nx2456), .A (FilterDout_4__1__6)) ;
    inv01 ix2457 (.Y (nx2458), .A (L0_3_L1_1_Fij_nx333)) ;
    oai32 L0_3_L1_1_Fij_ix283 (.Y (L0_3_L1_1_Fij_nx282), .A0 (nx2460), .A1 (RST)
          , .A2 (nx2458), .B0 (nx2240), .B1 (nx2886)) ;
    inv01 ix2459 (.Y (nx2460), .A (FilterDout_4__1__7)) ;
    oai32 L0_3_L1_1_Wij_ix213 (.Y (L0_3_L1_1_Wij_nx212), .A0 (nx2462), .A1 (RST)
          , .A2 (nx2464), .B0 (nx2242), .B1 (nx2888)) ;
    inv01 ix2461 (.Y (nx2462), .A (WindowDout_4__1__0)) ;
    inv02 ix2463 (.Y (nx2464), .A (L0_3_L1_1_Wij_nx331)) ;
    oai32 L0_3_L1_1_Wij_ix223 (.Y (L0_3_L1_1_Wij_nx222), .A0 (nx2468), .A1 (RST)
          , .A2 (nx2464), .B0 (nx2248), .B1 (nx2888)) ;
    inv01 ix2467 (.Y (nx2468), .A (WindowDout_4__1__1)) ;
    oai32 L0_3_L1_1_Wij_ix233 (.Y (L0_3_L1_1_Wij_nx232), .A0 (nx2470), .A1 (RST)
          , .A2 (nx2464), .B0 (nx2250), .B1 (nx2888)) ;
    inv01 ix2469 (.Y (nx2470), .A (WindowDout_4__1__2)) ;
    oai32 L0_3_L1_1_Wij_ix243 (.Y (L0_3_L1_1_Wij_nx242), .A0 (nx2472), .A1 (RST)
          , .A2 (nx2464), .B0 (nx2252), .B1 (nx2888)) ;
    inv01 ix2471 (.Y (nx2472), .A (WindowDout_4__1__3)) ;
    oai32 L0_3_L1_1_Wij_ix253 (.Y (L0_3_L1_1_Wij_nx252), .A0 (nx2474), .A1 (RST)
          , .A2 (nx2464), .B0 (nx2254), .B1 (nx2888)) ;
    inv01 ix2473 (.Y (nx2474), .A (WindowDout_4__1__4)) ;
    oai32 L0_3_L1_1_Wij_ix263 (.Y (L0_3_L1_1_Wij_nx262), .A0 (nx2476), .A1 (RST)
          , .A2 (nx2464), .B0 (nx2256), .B1 (nx2888)) ;
    inv01 ix2475 (.Y (nx2476), .A (WindowDout_4__1__5)) ;
    oai32 L0_3_L1_1_Wij_ix273 (.Y (L0_3_L1_1_Wij_nx272), .A0 (nx2478), .A1 (RST)
          , .A2 (nx2480), .B0 (nx2258), .B1 (nx2888)) ;
    inv01 ix2477 (.Y (nx2478), .A (WindowDout_4__1__6)) ;
    inv01 ix2479 (.Y (nx2480), .A (L0_3_L1_1_Wij_nx333)) ;
    oai32 L0_3_L1_1_Wij_ix283 (.Y (L0_3_L1_1_Wij_nx282), .A0 (nx2482), .A1 (RST)
          , .A2 (nx2480), .B0 (nx2262), .B1 (nx2890)) ;
    inv01 ix2481 (.Y (nx2482), .A (WindowDout_4__1__7)) ;
    oai32 L0_3_L1_2_Fij_ix213 (.Y (L0_3_L1_2_Fij_nx212), .A0 (nx2484), .A1 (RST)
          , .A2 (nx2486), .B0 (nx2264), .B1 (nx2892)) ;
    inv01 ix2483 (.Y (nx2484), .A (FilterDout_4__2__0)) ;
    inv02 ix2485 (.Y (nx2486), .A (L0_3_L1_2_Fij_nx331)) ;
    oai32 L0_3_L1_2_Fij_ix223 (.Y (L0_3_L1_2_Fij_nx222), .A0 (nx2490), .A1 (RST)
          , .A2 (nx2486), .B0 (nx2270), .B1 (nx2892)) ;
    inv01 ix2489 (.Y (nx2490), .A (FilterDout_4__2__1)) ;
    oai32 L0_3_L1_2_Fij_ix233 (.Y (L0_3_L1_2_Fij_nx232), .A0 (nx2492), .A1 (RST)
          , .A2 (nx2486), .B0 (nx2272), .B1 (nx2892)) ;
    inv01 ix2491 (.Y (nx2492), .A (FilterDout_4__2__2)) ;
    oai32 L0_3_L1_2_Fij_ix243 (.Y (L0_3_L1_2_Fij_nx242), .A0 (nx2494), .A1 (RST)
          , .A2 (nx2486), .B0 (nx2274), .B1 (nx2892)) ;
    inv01 ix2493 (.Y (nx2494), .A (FilterDout_4__2__3)) ;
    oai32 L0_3_L1_2_Fij_ix253 (.Y (L0_3_L1_2_Fij_nx252), .A0 (nx2496), .A1 (RST)
          , .A2 (nx2486), .B0 (nx2276), .B1 (nx2892)) ;
    inv01 ix2495 (.Y (nx2496), .A (FilterDout_4__2__4)) ;
    oai32 L0_3_L1_2_Fij_ix263 (.Y (L0_3_L1_2_Fij_nx262), .A0 (nx2498), .A1 (RST)
          , .A2 (nx2486), .B0 (nx2278), .B1 (nx2892)) ;
    inv01 ix2497 (.Y (nx2498), .A (FilterDout_4__2__5)) ;
    oai32 L0_3_L1_2_Fij_ix273 (.Y (L0_3_L1_2_Fij_nx272), .A0 (nx2500), .A1 (RST)
          , .A2 (nx2502), .B0 (nx2280), .B1 (nx2892)) ;
    inv01 ix2499 (.Y (nx2500), .A (FilterDout_4__2__6)) ;
    inv01 ix2501 (.Y (nx2502), .A (L0_3_L1_2_Fij_nx333)) ;
    oai32 L0_3_L1_2_Fij_ix283 (.Y (L0_3_L1_2_Fij_nx282), .A0 (nx2504), .A1 (RST)
          , .A2 (nx2502), .B0 (nx2284), .B1 (nx2894)) ;
    inv01 ix2503 (.Y (nx2504), .A (FilterDout_4__2__7)) ;
    oai32 L0_3_L1_2_Wij_ix213 (.Y (L0_3_L1_2_Wij_nx212), .A0 (nx2506), .A1 (RST)
          , .A2 (nx2508), .B0 (nx2286), .B1 (nx2896)) ;
    inv01 ix2505 (.Y (nx2506), .A (WindowDout_4__2__0)) ;
    inv02 ix2507 (.Y (nx2508), .A (L0_3_L1_2_Wij_nx331)) ;
    oai32 L0_3_L1_2_Wij_ix223 (.Y (L0_3_L1_2_Wij_nx222), .A0 (nx2512), .A1 (RST)
          , .A2 (nx2508), .B0 (nx2292), .B1 (nx2896)) ;
    inv01 ix2511 (.Y (nx2512), .A (WindowDout_4__2__1)) ;
    oai32 L0_3_L1_2_Wij_ix233 (.Y (L0_3_L1_2_Wij_nx232), .A0 (nx2514), .A1 (RST)
          , .A2 (nx2508), .B0 (nx2294), .B1 (nx2896)) ;
    inv01 ix2513 (.Y (nx2514), .A (WindowDout_4__2__2)) ;
    oai32 L0_3_L1_2_Wij_ix243 (.Y (L0_3_L1_2_Wij_nx242), .A0 (nx2516), .A1 (RST)
          , .A2 (nx2508), .B0 (nx2296), .B1 (nx2896)) ;
    inv01 ix2515 (.Y (nx2516), .A (WindowDout_4__2__3)) ;
    oai32 L0_3_L1_2_Wij_ix253 (.Y (L0_3_L1_2_Wij_nx252), .A0 (nx2518), .A1 (RST)
          , .A2 (nx2508), .B0 (nx2298), .B1 (nx2896)) ;
    inv01 ix2517 (.Y (nx2518), .A (WindowDout_4__2__4)) ;
    oai32 L0_3_L1_2_Wij_ix263 (.Y (L0_3_L1_2_Wij_nx262), .A0 (nx2520), .A1 (RST)
          , .A2 (nx2508), .B0 (nx2300), .B1 (nx2896)) ;
    inv01 ix2519 (.Y (nx2520), .A (WindowDout_4__2__5)) ;
    oai32 L0_3_L1_2_Wij_ix273 (.Y (L0_3_L1_2_Wij_nx272), .A0 (nx2522), .A1 (RST)
          , .A2 (nx2524), .B0 (nx2302), .B1 (nx2896)) ;
    inv01 ix2521 (.Y (nx2522), .A (WindowDout_4__2__6)) ;
    inv01 ix2523 (.Y (nx2524), .A (L0_3_L1_2_Wij_nx333)) ;
    oai32 L0_3_L1_2_Wij_ix283 (.Y (L0_3_L1_2_Wij_nx282), .A0 (nx2526), .A1 (RST)
          , .A2 (nx2524), .B0 (nx2306), .B1 (nx2898)) ;
    inv01 ix2525 (.Y (nx2526), .A (WindowDout_4__2__7)) ;
    oai32 L0_3_L1_3_Fij_ix213 (.Y (L0_3_L1_3_Fij_nx212), .A0 (nx2528), .A1 (RST)
          , .A2 (nx2530), .B0 (nx2308), .B1 (nx2900)) ;
    inv01 ix2527 (.Y (nx2528), .A (FilterDout_4__3__0)) ;
    inv02 ix2529 (.Y (nx2530), .A (L0_3_L1_3_Fij_nx331)) ;
    oai32 L0_3_L1_3_Fij_ix223 (.Y (L0_3_L1_3_Fij_nx222), .A0 (nx2534), .A1 (RST)
          , .A2 (nx2530), .B0 (nx2314), .B1 (nx2900)) ;
    inv01 ix2533 (.Y (nx2534), .A (FilterDout_4__3__1)) ;
    oai32 L0_3_L1_3_Fij_ix233 (.Y (L0_3_L1_3_Fij_nx232), .A0 (nx2536), .A1 (RST)
          , .A2 (nx2530), .B0 (nx2316), .B1 (nx2900)) ;
    inv01 ix2535 (.Y (nx2536), .A (FilterDout_4__3__2)) ;
    oai32 L0_3_L1_3_Fij_ix243 (.Y (L0_3_L1_3_Fij_nx242), .A0 (nx2538), .A1 (RST)
          , .A2 (nx2530), .B0 (nx2318), .B1 (nx2900)) ;
    inv01 ix2537 (.Y (nx2538), .A (FilterDout_4__3__3)) ;
    oai32 L0_3_L1_3_Fij_ix253 (.Y (L0_3_L1_3_Fij_nx252), .A0 (nx2540), .A1 (RST)
          , .A2 (nx2530), .B0 (nx2320), .B1 (nx2900)) ;
    inv01 ix2539 (.Y (nx2540), .A (FilterDout_4__3__4)) ;
    oai32 L0_3_L1_3_Fij_ix263 (.Y (L0_3_L1_3_Fij_nx262), .A0 (nx2542), .A1 (RST)
          , .A2 (nx2530), .B0 (nx2322), .B1 (nx2900)) ;
    inv01 ix2541 (.Y (nx2542), .A (FilterDout_4__3__5)) ;
    oai32 L0_3_L1_3_Fij_ix273 (.Y (L0_3_L1_3_Fij_nx272), .A0 (nx2544), .A1 (RST)
          , .A2 (nx2546), .B0 (nx2324), .B1 (nx2900)) ;
    inv01 ix2543 (.Y (nx2544), .A (FilterDout_4__3__6)) ;
    inv01 ix2545 (.Y (nx2546), .A (L0_3_L1_3_Fij_nx333)) ;
    oai32 L0_3_L1_3_Fij_ix283 (.Y (L0_3_L1_3_Fij_nx282), .A0 (nx2548), .A1 (RST)
          , .A2 (nx2546), .B0 (nx2328), .B1 (nx2902)) ;
    inv01 ix2547 (.Y (nx2548), .A (FilterDout_4__3__7)) ;
    oai32 L0_3_L1_3_Wij_ix213 (.Y (L0_3_L1_3_Wij_nx212), .A0 (nx2550), .A1 (RST)
          , .A2 (nx2552), .B0 (nx2330), .B1 (nx2904)) ;
    inv01 ix2549 (.Y (nx2550), .A (WindowDout_4__3__0)) ;
    inv02 ix2551 (.Y (nx2552), .A (L0_3_L1_3_Wij_nx331)) ;
    oai32 L0_3_L1_3_Wij_ix223 (.Y (L0_3_L1_3_Wij_nx222), .A0 (nx2556), .A1 (RST)
          , .A2 (nx2552), .B0 (nx2336), .B1 (nx2904)) ;
    inv01 ix2555 (.Y (nx2556), .A (WindowDout_4__3__1)) ;
    oai32 L0_3_L1_3_Wij_ix233 (.Y (L0_3_L1_3_Wij_nx232), .A0 (nx2558), .A1 (RST)
          , .A2 (nx2552), .B0 (nx2338), .B1 (nx2904)) ;
    inv01 ix2557 (.Y (nx2558), .A (WindowDout_4__3__2)) ;
    oai32 L0_3_L1_3_Wij_ix243 (.Y (L0_3_L1_3_Wij_nx242), .A0 (nx2560), .A1 (RST)
          , .A2 (nx2552), .B0 (nx2340), .B1 (nx2904)) ;
    inv01 ix2559 (.Y (nx2560), .A (WindowDout_4__3__3)) ;
    oai32 L0_3_L1_3_Wij_ix253 (.Y (L0_3_L1_3_Wij_nx252), .A0 (nx2562), .A1 (RST)
          , .A2 (nx2552), .B0 (nx2342), .B1 (nx2904)) ;
    inv01 ix2561 (.Y (nx2562), .A (WindowDout_4__3__4)) ;
    oai32 L0_3_L1_3_Wij_ix263 (.Y (L0_3_L1_3_Wij_nx262), .A0 (nx2564), .A1 (RST)
          , .A2 (nx2552), .B0 (nx2344), .B1 (nx2904)) ;
    inv01 ix2563 (.Y (nx2564), .A (WindowDout_4__3__5)) ;
    oai32 L0_3_L1_3_Wij_ix273 (.Y (L0_3_L1_3_Wij_nx272), .A0 (nx2566), .A1 (RST)
          , .A2 (nx2568), .B0 (nx2346), .B1 (nx2904)) ;
    inv01 ix2565 (.Y (nx2566), .A (WindowDout_4__3__6)) ;
    inv01 ix2567 (.Y (nx2568), .A (L0_3_L1_3_Wij_nx333)) ;
    oai32 L0_3_L1_3_Wij_ix283 (.Y (L0_3_L1_3_Wij_nx282), .A0 (nx2570), .A1 (RST)
          , .A2 (nx2568), .B0 (nx2350), .B1 (nx2906)) ;
    inv01 ix2569 (.Y (nx2570), .A (WindowDout_4__3__7)) ;
    oai32 L0_3_L1_4_Fij_ix213 (.Y (L0_3_L1_4_Fij_nx212), .A0 (nx2572), .A1 (RST)
          , .A2 (nx2574), .B0 (nx2352), .B1 (nx2908)) ;
    inv01 ix2571 (.Y (nx2572), .A (FilterDout_4__4__0)) ;
    inv02 ix2573 (.Y (nx2574), .A (L0_3_L1_4_Fij_nx331)) ;
    oai32 L0_3_L1_4_Fij_ix223 (.Y (L0_3_L1_4_Fij_nx222), .A0 (nx2578), .A1 (RST)
          , .A2 (nx2574), .B0 (nx2358), .B1 (nx2908)) ;
    inv01 ix2577 (.Y (nx2578), .A (FilterDout_4__4__1)) ;
    oai32 L0_3_L1_4_Fij_ix233 (.Y (L0_3_L1_4_Fij_nx232), .A0 (nx2580), .A1 (RST)
          , .A2 (nx2574), .B0 (nx2360), .B1 (nx2908)) ;
    inv01 ix2579 (.Y (nx2580), .A (FilterDout_4__4__2)) ;
    oai32 L0_3_L1_4_Fij_ix243 (.Y (L0_3_L1_4_Fij_nx242), .A0 (nx2582), .A1 (RST)
          , .A2 (nx2574), .B0 (nx2362), .B1 (nx2908)) ;
    inv01 ix2581 (.Y (nx2582), .A (FilterDout_4__4__3)) ;
    oai32 L0_3_L1_4_Fij_ix253 (.Y (L0_3_L1_4_Fij_nx252), .A0 (nx2584), .A1 (RST)
          , .A2 (nx2574), .B0 (nx2364), .B1 (nx2908)) ;
    inv01 ix2583 (.Y (nx2584), .A (FilterDout_4__4__4)) ;
    oai32 L0_3_L1_4_Fij_ix263 (.Y (L0_3_L1_4_Fij_nx262), .A0 (nx2586), .A1 (RST)
          , .A2 (nx2574), .B0 (nx2366), .B1 (nx2908)) ;
    inv01 ix2585 (.Y (nx2586), .A (FilterDout_4__4__5)) ;
    oai32 L0_3_L1_4_Fij_ix273 (.Y (L0_3_L1_4_Fij_nx272), .A0 (nx2588), .A1 (RST)
          , .A2 (nx2590), .B0 (nx2368), .B1 (nx2908)) ;
    inv01 ix2587 (.Y (nx2588), .A (FilterDout_4__4__6)) ;
    inv01 ix2589 (.Y (nx2590), .A (L0_3_L1_4_Fij_nx333)) ;
    oai32 L0_3_L1_4_Fij_ix283 (.Y (L0_3_L1_4_Fij_nx282), .A0 (nx2592), .A1 (RST)
          , .A2 (nx2590), .B0 (nx2372), .B1 (nx2910)) ;
    inv01 ix2591 (.Y (nx2592), .A (FilterDout_4__4__7)) ;
    oai32 L0_3_L1_4_Wij_ix213 (.Y (L0_3_L1_4_Wij_nx212), .A0 (nx2594), .A1 (RST)
          , .A2 (nx2596), .B0 (nx2374), .B1 (nx2912)) ;
    inv01 ix2593 (.Y (nx2594), .A (WindowDout_4__4__0)) ;
    inv02 ix2595 (.Y (nx2596), .A (L0_3_L1_4_Wij_nx331)) ;
    oai32 L0_3_L1_4_Wij_ix223 (.Y (L0_3_L1_4_Wij_nx222), .A0 (nx2600), .A1 (RST)
          , .A2 (nx2596), .B0 (nx2380), .B1 (nx2912)) ;
    inv01 ix2599 (.Y (nx2600), .A (WindowDout_4__4__1)) ;
    oai32 L0_3_L1_4_Wij_ix233 (.Y (L0_3_L1_4_Wij_nx232), .A0 (nx2602), .A1 (RST)
          , .A2 (nx2596), .B0 (nx2382), .B1 (nx2912)) ;
    inv01 ix2601 (.Y (nx2602), .A (WindowDout_4__4__2)) ;
    oai32 L0_3_L1_4_Wij_ix243 (.Y (L0_3_L1_4_Wij_nx242), .A0 (nx2604), .A1 (RST)
          , .A2 (nx2596), .B0 (nx2384), .B1 (nx2912)) ;
    inv01 ix2603 (.Y (nx2604), .A (WindowDout_4__4__3)) ;
    oai32 L0_3_L1_4_Wij_ix253 (.Y (L0_3_L1_4_Wij_nx252), .A0 (nx2606), .A1 (RST)
          , .A2 (nx2596), .B0 (nx2386), .B1 (nx2912)) ;
    inv01 ix2605 (.Y (nx2606), .A (WindowDout_4__4__4)) ;
    oai32 L0_3_L1_4_Wij_ix263 (.Y (L0_3_L1_4_Wij_nx262), .A0 (nx2608), .A1 (RST)
          , .A2 (nx2596), .B0 (nx2388), .B1 (nx2912)) ;
    inv01 ix2607 (.Y (nx2608), .A (WindowDout_4__4__5)) ;
    oai32 L0_3_L1_4_Wij_ix273 (.Y (L0_3_L1_4_Wij_nx272), .A0 (nx2610), .A1 (RST)
          , .A2 (nx2612), .B0 (nx2390), .B1 (nx2912)) ;
    inv01 ix2609 (.Y (nx2610), .A (WindowDout_4__4__6)) ;
    inv01 ix2611 (.Y (nx2612), .A (L0_3_L1_4_Wij_nx333)) ;
    oai32 L0_3_L1_4_Wij_ix283 (.Y (L0_3_L1_4_Wij_nx282), .A0 (nx2614), .A1 (RST)
          , .A2 (nx2612), .B0 (nx2394), .B1 (nx2914)) ;
    inv01 ix2613 (.Y (nx2614), .A (WindowDout_4__4__7)) ;
    oai32 L0_4_L1_0_Fij_ix213 (.Y (L0_4_L1_0_Fij_nx212), .A0 (nx2616), .A1 (RST)
          , .A2 (nx2618), .B0 (nx2396), .B1 (nx2916)) ;
    inv01 ix2615 (.Y (nx2616), .A (Din[0])) ;
    inv02 ix2617 (.Y (nx2618), .A (L0_4_L1_0_Fij_nx331)) ;
    oai32 L0_4_L1_0_Fij_ix223 (.Y (L0_4_L1_0_Fij_nx222), .A0 (nx2622), .A1 (RST)
          , .A2 (nx2618), .B0 (nx2402), .B1 (nx2916)) ;
    inv01 ix2621 (.Y (nx2622), .A (Din[1])) ;
    oai32 L0_4_L1_0_Fij_ix233 (.Y (L0_4_L1_0_Fij_nx232), .A0 (nx2624), .A1 (RST)
          , .A2 (nx2618), .B0 (nx2404), .B1 (nx2916)) ;
    inv01 ix2623 (.Y (nx2624), .A (Din[2])) ;
    oai32 L0_4_L1_0_Fij_ix243 (.Y (L0_4_L1_0_Fij_nx242), .A0 (nx2626), .A1 (RST)
          , .A2 (nx2618), .B0 (nx2406), .B1 (nx2916)) ;
    inv01 ix2625 (.Y (nx2626), .A (Din[3])) ;
    oai32 L0_4_L1_0_Fij_ix253 (.Y (L0_4_L1_0_Fij_nx252), .A0 (nx2628), .A1 (RST)
          , .A2 (nx2618), .B0 (nx2408), .B1 (nx2916)) ;
    inv01 ix2627 (.Y (nx2628), .A (Din[4])) ;
    oai32 L0_4_L1_0_Fij_ix263 (.Y (L0_4_L1_0_Fij_nx262), .A0 (nx2630), .A1 (RST)
          , .A2 (nx2618), .B0 (nx2410), .B1 (nx2916)) ;
    inv01 ix2629 (.Y (nx2630), .A (Din[5])) ;
    oai32 L0_4_L1_0_Fij_ix273 (.Y (L0_4_L1_0_Fij_nx272), .A0 (nx2632), .A1 (RST)
          , .A2 (nx2634), .B0 (nx2412), .B1 (nx2916)) ;
    inv01 ix2631 (.Y (nx2632), .A (Din[6])) ;
    inv01 ix2633 (.Y (nx2634), .A (L0_4_L1_0_Fij_nx333)) ;
    oai32 L0_4_L1_0_Fij_ix283 (.Y (L0_4_L1_0_Fij_nx282), .A0 (nx2636), .A1 (RST)
          , .A2 (nx2634), .B0 (nx2416), .B1 (nx2918)) ;
    inv01 ix2635 (.Y (nx2636), .A (Din[7])) ;
    oai32 L0_4_L1_0_Wij_ix213 (.Y (L0_4_L1_0_Wij_nx212), .A0 (nx2616), .A1 (RST)
          , .A2 (nx2638), .B0 (nx2418), .B1 (nx2920)) ;
    inv02 ix2637 (.Y (nx2638), .A (L0_4_L1_0_Wij_nx331)) ;
    oai32 L0_4_L1_0_Wij_ix223 (.Y (L0_4_L1_0_Wij_nx222), .A0 (nx2622), .A1 (RST)
          , .A2 (nx2638), .B0 (nx2424), .B1 (nx2920)) ;
    oai32 L0_4_L1_0_Wij_ix233 (.Y (L0_4_L1_0_Wij_nx232), .A0 (nx2624), .A1 (RST)
          , .A2 (nx2638), .B0 (nx2426), .B1 (nx2920)) ;
    oai32 L0_4_L1_0_Wij_ix243 (.Y (L0_4_L1_0_Wij_nx242), .A0 (nx2626), .A1 (RST)
          , .A2 (nx2638), .B0 (nx2428), .B1 (nx2920)) ;
    oai32 L0_4_L1_0_Wij_ix253 (.Y (L0_4_L1_0_Wij_nx252), .A0 (nx2628), .A1 (RST)
          , .A2 (nx2638), .B0 (nx2430), .B1 (nx2920)) ;
    oai32 L0_4_L1_0_Wij_ix263 (.Y (L0_4_L1_0_Wij_nx262), .A0 (nx2630), .A1 (RST)
          , .A2 (nx2638), .B0 (nx2432), .B1 (nx2920)) ;
    oai32 L0_4_L1_0_Wij_ix273 (.Y (L0_4_L1_0_Wij_nx272), .A0 (nx2632), .A1 (RST)
          , .A2 (nx2642), .B0 (nx2434), .B1 (nx2920)) ;
    inv01 ix2641 (.Y (nx2642), .A (L0_4_L1_0_Wij_nx333)) ;
    oai32 L0_4_L1_0_Wij_ix283 (.Y (L0_4_L1_0_Wij_nx282), .A0 (nx2636), .A1 (RST)
          , .A2 (nx2642), .B0 (nx2438), .B1 (nx2922)) ;
    oai32 L0_4_L1_1_Fij_ix213 (.Y (L0_4_L1_1_Fij_nx212), .A0 (nx2644), .A1 (RST)
          , .A2 (nx2646), .B0 (nx2440), .B1 (nx2924)) ;
    inv01 ix2643 (.Y (nx2644), .A (Din[8])) ;
    inv02 ix2645 (.Y (nx2646), .A (L0_4_L1_1_Fij_nx331)) ;
    oai32 L0_4_L1_1_Fij_ix223 (.Y (L0_4_L1_1_Fij_nx222), .A0 (nx2650), .A1 (RST)
          , .A2 (nx2646), .B0 (nx2446), .B1 (nx2924)) ;
    inv01 ix2649 (.Y (nx2650), .A (Din[9])) ;
    oai32 L0_4_L1_1_Fij_ix233 (.Y (L0_4_L1_1_Fij_nx232), .A0 (nx2652), .A1 (RST)
          , .A2 (nx2646), .B0 (nx2448), .B1 (nx2924)) ;
    inv01 ix2651 (.Y (nx2652), .A (Din[10])) ;
    oai32 L0_4_L1_1_Fij_ix243 (.Y (L0_4_L1_1_Fij_nx242), .A0 (nx2654), .A1 (RST)
          , .A2 (nx2646), .B0 (nx2450), .B1 (nx2924)) ;
    inv01 ix2653 (.Y (nx2654), .A (Din[11])) ;
    oai32 L0_4_L1_1_Fij_ix253 (.Y (L0_4_L1_1_Fij_nx252), .A0 (nx2656), .A1 (RST)
          , .A2 (nx2646), .B0 (nx2452), .B1 (nx2924)) ;
    inv01 ix2655 (.Y (nx2656), .A (Din[12])) ;
    oai32 L0_4_L1_1_Fij_ix263 (.Y (L0_4_L1_1_Fij_nx262), .A0 (nx2658), .A1 (RST)
          , .A2 (nx2646), .B0 (nx2454), .B1 (nx2924)) ;
    inv01 ix2657 (.Y (nx2658), .A (Din[13])) ;
    oai32 L0_4_L1_1_Fij_ix273 (.Y (L0_4_L1_1_Fij_nx272), .A0 (nx2660), .A1 (RST)
          , .A2 (nx2662), .B0 (nx2456), .B1 (nx2924)) ;
    inv01 ix2659 (.Y (nx2660), .A (Din[14])) ;
    inv01 ix2661 (.Y (nx2662), .A (L0_4_L1_1_Fij_nx333)) ;
    oai32 L0_4_L1_1_Fij_ix283 (.Y (L0_4_L1_1_Fij_nx282), .A0 (nx2664), .A1 (RST)
          , .A2 (nx2662), .B0 (nx2460), .B1 (nx2926)) ;
    inv01 ix2663 (.Y (nx2664), .A (Din[15])) ;
    oai32 L0_4_L1_1_Wij_ix213 (.Y (L0_4_L1_1_Wij_nx212), .A0 (nx2644), .A1 (RST)
          , .A2 (nx2666), .B0 (nx2462), .B1 (nx2928)) ;
    inv02 ix2665 (.Y (nx2666), .A (L0_4_L1_1_Wij_nx331)) ;
    oai32 L0_4_L1_1_Wij_ix223 (.Y (L0_4_L1_1_Wij_nx222), .A0 (nx2650), .A1 (RST)
          , .A2 (nx2666), .B0 (nx2468), .B1 (nx2928)) ;
    oai32 L0_4_L1_1_Wij_ix233 (.Y (L0_4_L1_1_Wij_nx232), .A0 (nx2652), .A1 (RST)
          , .A2 (nx2666), .B0 (nx2470), .B1 (nx2928)) ;
    oai32 L0_4_L1_1_Wij_ix243 (.Y (L0_4_L1_1_Wij_nx242), .A0 (nx2654), .A1 (RST)
          , .A2 (nx2666), .B0 (nx2472), .B1 (nx2928)) ;
    oai32 L0_4_L1_1_Wij_ix253 (.Y (L0_4_L1_1_Wij_nx252), .A0 (nx2656), .A1 (RST)
          , .A2 (nx2666), .B0 (nx2474), .B1 (nx2928)) ;
    oai32 L0_4_L1_1_Wij_ix263 (.Y (L0_4_L1_1_Wij_nx262), .A0 (nx2658), .A1 (RST)
          , .A2 (nx2666), .B0 (nx2476), .B1 (nx2928)) ;
    oai32 L0_4_L1_1_Wij_ix273 (.Y (L0_4_L1_1_Wij_nx272), .A0 (nx2660), .A1 (RST)
          , .A2 (nx2670), .B0 (nx2478), .B1 (nx2928)) ;
    inv01 ix2669 (.Y (nx2670), .A (L0_4_L1_1_Wij_nx333)) ;
    oai32 L0_4_L1_1_Wij_ix283 (.Y (L0_4_L1_1_Wij_nx282), .A0 (nx2664), .A1 (RST)
          , .A2 (nx2670), .B0 (nx2482), .B1 (nx2930)) ;
    oai32 L0_4_L1_2_Fij_ix213 (.Y (L0_4_L1_2_Fij_nx212), .A0 (nx2672), .A1 (RST)
          , .A2 (nx2674), .B0 (nx2484), .B1 (nx2932)) ;
    inv01 ix2671 (.Y (nx2672), .A (Din[16])) ;
    inv02 ix2673 (.Y (nx2674), .A (L0_4_L1_2_Fij_nx331)) ;
    oai32 L0_4_L1_2_Fij_ix223 (.Y (L0_4_L1_2_Fij_nx222), .A0 (nx2678), .A1 (RST)
          , .A2 (nx2674), .B0 (nx2490), .B1 (nx2932)) ;
    inv01 ix2677 (.Y (nx2678), .A (Din[17])) ;
    oai32 L0_4_L1_2_Fij_ix233 (.Y (L0_4_L1_2_Fij_nx232), .A0 (nx2680), .A1 (RST)
          , .A2 (nx2674), .B0 (nx2492), .B1 (nx2932)) ;
    inv01 ix2679 (.Y (nx2680), .A (Din[18])) ;
    oai32 L0_4_L1_2_Fij_ix243 (.Y (L0_4_L1_2_Fij_nx242), .A0 (nx2682), .A1 (RST)
          , .A2 (nx2674), .B0 (nx2494), .B1 (nx2932)) ;
    inv01 ix2681 (.Y (nx2682), .A (Din[19])) ;
    oai32 L0_4_L1_2_Fij_ix253 (.Y (L0_4_L1_2_Fij_nx252), .A0 (nx2684), .A1 (RST)
          , .A2 (nx2674), .B0 (nx2496), .B1 (nx2932)) ;
    inv01 ix2683 (.Y (nx2684), .A (Din[20])) ;
    oai32 L0_4_L1_2_Fij_ix263 (.Y (L0_4_L1_2_Fij_nx262), .A0 (nx2686), .A1 (RST)
          , .A2 (nx2674), .B0 (nx2498), .B1 (nx2932)) ;
    inv01 ix2685 (.Y (nx2686), .A (Din[21])) ;
    oai32 L0_4_L1_2_Fij_ix273 (.Y (L0_4_L1_2_Fij_nx272), .A0 (nx2688), .A1 (RST)
          , .A2 (nx2690), .B0 (nx2500), .B1 (nx2932)) ;
    inv01 ix2687 (.Y (nx2688), .A (Din[22])) ;
    inv01 ix2689 (.Y (nx2690), .A (L0_4_L1_2_Fij_nx333)) ;
    oai32 L0_4_L1_2_Fij_ix283 (.Y (L0_4_L1_2_Fij_nx282), .A0 (nx2692), .A1 (RST)
          , .A2 (nx2690), .B0 (nx2504), .B1 (nx2934)) ;
    inv01 ix2691 (.Y (nx2692), .A (Din[23])) ;
    oai32 L0_4_L1_2_Wij_ix213 (.Y (L0_4_L1_2_Wij_nx212), .A0 (nx2672), .A1 (RST)
          , .A2 (nx2694), .B0 (nx2506), .B1 (nx2936)) ;
    inv02 ix2693 (.Y (nx2694), .A (L0_4_L1_2_Wij_nx331)) ;
    oai32 L0_4_L1_2_Wij_ix223 (.Y (L0_4_L1_2_Wij_nx222), .A0 (nx2678), .A1 (RST)
          , .A2 (nx2694), .B0 (nx2512), .B1 (nx2936)) ;
    oai32 L0_4_L1_2_Wij_ix233 (.Y (L0_4_L1_2_Wij_nx232), .A0 (nx2680), .A1 (RST)
          , .A2 (nx2694), .B0 (nx2514), .B1 (nx2936)) ;
    oai32 L0_4_L1_2_Wij_ix243 (.Y (L0_4_L1_2_Wij_nx242), .A0 (nx2682), .A1 (RST)
          , .A2 (nx2694), .B0 (nx2516), .B1 (nx2936)) ;
    oai32 L0_4_L1_2_Wij_ix253 (.Y (L0_4_L1_2_Wij_nx252), .A0 (nx2684), .A1 (RST)
          , .A2 (nx2694), .B0 (nx2518), .B1 (nx2936)) ;
    oai32 L0_4_L1_2_Wij_ix263 (.Y (L0_4_L1_2_Wij_nx262), .A0 (nx2686), .A1 (RST)
          , .A2 (nx2694), .B0 (nx2520), .B1 (nx2936)) ;
    oai32 L0_4_L1_2_Wij_ix273 (.Y (L0_4_L1_2_Wij_nx272), .A0 (nx2688), .A1 (RST)
          , .A2 (nx2698), .B0 (nx2522), .B1 (nx2936)) ;
    inv01 ix2697 (.Y (nx2698), .A (L0_4_L1_2_Wij_nx333)) ;
    oai32 L0_4_L1_2_Wij_ix283 (.Y (L0_4_L1_2_Wij_nx282), .A0 (nx2692), .A1 (RST)
          , .A2 (nx2698), .B0 (nx2526), .B1 (nx2938)) ;
    oai32 L0_4_L1_3_Fij_ix213 (.Y (L0_4_L1_3_Fij_nx212), .A0 (nx2700), .A1 (RST)
          , .A2 (nx2702), .B0 (nx2528), .B1 (nx2940)) ;
    inv01 ix2699 (.Y (nx2700), .A (Din[24])) ;
    inv02 ix2701 (.Y (nx2702), .A (L0_4_L1_3_Fij_nx331)) ;
    oai32 L0_4_L1_3_Fij_ix223 (.Y (L0_4_L1_3_Fij_nx222), .A0 (nx2706), .A1 (RST)
          , .A2 (nx2702), .B0 (nx2534), .B1 (nx2940)) ;
    inv01 ix2705 (.Y (nx2706), .A (Din[25])) ;
    oai32 L0_4_L1_3_Fij_ix233 (.Y (L0_4_L1_3_Fij_nx232), .A0 (nx2708), .A1 (RST)
          , .A2 (nx2702), .B0 (nx2536), .B1 (nx2940)) ;
    inv01 ix2707 (.Y (nx2708), .A (Din[26])) ;
    oai32 L0_4_L1_3_Fij_ix243 (.Y (L0_4_L1_3_Fij_nx242), .A0 (nx2710), .A1 (RST)
          , .A2 (nx2702), .B0 (nx2538), .B1 (nx2940)) ;
    inv01 ix2709 (.Y (nx2710), .A (Din[27])) ;
    oai32 L0_4_L1_3_Fij_ix253 (.Y (L0_4_L1_3_Fij_nx252), .A0 (nx2712), .A1 (RST)
          , .A2 (nx2702), .B0 (nx2540), .B1 (nx2940)) ;
    inv01 ix2711 (.Y (nx2712), .A (Din[28])) ;
    oai32 L0_4_L1_3_Fij_ix263 (.Y (L0_4_L1_3_Fij_nx262), .A0 (nx2714), .A1 (RST)
          , .A2 (nx2702), .B0 (nx2542), .B1 (nx2940)) ;
    inv01 ix2713 (.Y (nx2714), .A (Din[29])) ;
    oai32 L0_4_L1_3_Fij_ix273 (.Y (L0_4_L1_3_Fij_nx272), .A0 (nx2716), .A1 (RST)
          , .A2 (nx2718), .B0 (nx2544), .B1 (nx2940)) ;
    inv01 ix2715 (.Y (nx2716), .A (Din[30])) ;
    inv01 ix2717 (.Y (nx2718), .A (L0_4_L1_3_Fij_nx333)) ;
    oai32 L0_4_L1_3_Fij_ix283 (.Y (L0_4_L1_3_Fij_nx282), .A0 (nx2720), .A1 (RST)
          , .A2 (nx2718), .B0 (nx2548), .B1 (nx2942)) ;
    inv01 ix2719 (.Y (nx2720), .A (Din[31])) ;
    oai32 L0_4_L1_3_Wij_ix213 (.Y (L0_4_L1_3_Wij_nx212), .A0 (nx2700), .A1 (RST)
          , .A2 (nx2722), .B0 (nx2550), .B1 (nx2944)) ;
    inv02 ix2721 (.Y (nx2722), .A (L0_4_L1_3_Wij_nx331)) ;
    oai32 L0_4_L1_3_Wij_ix223 (.Y (L0_4_L1_3_Wij_nx222), .A0 (nx2706), .A1 (RST)
          , .A2 (nx2722), .B0 (nx2556), .B1 (nx2944)) ;
    oai32 L0_4_L1_3_Wij_ix233 (.Y (L0_4_L1_3_Wij_nx232), .A0 (nx2708), .A1 (RST)
          , .A2 (nx2722), .B0 (nx2558), .B1 (nx2944)) ;
    oai32 L0_4_L1_3_Wij_ix243 (.Y (L0_4_L1_3_Wij_nx242), .A0 (nx2710), .A1 (RST)
          , .A2 (nx2722), .B0 (nx2560), .B1 (nx2944)) ;
    oai32 L0_4_L1_3_Wij_ix253 (.Y (L0_4_L1_3_Wij_nx252), .A0 (nx2712), .A1 (RST)
          , .A2 (nx2722), .B0 (nx2562), .B1 (nx2944)) ;
    oai32 L0_4_L1_3_Wij_ix263 (.Y (L0_4_L1_3_Wij_nx262), .A0 (nx2714), .A1 (RST)
          , .A2 (nx2722), .B0 (nx2564), .B1 (nx2944)) ;
    oai32 L0_4_L1_3_Wij_ix273 (.Y (L0_4_L1_3_Wij_nx272), .A0 (nx2716), .A1 (RST)
          , .A2 (nx2726), .B0 (nx2566), .B1 (nx2944)) ;
    inv01 ix2725 (.Y (nx2726), .A (L0_4_L1_3_Wij_nx333)) ;
    oai32 L0_4_L1_3_Wij_ix283 (.Y (L0_4_L1_3_Wij_nx282), .A0 (nx2720), .A1 (RST)
          , .A2 (nx2726), .B0 (nx2570), .B1 (nx2946)) ;
    oai32 L0_4_L1_4_Fij_ix213 (.Y (L0_4_L1_4_Fij_nx212), .A0 (nx2728), .A1 (RST)
          , .A2 (nx2730), .B0 (nx2572), .B1 (nx2948)) ;
    inv01 ix2727 (.Y (nx2728), .A (Din[32])) ;
    inv02 ix2729 (.Y (nx2730), .A (L0_4_L1_4_Fij_nx331)) ;
    oai32 L0_4_L1_4_Fij_ix223 (.Y (L0_4_L1_4_Fij_nx222), .A0 (nx2734), .A1 (RST)
          , .A2 (nx2730), .B0 (nx2578), .B1 (nx2948)) ;
    inv01 ix2733 (.Y (nx2734), .A (Din[33])) ;
    oai32 L0_4_L1_4_Fij_ix233 (.Y (L0_4_L1_4_Fij_nx232), .A0 (nx2736), .A1 (RST)
          , .A2 (nx2730), .B0 (nx2580), .B1 (nx2948)) ;
    inv01 ix2735 (.Y (nx2736), .A (Din[34])) ;
    oai32 L0_4_L1_4_Fij_ix243 (.Y (L0_4_L1_4_Fij_nx242), .A0 (nx2738), .A1 (RST)
          , .A2 (nx2730), .B0 (nx2582), .B1 (nx2948)) ;
    inv01 ix2737 (.Y (nx2738), .A (Din[35])) ;
    oai32 L0_4_L1_4_Fij_ix253 (.Y (L0_4_L1_4_Fij_nx252), .A0 (nx2740), .A1 (RST)
          , .A2 (nx2730), .B0 (nx2584), .B1 (nx2948)) ;
    inv01 ix2739 (.Y (nx2740), .A (Din[36])) ;
    oai32 L0_4_L1_4_Fij_ix263 (.Y (L0_4_L1_4_Fij_nx262), .A0 (nx2742), .A1 (RST)
          , .A2 (nx2730), .B0 (nx2586), .B1 (nx2948)) ;
    inv01 ix2741 (.Y (nx2742), .A (Din[37])) ;
    oai32 L0_4_L1_4_Fij_ix273 (.Y (L0_4_L1_4_Fij_nx272), .A0 (nx2744), .A1 (RST)
          , .A2 (nx2746), .B0 (nx2588), .B1 (nx2948)) ;
    inv01 ix2743 (.Y (nx2744), .A (Din[38])) ;
    inv01 ix2745 (.Y (nx2746), .A (L0_4_L1_4_Fij_nx333)) ;
    oai32 L0_4_L1_4_Fij_ix283 (.Y (L0_4_L1_4_Fij_nx282), .A0 (nx2748), .A1 (RST)
          , .A2 (nx2746), .B0 (nx2592), .B1 (nx2950)) ;
    inv01 ix2747 (.Y (nx2748), .A (Din[39])) ;
    oai32 L0_4_L1_4_Wij_ix213 (.Y (L0_4_L1_4_Wij_nx212), .A0 (nx2728), .A1 (RST)
          , .A2 (nx2750), .B0 (nx2594), .B1 (nx2952)) ;
    inv02 ix2749 (.Y (nx2750), .A (L0_4_L1_4_Wij_nx331)) ;
    oai32 L0_4_L1_4_Wij_ix223 (.Y (L0_4_L1_4_Wij_nx222), .A0 (nx2734), .A1 (RST)
          , .A2 (nx2750), .B0 (nx2600), .B1 (nx2952)) ;
    oai32 L0_4_L1_4_Wij_ix233 (.Y (L0_4_L1_4_Wij_nx232), .A0 (nx2736), .A1 (RST)
          , .A2 (nx2750), .B0 (nx2602), .B1 (nx2952)) ;
    oai32 L0_4_L1_4_Wij_ix243 (.Y (L0_4_L1_4_Wij_nx242), .A0 (nx2738), .A1 (RST)
          , .A2 (nx2750), .B0 (nx2604), .B1 (nx2952)) ;
    oai32 L0_4_L1_4_Wij_ix253 (.Y (L0_4_L1_4_Wij_nx252), .A0 (nx2740), .A1 (RST)
          , .A2 (nx2750), .B0 (nx2606), .B1 (nx2952)) ;
    oai32 L0_4_L1_4_Wij_ix263 (.Y (L0_4_L1_4_Wij_nx262), .A0 (nx2742), .A1 (RST)
          , .A2 (nx2750), .B0 (nx2608), .B1 (nx2952)) ;
    oai32 L0_4_L1_4_Wij_ix273 (.Y (L0_4_L1_4_Wij_nx272), .A0 (nx2744), .A1 (RST)
          , .A2 (nx2754), .B0 (nx2610), .B1 (nx2952)) ;
    inv01 ix2753 (.Y (nx2754), .A (L0_4_L1_4_Wij_nx333)) ;
    oai32 L0_4_L1_4_Wij_ix283 (.Y (L0_4_L1_4_Wij_nx282), .A0 (nx2748), .A1 (RST)
          , .A2 (nx2754), .B0 (nx2614), .B1 (nx2954)) ;
    inv02 ix2755 (.Y (nx2756), .A (L0_0_L1_0_Fij_nx296)) ;
    inv02 ix2757 (.Y (nx2758), .A (L0_0_L1_0_Fij_nx296)) ;
    inv02 ix2759 (.Y (nx2760), .A (L0_0_L1_0_Wij_nx296)) ;
    inv02 ix2761 (.Y (nx2762), .A (L0_0_L1_0_Wij_nx296)) ;
    inv02 ix2763 (.Y (nx2764), .A (L0_0_L1_1_Fij_nx296)) ;
    inv02 ix2765 (.Y (nx2766), .A (L0_0_L1_1_Fij_nx296)) ;
    inv02 ix2767 (.Y (nx2768), .A (L0_0_L1_1_Wij_nx296)) ;
    inv02 ix2769 (.Y (nx2770), .A (L0_0_L1_1_Wij_nx296)) ;
    inv02 ix2771 (.Y (nx2772), .A (L0_0_L1_2_Fij_nx296)) ;
    inv02 ix2773 (.Y (nx2774), .A (L0_0_L1_2_Fij_nx296)) ;
    inv02 ix2775 (.Y (nx2776), .A (L0_0_L1_2_Wij_nx296)) ;
    inv02 ix2777 (.Y (nx2778), .A (L0_0_L1_2_Wij_nx296)) ;
    inv02 ix2779 (.Y (nx2780), .A (L0_0_L1_3_Fij_nx296)) ;
    inv02 ix2781 (.Y (nx2782), .A (L0_0_L1_3_Fij_nx296)) ;
    inv02 ix2783 (.Y (nx2784), .A (L0_0_L1_3_Wij_nx296)) ;
    inv02 ix2785 (.Y (nx2786), .A (L0_0_L1_3_Wij_nx296)) ;
    inv02 ix2787 (.Y (nx2788), .A (L0_0_L1_4_Fij_nx296)) ;
    inv02 ix2789 (.Y (nx2790), .A (L0_0_L1_4_Fij_nx296)) ;
    inv02 ix2791 (.Y (nx2792), .A (L0_0_L1_4_Wij_nx296)) ;
    inv02 ix2793 (.Y (nx2794), .A (L0_0_L1_4_Wij_nx296)) ;
    inv02 ix2795 (.Y (nx2796), .A (L0_1_L1_0_Fij_nx296)) ;
    inv02 ix2797 (.Y (nx2798), .A (L0_1_L1_0_Fij_nx296)) ;
    inv02 ix2799 (.Y (nx2800), .A (L0_1_L1_0_Wij_nx296)) ;
    inv02 ix2801 (.Y (nx2802), .A (L0_1_L1_0_Wij_nx296)) ;
    inv02 ix2803 (.Y (nx2804), .A (L0_1_L1_1_Fij_nx296)) ;
    inv02 ix2805 (.Y (nx2806), .A (L0_1_L1_1_Fij_nx296)) ;
    inv02 ix2807 (.Y (nx2808), .A (L0_1_L1_1_Wij_nx296)) ;
    inv02 ix2809 (.Y (nx2810), .A (L0_1_L1_1_Wij_nx296)) ;
    inv02 ix2811 (.Y (nx2812), .A (L0_1_L1_2_Fij_nx296)) ;
    inv02 ix2813 (.Y (nx2814), .A (L0_1_L1_2_Fij_nx296)) ;
    inv02 ix2815 (.Y (nx2816), .A (L0_1_L1_2_Wij_nx296)) ;
    inv02 ix2817 (.Y (nx2818), .A (L0_1_L1_2_Wij_nx296)) ;
    inv02 ix2819 (.Y (nx2820), .A (L0_1_L1_3_Fij_nx296)) ;
    inv02 ix2821 (.Y (nx2822), .A (L0_1_L1_3_Fij_nx296)) ;
    inv02 ix2823 (.Y (nx2824), .A (L0_1_L1_3_Wij_nx296)) ;
    inv02 ix2825 (.Y (nx2826), .A (L0_1_L1_3_Wij_nx296)) ;
    inv02 ix2827 (.Y (nx2828), .A (L0_1_L1_4_Fij_nx296)) ;
    inv02 ix2829 (.Y (nx2830), .A (L0_1_L1_4_Fij_nx296)) ;
    inv02 ix2831 (.Y (nx2832), .A (L0_1_L1_4_Wij_nx296)) ;
    inv02 ix2833 (.Y (nx2834), .A (L0_1_L1_4_Wij_nx296)) ;
    inv02 ix2835 (.Y (nx2836), .A (L0_2_L1_0_Fij_nx296)) ;
    inv02 ix2837 (.Y (nx2838), .A (L0_2_L1_0_Fij_nx296)) ;
    inv02 ix2839 (.Y (nx2840), .A (L0_2_L1_0_Wij_nx296)) ;
    inv02 ix2841 (.Y (nx2842), .A (L0_2_L1_0_Wij_nx296)) ;
    inv02 ix2843 (.Y (nx2844), .A (L0_2_L1_1_Fij_nx296)) ;
    inv02 ix2845 (.Y (nx2846), .A (L0_2_L1_1_Fij_nx296)) ;
    inv02 ix2847 (.Y (nx2848), .A (L0_2_L1_1_Wij_nx296)) ;
    inv02 ix2849 (.Y (nx2850), .A (L0_2_L1_1_Wij_nx296)) ;
    inv02 ix2851 (.Y (nx2852), .A (L0_2_L1_2_Fij_nx296)) ;
    inv02 ix2853 (.Y (nx2854), .A (L0_2_L1_2_Fij_nx296)) ;
    inv02 ix2855 (.Y (nx2856), .A (L0_2_L1_2_Wij_nx296)) ;
    inv02 ix2857 (.Y (nx2858), .A (L0_2_L1_2_Wij_nx296)) ;
    inv02 ix2859 (.Y (nx2860), .A (L0_2_L1_3_Fij_nx296)) ;
    inv02 ix2861 (.Y (nx2862), .A (L0_2_L1_3_Fij_nx296)) ;
    inv02 ix2863 (.Y (nx2864), .A (L0_2_L1_3_Wij_nx296)) ;
    inv02 ix2865 (.Y (nx2866), .A (L0_2_L1_3_Wij_nx296)) ;
    inv02 ix2867 (.Y (nx2868), .A (L0_2_L1_4_Fij_nx296)) ;
    inv02 ix2869 (.Y (nx2870), .A (L0_2_L1_4_Fij_nx296)) ;
    inv02 ix2871 (.Y (nx2872), .A (L0_2_L1_4_Wij_nx296)) ;
    inv02 ix2873 (.Y (nx2874), .A (L0_2_L1_4_Wij_nx296)) ;
    inv02 ix2875 (.Y (nx2876), .A (L0_3_L1_0_Fij_nx296)) ;
    inv02 ix2877 (.Y (nx2878), .A (L0_3_L1_0_Fij_nx296)) ;
    inv02 ix2879 (.Y (nx2880), .A (L0_3_L1_0_Wij_nx296)) ;
    inv02 ix2881 (.Y (nx2882), .A (L0_3_L1_0_Wij_nx296)) ;
    inv02 ix2883 (.Y (nx2884), .A (L0_3_L1_1_Fij_nx296)) ;
    inv02 ix2885 (.Y (nx2886), .A (L0_3_L1_1_Fij_nx296)) ;
    inv02 ix2887 (.Y (nx2888), .A (L0_3_L1_1_Wij_nx296)) ;
    inv02 ix2889 (.Y (nx2890), .A (L0_3_L1_1_Wij_nx296)) ;
    inv02 ix2891 (.Y (nx2892), .A (L0_3_L1_2_Fij_nx296)) ;
    inv02 ix2893 (.Y (nx2894), .A (L0_3_L1_2_Fij_nx296)) ;
    inv02 ix2895 (.Y (nx2896), .A (L0_3_L1_2_Wij_nx296)) ;
    inv02 ix2897 (.Y (nx2898), .A (L0_3_L1_2_Wij_nx296)) ;
    inv02 ix2899 (.Y (nx2900), .A (L0_3_L1_3_Fij_nx296)) ;
    inv02 ix2901 (.Y (nx2902), .A (L0_3_L1_3_Fij_nx296)) ;
    inv02 ix2903 (.Y (nx2904), .A (L0_3_L1_3_Wij_nx296)) ;
    inv02 ix2905 (.Y (nx2906), .A (L0_3_L1_3_Wij_nx296)) ;
    inv02 ix2907 (.Y (nx2908), .A (L0_3_L1_4_Fij_nx296)) ;
    inv02 ix2909 (.Y (nx2910), .A (L0_3_L1_4_Fij_nx296)) ;
    inv02 ix2911 (.Y (nx2912), .A (L0_3_L1_4_Wij_nx296)) ;
    inv02 ix2913 (.Y (nx2914), .A (L0_3_L1_4_Wij_nx296)) ;
    inv02 ix2915 (.Y (nx2916), .A (L0_4_L1_0_Fij_nx296)) ;
    inv02 ix2917 (.Y (nx2918), .A (L0_4_L1_0_Fij_nx296)) ;
    inv02 ix2919 (.Y (nx2920), .A (L0_4_L1_0_Wij_nx296)) ;
    inv02 ix2921 (.Y (nx2922), .A (L0_4_L1_0_Wij_nx296)) ;
    inv02 ix2923 (.Y (nx2924), .A (L0_4_L1_1_Fij_nx296)) ;
    inv02 ix2925 (.Y (nx2926), .A (L0_4_L1_1_Fij_nx296)) ;
    inv02 ix2927 (.Y (nx2928), .A (L0_4_L1_1_Wij_nx296)) ;
    inv02 ix2929 (.Y (nx2930), .A (L0_4_L1_1_Wij_nx296)) ;
    inv02 ix2931 (.Y (nx2932), .A (L0_4_L1_2_Fij_nx296)) ;
    inv02 ix2933 (.Y (nx2934), .A (L0_4_L1_2_Fij_nx296)) ;
    inv02 ix2935 (.Y (nx2936), .A (L0_4_L1_2_Wij_nx296)) ;
    inv02 ix2937 (.Y (nx2938), .A (L0_4_L1_2_Wij_nx296)) ;
    inv02 ix2939 (.Y (nx2940), .A (L0_4_L1_3_Fij_nx296)) ;
    inv02 ix2941 (.Y (nx2942), .A (L0_4_L1_3_Fij_nx296)) ;
    inv02 ix2943 (.Y (nx2944), .A (L0_4_L1_3_Wij_nx296)) ;
    inv02 ix2945 (.Y (nx2946), .A (L0_4_L1_3_Wij_nx296)) ;
    inv02 ix2947 (.Y (nx2948), .A (L0_4_L1_4_Fij_nx296)) ;
    inv02 ix2949 (.Y (nx2950), .A (L0_4_L1_4_Fij_nx296)) ;
    inv02 ix2951 (.Y (nx2952), .A (L0_4_L1_4_Wij_nx296)) ;
    inv02 ix2953 (.Y (nx2954), .A (L0_4_L1_4_Wij_nx296)) ;
endmodule

