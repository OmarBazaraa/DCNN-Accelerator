//
// Verilog description for cell cache, 
// Wed May  2 09:48:18 2018
//
// LeonardoSpectrum Level 3, 2017a.2 
//


module cache ( CLK, RST, FilterSize, FilterWR, WindowWR, Din, FilterDout_0__0__7, 
               FilterDout_0__0__6, FilterDout_0__0__5, FilterDout_0__0__4, 
               FilterDout_0__0__3, FilterDout_0__0__2, FilterDout_0__0__1, 
               FilterDout_0__0__0, FilterDout_0__1__7, FilterDout_0__1__6, 
               FilterDout_0__1__5, FilterDout_0__1__4, FilterDout_0__1__3, 
               FilterDout_0__1__2, FilterDout_0__1__1, FilterDout_0__1__0, 
               FilterDout_0__2__7, FilterDout_0__2__6, FilterDout_0__2__5, 
               FilterDout_0__2__4, FilterDout_0__2__3, FilterDout_0__2__2, 
               FilterDout_0__2__1, FilterDout_0__2__0, FilterDout_0__3__7, 
               FilterDout_0__3__6, FilterDout_0__3__5, FilterDout_0__3__4, 
               FilterDout_0__3__3, FilterDout_0__3__2, FilterDout_0__3__1, 
               FilterDout_0__3__0, FilterDout_0__4__7, FilterDout_0__4__6, 
               FilterDout_0__4__5, FilterDout_0__4__4, FilterDout_0__4__3, 
               FilterDout_0__4__2, FilterDout_0__4__1, FilterDout_0__4__0, 
               FilterDout_1__0__7, FilterDout_1__0__6, FilterDout_1__0__5, 
               FilterDout_1__0__4, FilterDout_1__0__3, FilterDout_1__0__2, 
               FilterDout_1__0__1, FilterDout_1__0__0, FilterDout_1__1__7, 
               FilterDout_1__1__6, FilterDout_1__1__5, FilterDout_1__1__4, 
               FilterDout_1__1__3, FilterDout_1__1__2, FilterDout_1__1__1, 
               FilterDout_1__1__0, FilterDout_1__2__7, FilterDout_1__2__6, 
               FilterDout_1__2__5, FilterDout_1__2__4, FilterDout_1__2__3, 
               FilterDout_1__2__2, FilterDout_1__2__1, FilterDout_1__2__0, 
               FilterDout_1__3__7, FilterDout_1__3__6, FilterDout_1__3__5, 
               FilterDout_1__3__4, FilterDout_1__3__3, FilterDout_1__3__2, 
               FilterDout_1__3__1, FilterDout_1__3__0, FilterDout_1__4__7, 
               FilterDout_1__4__6, FilterDout_1__4__5, FilterDout_1__4__4, 
               FilterDout_1__4__3, FilterDout_1__4__2, FilterDout_1__4__1, 
               FilterDout_1__4__0, FilterDout_2__0__7, FilterDout_2__0__6, 
               FilterDout_2__0__5, FilterDout_2__0__4, FilterDout_2__0__3, 
               FilterDout_2__0__2, FilterDout_2__0__1, FilterDout_2__0__0, 
               FilterDout_2__1__7, FilterDout_2__1__6, FilterDout_2__1__5, 
               FilterDout_2__1__4, FilterDout_2__1__3, FilterDout_2__1__2, 
               FilterDout_2__1__1, FilterDout_2__1__0, FilterDout_2__2__7, 
               FilterDout_2__2__6, FilterDout_2__2__5, FilterDout_2__2__4, 
               FilterDout_2__2__3, FilterDout_2__2__2, FilterDout_2__2__1, 
               FilterDout_2__2__0, FilterDout_2__3__7, FilterDout_2__3__6, 
               FilterDout_2__3__5, FilterDout_2__3__4, FilterDout_2__3__3, 
               FilterDout_2__3__2, FilterDout_2__3__1, FilterDout_2__3__0, 
               FilterDout_2__4__7, FilterDout_2__4__6, FilterDout_2__4__5, 
               FilterDout_2__4__4, FilterDout_2__4__3, FilterDout_2__4__2, 
               FilterDout_2__4__1, FilterDout_2__4__0, FilterDout_3__0__7, 
               FilterDout_3__0__6, FilterDout_3__0__5, FilterDout_3__0__4, 
               FilterDout_3__0__3, FilterDout_3__0__2, FilterDout_3__0__1, 
               FilterDout_3__0__0, FilterDout_3__1__7, FilterDout_3__1__6, 
               FilterDout_3__1__5, FilterDout_3__1__4, FilterDout_3__1__3, 
               FilterDout_3__1__2, FilterDout_3__1__1, FilterDout_3__1__0, 
               FilterDout_3__2__7, FilterDout_3__2__6, FilterDout_3__2__5, 
               FilterDout_3__2__4, FilterDout_3__2__3, FilterDout_3__2__2, 
               FilterDout_3__2__1, FilterDout_3__2__0, FilterDout_3__3__7, 
               FilterDout_3__3__6, FilterDout_3__3__5, FilterDout_3__3__4, 
               FilterDout_3__3__3, FilterDout_3__3__2, FilterDout_3__3__1, 
               FilterDout_3__3__0, FilterDout_3__4__7, FilterDout_3__4__6, 
               FilterDout_3__4__5, FilterDout_3__4__4, FilterDout_3__4__3, 
               FilterDout_3__4__2, FilterDout_3__4__1, FilterDout_3__4__0, 
               FilterDout_4__0__7, FilterDout_4__0__6, FilterDout_4__0__5, 
               FilterDout_4__0__4, FilterDout_4__0__3, FilterDout_4__0__2, 
               FilterDout_4__0__1, FilterDout_4__0__0, FilterDout_4__1__7, 
               FilterDout_4__1__6, FilterDout_4__1__5, FilterDout_4__1__4, 
               FilterDout_4__1__3, FilterDout_4__1__2, FilterDout_4__1__1, 
               FilterDout_4__1__0, FilterDout_4__2__7, FilterDout_4__2__6, 
               FilterDout_4__2__5, FilterDout_4__2__4, FilterDout_4__2__3, 
               FilterDout_4__2__2, FilterDout_4__2__1, FilterDout_4__2__0, 
               FilterDout_4__3__7, FilterDout_4__3__6, FilterDout_4__3__5, 
               FilterDout_4__3__4, FilterDout_4__3__3, FilterDout_4__3__2, 
               FilterDout_4__3__1, FilterDout_4__3__0, FilterDout_4__4__7, 
               FilterDout_4__4__6, FilterDout_4__4__5, FilterDout_4__4__4, 
               FilterDout_4__4__3, FilterDout_4__4__2, FilterDout_4__4__1, 
               FilterDout_4__4__0, WindowDout_0__0__7, WindowDout_0__0__6, 
               WindowDout_0__0__5, WindowDout_0__0__4, WindowDout_0__0__3, 
               WindowDout_0__0__2, WindowDout_0__0__1, WindowDout_0__0__0, 
               WindowDout_0__1__7, WindowDout_0__1__6, WindowDout_0__1__5, 
               WindowDout_0__1__4, WindowDout_0__1__3, WindowDout_0__1__2, 
               WindowDout_0__1__1, WindowDout_0__1__0, WindowDout_0__2__7, 
               WindowDout_0__2__6, WindowDout_0__2__5, WindowDout_0__2__4, 
               WindowDout_0__2__3, WindowDout_0__2__2, WindowDout_0__2__1, 
               WindowDout_0__2__0, WindowDout_0__3__7, WindowDout_0__3__6, 
               WindowDout_0__3__5, WindowDout_0__3__4, WindowDout_0__3__3, 
               WindowDout_0__3__2, WindowDout_0__3__1, WindowDout_0__3__0, 
               WindowDout_0__4__7, WindowDout_0__4__6, WindowDout_0__4__5, 
               WindowDout_0__4__4, WindowDout_0__4__3, WindowDout_0__4__2, 
               WindowDout_0__4__1, WindowDout_0__4__0, WindowDout_1__0__7, 
               WindowDout_1__0__6, WindowDout_1__0__5, WindowDout_1__0__4, 
               WindowDout_1__0__3, WindowDout_1__0__2, WindowDout_1__0__1, 
               WindowDout_1__0__0, WindowDout_1__1__7, WindowDout_1__1__6, 
               WindowDout_1__1__5, WindowDout_1__1__4, WindowDout_1__1__3, 
               WindowDout_1__1__2, WindowDout_1__1__1, WindowDout_1__1__0, 
               WindowDout_1__2__7, WindowDout_1__2__6, WindowDout_1__2__5, 
               WindowDout_1__2__4, WindowDout_1__2__3, WindowDout_1__2__2, 
               WindowDout_1__2__1, WindowDout_1__2__0, WindowDout_1__3__7, 
               WindowDout_1__3__6, WindowDout_1__3__5, WindowDout_1__3__4, 
               WindowDout_1__3__3, WindowDout_1__3__2, WindowDout_1__3__1, 
               WindowDout_1__3__0, WindowDout_1__4__7, WindowDout_1__4__6, 
               WindowDout_1__4__5, WindowDout_1__4__4, WindowDout_1__4__3, 
               WindowDout_1__4__2, WindowDout_1__4__1, WindowDout_1__4__0, 
               WindowDout_2__0__7, WindowDout_2__0__6, WindowDout_2__0__5, 
               WindowDout_2__0__4, WindowDout_2__0__3, WindowDout_2__0__2, 
               WindowDout_2__0__1, WindowDout_2__0__0, WindowDout_2__1__7, 
               WindowDout_2__1__6, WindowDout_2__1__5, WindowDout_2__1__4, 
               WindowDout_2__1__3, WindowDout_2__1__2, WindowDout_2__1__1, 
               WindowDout_2__1__0, WindowDout_2__2__7, WindowDout_2__2__6, 
               WindowDout_2__2__5, WindowDout_2__2__4, WindowDout_2__2__3, 
               WindowDout_2__2__2, WindowDout_2__2__1, WindowDout_2__2__0, 
               WindowDout_2__3__7, WindowDout_2__3__6, WindowDout_2__3__5, 
               WindowDout_2__3__4, WindowDout_2__3__3, WindowDout_2__3__2, 
               WindowDout_2__3__1, WindowDout_2__3__0, WindowDout_2__4__7, 
               WindowDout_2__4__6, WindowDout_2__4__5, WindowDout_2__4__4, 
               WindowDout_2__4__3, WindowDout_2__4__2, WindowDout_2__4__1, 
               WindowDout_2__4__0, WindowDout_3__0__7, WindowDout_3__0__6, 
               WindowDout_3__0__5, WindowDout_3__0__4, WindowDout_3__0__3, 
               WindowDout_3__0__2, WindowDout_3__0__1, WindowDout_3__0__0, 
               WindowDout_3__1__7, WindowDout_3__1__6, WindowDout_3__1__5, 
               WindowDout_3__1__4, WindowDout_3__1__3, WindowDout_3__1__2, 
               WindowDout_3__1__1, WindowDout_3__1__0, WindowDout_3__2__7, 
               WindowDout_3__2__6, WindowDout_3__2__5, WindowDout_3__2__4, 
               WindowDout_3__2__3, WindowDout_3__2__2, WindowDout_3__2__1, 
               WindowDout_3__2__0, WindowDout_3__3__7, WindowDout_3__3__6, 
               WindowDout_3__3__5, WindowDout_3__3__4, WindowDout_3__3__3, 
               WindowDout_3__3__2, WindowDout_3__3__1, WindowDout_3__3__0, 
               WindowDout_3__4__7, WindowDout_3__4__6, WindowDout_3__4__5, 
               WindowDout_3__4__4, WindowDout_3__4__3, WindowDout_3__4__2, 
               WindowDout_3__4__1, WindowDout_3__4__0, WindowDout_4__0__7, 
               WindowDout_4__0__6, WindowDout_4__0__5, WindowDout_4__0__4, 
               WindowDout_4__0__3, WindowDout_4__0__2, WindowDout_4__0__1, 
               WindowDout_4__0__0, WindowDout_4__1__7, WindowDout_4__1__6, 
               WindowDout_4__1__5, WindowDout_4__1__4, WindowDout_4__1__3, 
               WindowDout_4__1__2, WindowDout_4__1__1, WindowDout_4__1__0, 
               WindowDout_4__2__7, WindowDout_4__2__6, WindowDout_4__2__5, 
               WindowDout_4__2__4, WindowDout_4__2__3, WindowDout_4__2__2, 
               WindowDout_4__2__1, WindowDout_4__2__0, WindowDout_4__3__7, 
               WindowDout_4__3__6, WindowDout_4__3__5, WindowDout_4__3__4, 
               WindowDout_4__3__3, WindowDout_4__3__2, WindowDout_4__3__1, 
               WindowDout_4__3__0, WindowDout_4__4__7, WindowDout_4__4__6, 
               WindowDout_4__4__5, WindowDout_4__4__4, WindowDout_4__4__3, 
               WindowDout_4__4__2, WindowDout_4__4__1, WindowDout_4__4__0, 
               ResultWR, ResultDin, ResultDout ) ;

    input CLK ;
    input RST ;
    input FilterSize ;
    input FilterWR ;
    input WindowWR ;
    input [39:0]Din ;
    output FilterDout_0__0__7 ;
    output FilterDout_0__0__6 ;
    output FilterDout_0__0__5 ;
    output FilterDout_0__0__4 ;
    output FilterDout_0__0__3 ;
    output FilterDout_0__0__2 ;
    output FilterDout_0__0__1 ;
    output FilterDout_0__0__0 ;
    output FilterDout_0__1__7 ;
    output FilterDout_0__1__6 ;
    output FilterDout_0__1__5 ;
    output FilterDout_0__1__4 ;
    output FilterDout_0__1__3 ;
    output FilterDout_0__1__2 ;
    output FilterDout_0__1__1 ;
    output FilterDout_0__1__0 ;
    output FilterDout_0__2__7 ;
    output FilterDout_0__2__6 ;
    output FilterDout_0__2__5 ;
    output FilterDout_0__2__4 ;
    output FilterDout_0__2__3 ;
    output FilterDout_0__2__2 ;
    output FilterDout_0__2__1 ;
    output FilterDout_0__2__0 ;
    output FilterDout_0__3__7 ;
    output FilterDout_0__3__6 ;
    output FilterDout_0__3__5 ;
    output FilterDout_0__3__4 ;
    output FilterDout_0__3__3 ;
    output FilterDout_0__3__2 ;
    output FilterDout_0__3__1 ;
    output FilterDout_0__3__0 ;
    output FilterDout_0__4__7 ;
    output FilterDout_0__4__6 ;
    output FilterDout_0__4__5 ;
    output FilterDout_0__4__4 ;
    output FilterDout_0__4__3 ;
    output FilterDout_0__4__2 ;
    output FilterDout_0__4__1 ;
    output FilterDout_0__4__0 ;
    output FilterDout_1__0__7 ;
    output FilterDout_1__0__6 ;
    output FilterDout_1__0__5 ;
    output FilterDout_1__0__4 ;
    output FilterDout_1__0__3 ;
    output FilterDout_1__0__2 ;
    output FilterDout_1__0__1 ;
    output FilterDout_1__0__0 ;
    output FilterDout_1__1__7 ;
    output FilterDout_1__1__6 ;
    output FilterDout_1__1__5 ;
    output FilterDout_1__1__4 ;
    output FilterDout_1__1__3 ;
    output FilterDout_1__1__2 ;
    output FilterDout_1__1__1 ;
    output FilterDout_1__1__0 ;
    output FilterDout_1__2__7 ;
    output FilterDout_1__2__6 ;
    output FilterDout_1__2__5 ;
    output FilterDout_1__2__4 ;
    output FilterDout_1__2__3 ;
    output FilterDout_1__2__2 ;
    output FilterDout_1__2__1 ;
    output FilterDout_1__2__0 ;
    output FilterDout_1__3__7 ;
    output FilterDout_1__3__6 ;
    output FilterDout_1__3__5 ;
    output FilterDout_1__3__4 ;
    output FilterDout_1__3__3 ;
    output FilterDout_1__3__2 ;
    output FilterDout_1__3__1 ;
    output FilterDout_1__3__0 ;
    output FilterDout_1__4__7 ;
    output FilterDout_1__4__6 ;
    output FilterDout_1__4__5 ;
    output FilterDout_1__4__4 ;
    output FilterDout_1__4__3 ;
    output FilterDout_1__4__2 ;
    output FilterDout_1__4__1 ;
    output FilterDout_1__4__0 ;
    output FilterDout_2__0__7 ;
    output FilterDout_2__0__6 ;
    output FilterDout_2__0__5 ;
    output FilterDout_2__0__4 ;
    output FilterDout_2__0__3 ;
    output FilterDout_2__0__2 ;
    output FilterDout_2__0__1 ;
    output FilterDout_2__0__0 ;
    output FilterDout_2__1__7 ;
    output FilterDout_2__1__6 ;
    output FilterDout_2__1__5 ;
    output FilterDout_2__1__4 ;
    output FilterDout_2__1__3 ;
    output FilterDout_2__1__2 ;
    output FilterDout_2__1__1 ;
    output FilterDout_2__1__0 ;
    output FilterDout_2__2__7 ;
    output FilterDout_2__2__6 ;
    output FilterDout_2__2__5 ;
    output FilterDout_2__2__4 ;
    output FilterDout_2__2__3 ;
    output FilterDout_2__2__2 ;
    output FilterDout_2__2__1 ;
    output FilterDout_2__2__0 ;
    output FilterDout_2__3__7 ;
    output FilterDout_2__3__6 ;
    output FilterDout_2__3__5 ;
    output FilterDout_2__3__4 ;
    output FilterDout_2__3__3 ;
    output FilterDout_2__3__2 ;
    output FilterDout_2__3__1 ;
    output FilterDout_2__3__0 ;
    output FilterDout_2__4__7 ;
    output FilterDout_2__4__6 ;
    output FilterDout_2__4__5 ;
    output FilterDout_2__4__4 ;
    output FilterDout_2__4__3 ;
    output FilterDout_2__4__2 ;
    output FilterDout_2__4__1 ;
    output FilterDout_2__4__0 ;
    output FilterDout_3__0__7 ;
    output FilterDout_3__0__6 ;
    output FilterDout_3__0__5 ;
    output FilterDout_3__0__4 ;
    output FilterDout_3__0__3 ;
    output FilterDout_3__0__2 ;
    output FilterDout_3__0__1 ;
    output FilterDout_3__0__0 ;
    output FilterDout_3__1__7 ;
    output FilterDout_3__1__6 ;
    output FilterDout_3__1__5 ;
    output FilterDout_3__1__4 ;
    output FilterDout_3__1__3 ;
    output FilterDout_3__1__2 ;
    output FilterDout_3__1__1 ;
    output FilterDout_3__1__0 ;
    output FilterDout_3__2__7 ;
    output FilterDout_3__2__6 ;
    output FilterDout_3__2__5 ;
    output FilterDout_3__2__4 ;
    output FilterDout_3__2__3 ;
    output FilterDout_3__2__2 ;
    output FilterDout_3__2__1 ;
    output FilterDout_3__2__0 ;
    output FilterDout_3__3__7 ;
    output FilterDout_3__3__6 ;
    output FilterDout_3__3__5 ;
    output FilterDout_3__3__4 ;
    output FilterDout_3__3__3 ;
    output FilterDout_3__3__2 ;
    output FilterDout_3__3__1 ;
    output FilterDout_3__3__0 ;
    output FilterDout_3__4__7 ;
    output FilterDout_3__4__6 ;
    output FilterDout_3__4__5 ;
    output FilterDout_3__4__4 ;
    output FilterDout_3__4__3 ;
    output FilterDout_3__4__2 ;
    output FilterDout_3__4__1 ;
    output FilterDout_3__4__0 ;
    output FilterDout_4__0__7 ;
    output FilterDout_4__0__6 ;
    output FilterDout_4__0__5 ;
    output FilterDout_4__0__4 ;
    output FilterDout_4__0__3 ;
    output FilterDout_4__0__2 ;
    output FilterDout_4__0__1 ;
    output FilterDout_4__0__0 ;
    output FilterDout_4__1__7 ;
    output FilterDout_4__1__6 ;
    output FilterDout_4__1__5 ;
    output FilterDout_4__1__4 ;
    output FilterDout_4__1__3 ;
    output FilterDout_4__1__2 ;
    output FilterDout_4__1__1 ;
    output FilterDout_4__1__0 ;
    output FilterDout_4__2__7 ;
    output FilterDout_4__2__6 ;
    output FilterDout_4__2__5 ;
    output FilterDout_4__2__4 ;
    output FilterDout_4__2__3 ;
    output FilterDout_4__2__2 ;
    output FilterDout_4__2__1 ;
    output FilterDout_4__2__0 ;
    output FilterDout_4__3__7 ;
    output FilterDout_4__3__6 ;
    output FilterDout_4__3__5 ;
    output FilterDout_4__3__4 ;
    output FilterDout_4__3__3 ;
    output FilterDout_4__3__2 ;
    output FilterDout_4__3__1 ;
    output FilterDout_4__3__0 ;
    output FilterDout_4__4__7 ;
    output FilterDout_4__4__6 ;
    output FilterDout_4__4__5 ;
    output FilterDout_4__4__4 ;
    output FilterDout_4__4__3 ;
    output FilterDout_4__4__2 ;
    output FilterDout_4__4__1 ;
    output FilterDout_4__4__0 ;
    output WindowDout_0__0__7 ;
    output WindowDout_0__0__6 ;
    output WindowDout_0__0__5 ;
    output WindowDout_0__0__4 ;
    output WindowDout_0__0__3 ;
    output WindowDout_0__0__2 ;
    output WindowDout_0__0__1 ;
    output WindowDout_0__0__0 ;
    output WindowDout_0__1__7 ;
    output WindowDout_0__1__6 ;
    output WindowDout_0__1__5 ;
    output WindowDout_0__1__4 ;
    output WindowDout_0__1__3 ;
    output WindowDout_0__1__2 ;
    output WindowDout_0__1__1 ;
    output WindowDout_0__1__0 ;
    output WindowDout_0__2__7 ;
    output WindowDout_0__2__6 ;
    output WindowDout_0__2__5 ;
    output WindowDout_0__2__4 ;
    output WindowDout_0__2__3 ;
    output WindowDout_0__2__2 ;
    output WindowDout_0__2__1 ;
    output WindowDout_0__2__0 ;
    output WindowDout_0__3__7 ;
    output WindowDout_0__3__6 ;
    output WindowDout_0__3__5 ;
    output WindowDout_0__3__4 ;
    output WindowDout_0__3__3 ;
    output WindowDout_0__3__2 ;
    output WindowDout_0__3__1 ;
    output WindowDout_0__3__0 ;
    output WindowDout_0__4__7 ;
    output WindowDout_0__4__6 ;
    output WindowDout_0__4__5 ;
    output WindowDout_0__4__4 ;
    output WindowDout_0__4__3 ;
    output WindowDout_0__4__2 ;
    output WindowDout_0__4__1 ;
    output WindowDout_0__4__0 ;
    output WindowDout_1__0__7 ;
    output WindowDout_1__0__6 ;
    output WindowDout_1__0__5 ;
    output WindowDout_1__0__4 ;
    output WindowDout_1__0__3 ;
    output WindowDout_1__0__2 ;
    output WindowDout_1__0__1 ;
    output WindowDout_1__0__0 ;
    output WindowDout_1__1__7 ;
    output WindowDout_1__1__6 ;
    output WindowDout_1__1__5 ;
    output WindowDout_1__1__4 ;
    output WindowDout_1__1__3 ;
    output WindowDout_1__1__2 ;
    output WindowDout_1__1__1 ;
    output WindowDout_1__1__0 ;
    output WindowDout_1__2__7 ;
    output WindowDout_1__2__6 ;
    output WindowDout_1__2__5 ;
    output WindowDout_1__2__4 ;
    output WindowDout_1__2__3 ;
    output WindowDout_1__2__2 ;
    output WindowDout_1__2__1 ;
    output WindowDout_1__2__0 ;
    output WindowDout_1__3__7 ;
    output WindowDout_1__3__6 ;
    output WindowDout_1__3__5 ;
    output WindowDout_1__3__4 ;
    output WindowDout_1__3__3 ;
    output WindowDout_1__3__2 ;
    output WindowDout_1__3__1 ;
    output WindowDout_1__3__0 ;
    output WindowDout_1__4__7 ;
    output WindowDout_1__4__6 ;
    output WindowDout_1__4__5 ;
    output WindowDout_1__4__4 ;
    output WindowDout_1__4__3 ;
    output WindowDout_1__4__2 ;
    output WindowDout_1__4__1 ;
    output WindowDout_1__4__0 ;
    output WindowDout_2__0__7 ;
    output WindowDout_2__0__6 ;
    output WindowDout_2__0__5 ;
    output WindowDout_2__0__4 ;
    output WindowDout_2__0__3 ;
    output WindowDout_2__0__2 ;
    output WindowDout_2__0__1 ;
    output WindowDout_2__0__0 ;
    output WindowDout_2__1__7 ;
    output WindowDout_2__1__6 ;
    output WindowDout_2__1__5 ;
    output WindowDout_2__1__4 ;
    output WindowDout_2__1__3 ;
    output WindowDout_2__1__2 ;
    output WindowDout_2__1__1 ;
    output WindowDout_2__1__0 ;
    output WindowDout_2__2__7 ;
    output WindowDout_2__2__6 ;
    output WindowDout_2__2__5 ;
    output WindowDout_2__2__4 ;
    output WindowDout_2__2__3 ;
    output WindowDout_2__2__2 ;
    output WindowDout_2__2__1 ;
    output WindowDout_2__2__0 ;
    output WindowDout_2__3__7 ;
    output WindowDout_2__3__6 ;
    output WindowDout_2__3__5 ;
    output WindowDout_2__3__4 ;
    output WindowDout_2__3__3 ;
    output WindowDout_2__3__2 ;
    output WindowDout_2__3__1 ;
    output WindowDout_2__3__0 ;
    output WindowDout_2__4__7 ;
    output WindowDout_2__4__6 ;
    output WindowDout_2__4__5 ;
    output WindowDout_2__4__4 ;
    output WindowDout_2__4__3 ;
    output WindowDout_2__4__2 ;
    output WindowDout_2__4__1 ;
    output WindowDout_2__4__0 ;
    output WindowDout_3__0__7 ;
    output WindowDout_3__0__6 ;
    output WindowDout_3__0__5 ;
    output WindowDout_3__0__4 ;
    output WindowDout_3__0__3 ;
    output WindowDout_3__0__2 ;
    output WindowDout_3__0__1 ;
    output WindowDout_3__0__0 ;
    output WindowDout_3__1__7 ;
    output WindowDout_3__1__6 ;
    output WindowDout_3__1__5 ;
    output WindowDout_3__1__4 ;
    output WindowDout_3__1__3 ;
    output WindowDout_3__1__2 ;
    output WindowDout_3__1__1 ;
    output WindowDout_3__1__0 ;
    output WindowDout_3__2__7 ;
    output WindowDout_3__2__6 ;
    output WindowDout_3__2__5 ;
    output WindowDout_3__2__4 ;
    output WindowDout_3__2__3 ;
    output WindowDout_3__2__2 ;
    output WindowDout_3__2__1 ;
    output WindowDout_3__2__0 ;
    output WindowDout_3__3__7 ;
    output WindowDout_3__3__6 ;
    output WindowDout_3__3__5 ;
    output WindowDout_3__3__4 ;
    output WindowDout_3__3__3 ;
    output WindowDout_3__3__2 ;
    output WindowDout_3__3__1 ;
    output WindowDout_3__3__0 ;
    output WindowDout_3__4__7 ;
    output WindowDout_3__4__6 ;
    output WindowDout_3__4__5 ;
    output WindowDout_3__4__4 ;
    output WindowDout_3__4__3 ;
    output WindowDout_3__4__2 ;
    output WindowDout_3__4__1 ;
    output WindowDout_3__4__0 ;
    output WindowDout_4__0__7 ;
    output WindowDout_4__0__6 ;
    output WindowDout_4__0__5 ;
    output WindowDout_4__0__4 ;
    output WindowDout_4__0__3 ;
    output WindowDout_4__0__2 ;
    output WindowDout_4__0__1 ;
    output WindowDout_4__0__0 ;
    output WindowDout_4__1__7 ;
    output WindowDout_4__1__6 ;
    output WindowDout_4__1__5 ;
    output WindowDout_4__1__4 ;
    output WindowDout_4__1__3 ;
    output WindowDout_4__1__2 ;
    output WindowDout_4__1__1 ;
    output WindowDout_4__1__0 ;
    output WindowDout_4__2__7 ;
    output WindowDout_4__2__6 ;
    output WindowDout_4__2__5 ;
    output WindowDout_4__2__4 ;
    output WindowDout_4__2__3 ;
    output WindowDout_4__2__2 ;
    output WindowDout_4__2__1 ;
    output WindowDout_4__2__0 ;
    output WindowDout_4__3__7 ;
    output WindowDout_4__3__6 ;
    output WindowDout_4__3__5 ;
    output WindowDout_4__3__4 ;
    output WindowDout_4__3__3 ;
    output WindowDout_4__3__2 ;
    output WindowDout_4__3__1 ;
    output WindowDout_4__3__0 ;
    output WindowDout_4__4__7 ;
    output WindowDout_4__4__6 ;
    output WindowDout_4__4__5 ;
    output WindowDout_4__4__4 ;
    output WindowDout_4__4__3 ;
    output WindowDout_4__4__2 ;
    output WindowDout_4__4__1 ;
    output WindowDout_4__4__0 ;
    input ResultWR ;
    input [7:0]ResultDin ;
    output [7:0]ResultDout ;

    wire nx84, nx88, nx98, nx108, nx118, nx128, nx138, nx148, nx158, nx168, 
         nx220, nx230, nx240, nx250, nx260, nx270, nx280, nx290, nx1931, nx1941, 
         nx1951, nx1961, nx1971, nx1981, nx1991, nx2001, nx2011, nx2021, nx2031, 
         nx2041, nx2051, nx2061, nx2071, nx2081, nx2091, nx2101, nx2111, nx2121, 
         nx2131, nx2141, nx2151, nx2161, nx2171, nx2181, nx2191, nx2201, nx2211, 
         nx2221, nx2231, nx2241, nx2251, nx2261, nx2271, nx2281, nx2291, nx2301, 
         nx2311, nx2321, nx2331, nx2341, nx2351, nx2361, nx2371, nx2381, nx2391, 
         nx2401, nx2411, nx2421, nx2431, nx2441, nx2451, nx2461, nx2471, nx2481, 
         nx2491, nx2501, nx2511, nx2521, nx2531, nx2541, nx2551, nx2561, nx2571, 
         nx2581, nx2591, nx2601, nx2611, nx2621, nx2631, nx2641, nx2651, nx2661, 
         nx2671, nx2681, nx2691, nx2701, nx2711, nx2721, nx2731, nx2741, nx2751, 
         nx2761, nx2771, nx2781, nx2791, nx2801, nx2811, nx2821, nx2831, nx2841, 
         nx2851, nx2861, nx2871, nx2881, nx2891, nx2901, nx2911, nx2921, nx2931, 
         nx2941, nx2951, nx2961, nx2971, nx2981, nx2991, nx3001, nx3011, nx3021, 
         nx3031, nx3041, nx3051, nx3061, nx3071, nx3081, nx3091, nx3101, nx3111, 
         nx3121, nx3131, nx3141, nx3151, nx3161, nx3171, nx3181, nx3191, nx3201, 
         nx3211, nx3221, nx3231, nx3241, nx3251, nx3261, nx3271, nx3281, nx3291, 
         nx3301, nx3311, nx3321, nx3331, nx3341, nx3351, nx3361, nx3371, nx3381, 
         nx3391, nx3401, nx3411, nx3421, nx3431, nx3441, nx3451, nx3461, nx3471, 
         nx3481, nx3491, nx3501, nx3511, nx3521, nx3531, nx3541, nx3551, nx3561, 
         nx3571, nx3581, nx3591, nx3601, nx3611, nx3621, nx3631, nx3641, nx3651, 
         nx3661, nx3671, nx3681, nx3691, nx3701, nx3711, nx3721, nx3731, nx3741, 
         nx3751, nx3761, nx3771, nx3781, nx3791, nx3801, nx3811, nx3821, nx3831, 
         nx3841, nx3851, nx3861, nx3871, nx3881, nx3891, nx3901, nx3911, nx3921, 
         nx3931, nx3941, nx3951, nx3961, nx3971, nx3981, nx3991, nx4001, nx4011, 
         nx4021, nx4031, nx4041, nx4051, nx4061, nx4071, nx4081, nx4091, nx4101, 
         nx4111, nx4121, nx4131, nx4141, nx4151, nx4161, nx4171, nx4181, nx4191, 
         nx4201, nx4211, nx4221, nx4231, nx4241, nx4251, nx4261, nx4271, nx4281, 
         nx4291, nx4301, nx4311, nx4321, nx4331, nx4341, nx4351, nx4361, nx4371, 
         nx4381, nx4391, nx4401, nx4411, nx4421, nx4431, nx4441, nx4451, nx4461, 
         nx4471, nx4481, nx4491, nx4501, nx4511, nx4521, nx4531, nx4541, nx4551, 
         nx4561, nx4571, nx4581, nx4591, nx4601, nx4611, nx4621, nx4631, nx4641, 
         nx4651, nx4661, nx4671, nx4681, nx4691, nx4701, nx4711, nx4721, nx4731, 
         nx4741, nx4751, nx4761, nx4771, nx4781, nx4791, nx4801, nx4811, nx4821, 
         nx4831, nx4841, nx4851, nx4861, nx4871, nx4881, nx4891, nx4901, nx4911, 
         nx4921, nx4931, nx4941, nx4951, nx4961, nx4971, nx4981, nx4991, nx5001, 
         nx5011, nx5021, nx5031, nx5041, nx5051, nx5061, nx5071, nx5081, nx5091, 
         nx5101, nx5111, nx5121, nx5131, nx5141, nx5151, nx5161, nx5171, nx5181, 
         nx5191, nx5201, nx5211, nx5221, nx5231, nx5241, nx5251, nx5261, nx5271, 
         nx5281, nx5291, nx5301, nx5311, nx5321, nx5331, nx5341, nx5351, nx5361, 
         nx5371, nx5381, nx5391, nx5401, nx5411, nx5421, nx5431, nx5441, nx5451, 
         nx5461, nx5471, nx5481, nx5491, nx5501, nx5511, nx5521, nx5531, nx5541, 
         nx5551, nx5561, nx5571, nx5581, nx5591, nx5601, nx5611, nx5621, nx5631, 
         nx5641, nx5651, nx5661, nx5671, nx5681, nx5691, nx5701, nx5711, nx5721, 
         nx5731, nx5741, nx5751, nx5761, nx5771, nx5781, nx5791, nx5801, nx5811, 
         nx5821, nx5831, nx5841, nx5851, nx5861, nx5871, nx5881, nx5891, nx5901, 
         nx5911, nx5921, nx5931, nx5941, nx5951, nx5961, nx5971, nx5981, nx5991, 
         nx6001, nx6015, nx6042, nx6107, nx6181, nx6184, nx6188, nx6190, nx6194, 
         nx6196, nx6200, nx6202, nx6206, nx6208, nx6212, nx6214, nx6218, nx6220, 
         nx6224, nx6226, nx6230, nx6232, nx6236, nx6238, nx6242, nx6244, nx6248, 
         nx6250, nx6254, nx6256, nx6260, nx6262, nx6266, nx6268, nx6272, nx6274, 
         nx6350, nx6352, nx6356, nx6358, nx6362, nx6364, nx6368, nx6370, nx6374, 
         nx6376, nx6380, nx6382, nx6386, nx6388, nx6392, nx6394, nx6398, nx6400, 
         nx6404, nx6406, nx6410, nx6412, nx6416, nx6418, nx6422, nx6424, nx6428, 
         nx6430, nx6434, nx6436, nx6440, nx6442, nx6518, nx6520, nx6524, nx6526, 
         nx6530, nx6532, nx6536, nx6538, nx6542, nx6544, nx6548, nx6550, nx6554, 
         nx6556, nx6560, nx6562, nx6566, nx6568, nx6572, nx6574, nx6578, nx6580, 
         nx6584, nx6586, nx6590, nx6592, nx6596, nx6598, nx6602, nx6604, nx6608, 
         nx6610, nx6614, nx6616, nx6620, nx6622, nx6626, nx6628, nx6632, nx6634, 
         nx6638, nx6640, nx6644, nx6646, nx6650, nx6652, nx6656, nx6658, nx6662, 
         nx6664, nx6668, nx6670, nx6674, nx6676, nx6680, nx6682, nx6686, nx6688, 
         nx6692, nx6694, nx6698, nx6700, nx6704, nx6706, nx6710, nx6712, nx6716, 
         nx6718, nx6722, nx6724, nx6728, nx6730, nx6734, nx6736, nx6740, nx6742, 
         nx6746, nx6748, nx6752, nx6754, nx6758, nx6760, nx6764, nx6766, nx6770, 
         nx6772, nx6776, nx6778, nx6782, nx6784, nx6788, nx6790, nx6794, nx6796, 
         nx6800, nx6802, nx6806, nx6808, nx6812, nx6814, nx6818, nx6820, nx6824, 
         nx6826, nx6830, nx6832, nx6836, nx6838, nx6842, nx6844, nx6848, nx6850, 
         nx6854, nx6856, nx6860, nx6862, nx6866, nx6868, nx6872, nx6874, nx6878, 
         nx6880, nx6884, nx6886, nx6890, nx6892, nx6896, nx6898, nx6902, nx6904, 
         nx6908, nx6910, nx6914, nx6916, nx6920, nx6922, nx6926, nx6928, nx6932, 
         nx6934, nx6938, nx6940, nx6944, nx6946, nx6950, nx6952, nx6956, nx6958, 
         nx6962, nx6964, nx6968, nx6970, nx6974, nx6976, nx6980, nx6982, nx6986, 
         nx6988, nx6992, nx6994, nx6998, nx7048, nx7122, nx7125, nx7129, nx7131, 
         nx7135, nx7137, nx7141, nx7143, nx7147, nx7149, nx7153, nx7155, nx7159, 
         nx7161, nx7165, nx7167, nx7171, nx7173, nx7177, nx7179, nx7183, nx7185, 
         nx7189, nx7191, nx7195, nx7197, nx7201, nx7203, nx7207, nx7209, nx7213, 
         nx7215, nx7291, nx7293, nx7297, nx7299, nx7303, nx7305, nx7309, nx7311, 
         nx7315, nx7317, nx7321, nx7323, nx7327, nx7329, nx7333, nx7335, nx7339, 
         nx7341, nx7345, nx7347, nx7351, nx7353, nx7357, nx7359, nx7363, nx7365, 
         nx7369, nx7371, nx7375, nx7377, nx7381, nx7383, nx7459, nx7461, nx7465, 
         nx7467, nx7471, nx7473, nx7477, nx7479, nx7483, nx7485, nx7489, nx7491, 
         nx7495, nx7497, nx7501, nx7503, nx7507, nx7509, nx7513, nx7515, nx7519, 
         nx7521, nx7525, nx7527, nx7531, nx7533, nx7537, nx7539, nx7543, nx7545, 
         nx7549, nx7551, nx7555, nx7557, nx7561, nx7563, nx7567, nx7569, nx7573, 
         nx7575, nx7579, nx7581, nx7585, nx7587, nx7591, nx7593, nx7597, nx7599, 
         nx7603, nx7605, nx7609, nx7611, nx7615, nx7617, nx7621, nx7623, nx7627, 
         nx7629, nx7633, nx7635, nx7639, nx7641, nx7645, nx7647, nx7651, nx7653, 
         nx7657, nx7659, nx7663, nx7665, nx7669, nx7671, nx7675, nx7677, nx7681, 
         nx7683, nx7687, nx7689, nx7693, nx7695, nx7699, nx7701, nx7705, nx7707, 
         nx7711, nx7713, nx7717, nx7719, nx7723, nx7725, nx7729, nx7731, nx7735, 
         nx7737, nx7741, nx7743, nx7747, nx7749, nx7753, nx7755, nx7759, nx7761, 
         nx7765, nx7767, nx7771, nx7773, nx7777, nx7779, nx7783, nx7785, nx7789, 
         nx7791, nx7795, nx7797, nx7801, nx7803, nx7807, nx7809, nx7813, nx7815, 
         nx7819, nx7821, nx7825, nx7827, nx7831, nx7833, nx7837, nx7839, nx7843, 
         nx7845, nx7849, nx7851, nx7855, nx7857, nx7861, nx7863, nx7867, nx7869, 
         nx7873, nx7875, nx7879, nx7881, nx7885, nx7887, nx7891, nx7893, nx7897, 
         nx7899, nx7903, nx7905, nx7909, nx7911, nx7915, nx7917, nx7921, nx7923, 
         nx7927, nx7929, nx7933, nx7935, nx7942, nx7944, nx7946, nx7948, nx7950, 
         nx7952, nx7954, nx7956, nx7958, nx7960, nx7962, nx7964, nx7966, nx7968, 
         nx7970, nx7972, nx7974, nx7976, nx7978, nx7980, nx7982, nx7984, nx7986, 
         nx7988, nx7990, nx7992, nx7994, nx7996, nx7998, nx8000, nx8002, nx8004, 
         nx8006, nx8008, nx8010, nx8012, nx8014, nx8016, nx8018, nx8020, nx8022, 
         nx8024, nx8026, nx8028, nx8030, nx8032, nx8034, nx8036, nx8038, nx8040, 
         nx8042, nx8044, nx8046, nx8048, nx8050, nx8052, nx8054, nx8056, nx8058, 
         nx8060, nx8062, nx8064, nx8066, nx8068, nx8070, nx8072, nx8074, nx8076, 
         nx8078, nx8080, nx8082, nx8084, nx8086, nx8088, nx8090, nx8094, nx8096, 
         nx8098, nx8100, nx8106, nx8108, nx8110, nx8112, nx8124, nx8126, nx8128, 
         nx8130, nx8132, nx8134, nx8136, nx8138, nx8140, nx8142, nx8146, nx8148, 
         nx8150, nx8152, nx8154, nx8158, nx8160, nx8162, nx8164, nx8182, nx8184, 
         nx8186, nx8188, nx8190, nx8194, nx8196, nx8198, nx8200, nx8202, nx8204, 
         nx8206, nx8208, nx8210, nx8212, nx8214, nx8220, nx8222, nx8224, nx8226, 
         nx8228, nx8232, nx8234, nx8236, nx8238, nx8240, nx8242, nx8244, nx8246, 
         nx8248, nx8250, nx8252, nx8254, nx8256, nx8258, nx8260, nx8270, nx8272, 
         nx8274, nx8276, nx8278, nx8280, nx8282, nx8284, nx8286, nx8288, nx8290, 
         nx8292, nx8294, nx8296, nx8298, nx8300, nx8302, nx8304, nx8306, nx8308, 
         nx8310, nx8312, nx8314, nx8316, nx8318, nx8320, nx8322, nx8324, nx8326, 
         nx8328, nx8334, nx8336;
    wire [183:0] \$dummy ;




    dff RESULT_REG_reg_Dout_0 (.Q (ResultDout[0]), .QB (\$dummy [0]), .D (nx1931
        ), .CLK (CLK)) ;
    ao32 ix1932 (.Y (nx1931), .A0 (ResultDin[0]), .A1 (nx8070), .A2 (ResultWR), 
         .B0 (ResultDout[0]), .B1 (nx6015)) ;
    nor02_2x ix6016 (.Y (nx6015), .A0 (RST), .A1 (ResultWR)) ;
    dff RESULT_REG_reg_Dout_1 (.Q (ResultDout[1]), .QB (\$dummy [1]), .D (nx1941
        ), .CLK (CLK)) ;
    ao32 ix1942 (.Y (nx1941), .A0 (ResultDin[1]), .A1 (nx8070), .A2 (ResultWR), 
         .B0 (ResultDout[1]), .B1 (nx6015)) ;
    dff RESULT_REG_reg_Dout_2 (.Q (ResultDout[2]), .QB (\$dummy [2]), .D (nx1951
        ), .CLK (CLK)) ;
    ao32 ix1952 (.Y (nx1951), .A0 (ResultDin[2]), .A1 (nx8070), .A2 (ResultWR), 
         .B0 (ResultDout[2]), .B1 (nx6015)) ;
    dff RESULT_REG_reg_Dout_3 (.Q (ResultDout[3]), .QB (\$dummy [3]), .D (nx1961
        ), .CLK (CLK)) ;
    ao32 ix1962 (.Y (nx1961), .A0 (ResultDin[3]), .A1 (nx8070), .A2 (ResultWR), 
         .B0 (ResultDout[3]), .B1 (nx6015)) ;
    dff RESULT_REG_reg_Dout_4 (.Q (ResultDout[4]), .QB (\$dummy [4]), .D (nx1971
        ), .CLK (CLK)) ;
    ao32 ix1972 (.Y (nx1971), .A0 (ResultDin[4]), .A1 (nx8070), .A2 (ResultWR), 
         .B0 (ResultDout[4]), .B1 (nx6015)) ;
    dff RESULT_REG_reg_Dout_5 (.Q (ResultDout[5]), .QB (\$dummy [5]), .D (nx1981
        ), .CLK (CLK)) ;
    ao32 ix1982 (.Y (nx1981), .A0 (ResultDin[5]), .A1 (nx8070), .A2 (ResultWR), 
         .B0 (ResultDout[5]), .B1 (nx6015)) ;
    dff RESULT_REG_reg_Dout_6 (.Q (ResultDout[6]), .QB (\$dummy [6]), .D (nx1991
        ), .CLK (CLK)) ;
    ao32 ix1992 (.Y (nx1991), .A0 (ResultDin[6]), .A1 (nx8070), .A2 (ResultWR), 
         .B0 (ResultDout[6]), .B1 (nx6015)) ;
    dff RESULT_REG_reg_Dout_7 (.Q (ResultDout[7]), .QB (\$dummy [7]), .D (nx2001
        ), .CLK (CLK)) ;
    ao32 ix2002 (.Y (nx2001), .A0 (ResultDin[7]), .A1 (nx8072), .A2 (ResultWR), 
         .B0 (ResultDout[7]), .B1 (nx6015)) ;
    dff L0_4_L1_4_Wij_reg_Dout_0 (.Q (WindowDout_4__4__0), .QB (\$dummy [8]), .D (
        nx2011), .CLK (CLK)) ;
    nor02ii ix89 (.Y (nx88), .A0 (RST), .A1 (Din[32])) ;
    aoi21 ix6043 (.Y (nx6042), .A0 (WindowWR), .A1 (FilterSize), .B0 (RST)) ;
    dff L0_4_L1_4_Wij_reg_Dout_1 (.Q (WindowDout_4__4__1), .QB (\$dummy [9]), .D (
        nx2021), .CLK (CLK)) ;
    nor02ii ix99 (.Y (nx98), .A0 (RST), .A1 (Din[33])) ;
    dff L0_4_L1_4_Wij_reg_Dout_2 (.Q (WindowDout_4__4__2), .QB (\$dummy [10]), .D (
        nx2031), .CLK (CLK)) ;
    nor02ii ix109 (.Y (nx108), .A0 (RST), .A1 (Din[34])) ;
    dff L0_4_L1_4_Wij_reg_Dout_3 (.Q (WindowDout_4__4__3), .QB (\$dummy [11]), .D (
        nx2041), .CLK (CLK)) ;
    nor02ii ix119 (.Y (nx118), .A0 (RST), .A1 (Din[35])) ;
    dff L0_4_L1_4_Wij_reg_Dout_4 (.Q (WindowDout_4__4__4), .QB (\$dummy [12]), .D (
        nx2051), .CLK (CLK)) ;
    nor02ii ix129 (.Y (nx128), .A0 (RST), .A1 (Din[36])) ;
    dff L0_4_L1_4_Wij_reg_Dout_5 (.Q (WindowDout_4__4__5), .QB (\$dummy [13]), .D (
        nx2061), .CLK (CLK)) ;
    nor02ii ix139 (.Y (nx138), .A0 (RST), .A1 (Din[37])) ;
    dff L0_4_L1_4_Wij_reg_Dout_6 (.Q (WindowDout_4__4__6), .QB (\$dummy [14]), .D (
        nx2071), .CLK (CLK)) ;
    nor02ii ix149 (.Y (nx148), .A0 (RST), .A1 (Din[38])) ;
    dff L0_4_L1_4_Wij_reg_Dout_7 (.Q (WindowDout_4__4__7), .QB (\$dummy [15]), .D (
        nx2081), .CLK (CLK)) ;
    nor02ii ix159 (.Y (nx158), .A0 (RST), .A1 (Din[39])) ;
    dff L0_4_L1_3_Wij_reg_Dout_0 (.Q (WindowDout_4__3__0), .QB (\$dummy [16]), .D (
        nx2171), .CLK (CLK)) ;
    nor02ii ix221 (.Y (nx220), .A0 (RST), .A1 (Din[24])) ;
    dff L0_4_L1_3_Wij_reg_Dout_1 (.Q (WindowDout_4__3__1), .QB (\$dummy [17]), .D (
        nx2181), .CLK (CLK)) ;
    nor02ii ix231 (.Y (nx230), .A0 (RST), .A1 (Din[25])) ;
    dff L0_4_L1_3_Wij_reg_Dout_2 (.Q (WindowDout_4__3__2), .QB (\$dummy [18]), .D (
        nx2191), .CLK (CLK)) ;
    nor02ii ix241 (.Y (nx240), .A0 (RST), .A1 (Din[26])) ;
    dff L0_4_L1_3_Wij_reg_Dout_3 (.Q (WindowDout_4__3__3), .QB (\$dummy [19]), .D (
        nx2201), .CLK (CLK)) ;
    nor02ii ix251 (.Y (nx250), .A0 (RST), .A1 (Din[27])) ;
    dff L0_4_L1_3_Wij_reg_Dout_4 (.Q (WindowDout_4__3__4), .QB (\$dummy [20]), .D (
        nx2211), .CLK (CLK)) ;
    nor02ii ix261 (.Y (nx260), .A0 (RST), .A1 (Din[28])) ;
    dff L0_4_L1_3_Wij_reg_Dout_5 (.Q (WindowDout_4__3__5), .QB (\$dummy [21]), .D (
        nx2221), .CLK (CLK)) ;
    nor02ii ix271 (.Y (nx270), .A0 (RST), .A1 (Din[29])) ;
    dff L0_4_L1_3_Wij_reg_Dout_6 (.Q (WindowDout_4__3__6), .QB (\$dummy [22]), .D (
        nx2231), .CLK (CLK)) ;
    nor02ii ix281 (.Y (nx280), .A0 (RST), .A1 (Din[30])) ;
    dff L0_4_L1_3_Wij_reg_Dout_7 (.Q (WindowDout_4__3__7), .QB (\$dummy [23]), .D (
        nx2241), .CLK (CLK)) ;
    nor02ii ix291 (.Y (nx290), .A0 (RST), .A1 (Din[31])) ;
    dff L0_4_L1_2_Wij_reg_Dout_0 (.Q (WindowDout_4__2__0), .QB (\$dummy [24]), .D (
        nx2331), .CLK (CLK)) ;
    ao32 ix2332 (.Y (nx2331), .A0 (Din[16]), .A1 (nx8072), .A2 (WindowWR), .B0 (
         WindowDout_4__2__0), .B1 (nx8194)) ;
    nor02_2x ix6108 (.Y (nx6107), .A0 (WindowWR), .A1 (RST)) ;
    dff L0_4_L1_2_Wij_reg_Dout_1 (.Q (WindowDout_4__2__1), .QB (\$dummy [25]), .D (
        nx2341), .CLK (CLK)) ;
    ao32 ix2342 (.Y (nx2341), .A0 (Din[17]), .A1 (nx8072), .A2 (WindowWR), .B0 (
         WindowDout_4__2__1), .B1 (nx8194)) ;
    dff L0_4_L1_2_Wij_reg_Dout_2 (.Q (WindowDout_4__2__2), .QB (\$dummy [26]), .D (
        nx2351), .CLK (CLK)) ;
    ao32 ix2352 (.Y (nx2351), .A0 (Din[18]), .A1 (nx8072), .A2 (WindowWR), .B0 (
         WindowDout_4__2__2), .B1 (nx8194)) ;
    dff L0_4_L1_2_Wij_reg_Dout_3 (.Q (WindowDout_4__2__3), .QB (\$dummy [27]), .D (
        nx2361), .CLK (CLK)) ;
    ao32 ix2362 (.Y (nx2361), .A0 (Din[19]), .A1 (nx8072), .A2 (WindowWR), .B0 (
         WindowDout_4__2__3), .B1 (nx8194)) ;
    dff L0_4_L1_2_Wij_reg_Dout_4 (.Q (WindowDout_4__2__4), .QB (\$dummy [28]), .D (
        nx2371), .CLK (CLK)) ;
    ao32 ix2372 (.Y (nx2371), .A0 (Din[20]), .A1 (nx8072), .A2 (WindowWR), .B0 (
         WindowDout_4__2__4), .B1 (nx8194)) ;
    dff L0_4_L1_2_Wij_reg_Dout_5 (.Q (WindowDout_4__2__5), .QB (\$dummy [29]), .D (
        nx2381), .CLK (CLK)) ;
    ao32 ix2382 (.Y (nx2381), .A0 (Din[21]), .A1 (nx8072), .A2 (WindowWR), .B0 (
         WindowDout_4__2__5), .B1 (nx8194)) ;
    dff L0_4_L1_2_Wij_reg_Dout_6 (.Q (WindowDout_4__2__6), .QB (\$dummy [30]), .D (
        nx2391), .CLK (CLK)) ;
    ao32 ix2392 (.Y (nx2391), .A0 (Din[22]), .A1 (nx8074), .A2 (WindowWR), .B0 (
         WindowDout_4__2__6), .B1 (nx8194)) ;
    dff L0_4_L1_2_Wij_reg_Dout_7 (.Q (WindowDout_4__2__7), .QB (\$dummy [31]), .D (
        nx2401), .CLK (CLK)) ;
    ao32 ix2402 (.Y (nx2401), .A0 (Din[23]), .A1 (nx8074), .A2 (WindowWR), .B0 (
         WindowDout_4__2__7), .B1 (nx8196)) ;
    dff L0_4_L1_1_Wij_reg_Dout_0 (.Q (WindowDout_4__1__0), .QB (\$dummy [32]), .D (
        nx2491), .CLK (CLK)) ;
    ao32 ix2492 (.Y (nx2491), .A0 (Din[8]), .A1 (nx8074), .A2 (WindowWR), .B0 (
         WindowDout_4__1__0), .B1 (nx8196)) ;
    dff L0_4_L1_1_Wij_reg_Dout_1 (.Q (WindowDout_4__1__1), .QB (\$dummy [33]), .D (
        nx2501), .CLK (CLK)) ;
    ao32 ix2502 (.Y (nx2501), .A0 (Din[9]), .A1 (nx8074), .A2 (WindowWR), .B0 (
         WindowDout_4__1__1), .B1 (nx8196)) ;
    dff L0_4_L1_1_Wij_reg_Dout_2 (.Q (WindowDout_4__1__2), .QB (\$dummy [34]), .D (
        nx2511), .CLK (CLK)) ;
    ao32 ix2512 (.Y (nx2511), .A0 (Din[10]), .A1 (nx8074), .A2 (WindowWR), .B0 (
         WindowDout_4__1__2), .B1 (nx8196)) ;
    dff L0_4_L1_1_Wij_reg_Dout_3 (.Q (WindowDout_4__1__3), .QB (\$dummy [35]), .D (
        nx2521), .CLK (CLK)) ;
    ao32 ix2522 (.Y (nx2521), .A0 (Din[11]), .A1 (nx8074), .A2 (WindowWR), .B0 (
         WindowDout_4__1__3), .B1 (nx8196)) ;
    dff L0_4_L1_1_Wij_reg_Dout_4 (.Q (WindowDout_4__1__4), .QB (\$dummy [36]), .D (
        nx2531), .CLK (CLK)) ;
    ao32 ix2532 (.Y (nx2531), .A0 (Din[12]), .A1 (nx8074), .A2 (WindowWR), .B0 (
         WindowDout_4__1__4), .B1 (nx8196)) ;
    dff L0_4_L1_1_Wij_reg_Dout_5 (.Q (WindowDout_4__1__5), .QB (\$dummy [37]), .D (
        nx2541), .CLK (CLK)) ;
    ao32 ix2542 (.Y (nx2541), .A0 (Din[13]), .A1 (nx8076), .A2 (WindowWR), .B0 (
         WindowDout_4__1__5), .B1 (nx8196)) ;
    dff L0_4_L1_1_Wij_reg_Dout_6 (.Q (WindowDout_4__1__6), .QB (\$dummy [38]), .D (
        nx2551), .CLK (CLK)) ;
    ao32 ix2552 (.Y (nx2551), .A0 (Din[14]), .A1 (nx8076), .A2 (WindowWR), .B0 (
         WindowDout_4__1__6), .B1 (nx8198)) ;
    dff L0_4_L1_1_Wij_reg_Dout_7 (.Q (WindowDout_4__1__7), .QB (\$dummy [39]), .D (
        nx2561), .CLK (CLK)) ;
    ao32 ix2562 (.Y (nx2561), .A0 (Din[15]), .A1 (nx8076), .A2 (WindowWR), .B0 (
         WindowDout_4__1__7), .B1 (nx8198)) ;
    dff L0_4_L1_0_Wij_reg_Dout_0 (.Q (WindowDout_4__0__0), .QB (\$dummy [40]), .D (
        nx2651), .CLK (CLK)) ;
    ao32 ix2652 (.Y (nx2651), .A0 (Din[0]), .A1 (nx8076), .A2 (WindowWR), .B0 (
         WindowDout_4__0__0), .B1 (nx8198)) ;
    dff L0_4_L1_0_Wij_reg_Dout_1 (.Q (WindowDout_4__0__1), .QB (\$dummy [41]), .D (
        nx2661), .CLK (CLK)) ;
    ao32 ix2662 (.Y (nx2661), .A0 (Din[1]), .A1 (nx8076), .A2 (WindowWR), .B0 (
         WindowDout_4__0__1), .B1 (nx8198)) ;
    dff L0_4_L1_0_Wij_reg_Dout_2 (.Q (WindowDout_4__0__2), .QB (\$dummy [42]), .D (
        nx2671), .CLK (CLK)) ;
    ao32 ix2672 (.Y (nx2671), .A0 (Din[2]), .A1 (nx8076), .A2 (WindowWR), .B0 (
         WindowDout_4__0__2), .B1 (nx8198)) ;
    dff L0_4_L1_0_Wij_reg_Dout_3 (.Q (WindowDout_4__0__3), .QB (\$dummy [43]), .D (
        nx2681), .CLK (CLK)) ;
    ao32 ix2682 (.Y (nx2681), .A0 (Din[3]), .A1 (nx8076), .A2 (WindowWR), .B0 (
         WindowDout_4__0__3), .B1 (nx8198)) ;
    dff L0_4_L1_0_Wij_reg_Dout_4 (.Q (WindowDout_4__0__4), .QB (\$dummy [44]), .D (
        nx2691), .CLK (CLK)) ;
    ao32 ix2692 (.Y (nx2691), .A0 (Din[4]), .A1 (nx8078), .A2 (WindowWR), .B0 (
         WindowDout_4__0__4), .B1 (nx8198)) ;
    dff L0_4_L1_0_Wij_reg_Dout_5 (.Q (WindowDout_4__0__5), .QB (\$dummy [45]), .D (
        nx2701), .CLK (CLK)) ;
    ao32 ix2702 (.Y (nx2701), .A0 (Din[5]), .A1 (nx8078), .A2 (WindowWR), .B0 (
         WindowDout_4__0__5), .B1 (nx8200)) ;
    dff L0_4_L1_0_Wij_reg_Dout_6 (.Q (WindowDout_4__0__6), .QB (\$dummy [46]), .D (
        nx2711), .CLK (CLK)) ;
    ao32 ix2712 (.Y (nx2711), .A0 (Din[6]), .A1 (nx8078), .A2 (WindowWR), .B0 (
         WindowDout_4__0__6), .B1 (nx8200)) ;
    dff L0_4_L1_0_Wij_reg_Dout_7 (.Q (WindowDout_4__0__7), .QB (\$dummy [47]), .D (
        nx2721), .CLK (CLK)) ;
    ao32 ix2722 (.Y (nx2721), .A0 (Din[7]), .A1 (nx8078), .A2 (WindowWR), .B0 (
         WindowDout_4__0__7), .B1 (nx8200)) ;
    oai21 ix2812 (.Y (nx2811), .A0 (nx6181), .A1 (nx7942), .B0 (nx6184)) ;
    dff L0_3_L1_4_Wij_reg_Dout_0 (.Q (WindowDout_3__4__0), .QB (nx6181), .D (
        nx2811), .CLK (CLK)) ;
    nand03 ix6185 (.Y (nx6184), .A0 (nx8078), .A1 (WindowDout_4__4__0), .A2 (
           nx7942)) ;
    oai21 ix2822 (.Y (nx2821), .A0 (nx6188), .A1 (nx7942), .B0 (nx6190)) ;
    dff L0_3_L1_4_Wij_reg_Dout_1 (.Q (WindowDout_3__4__1), .QB (nx6188), .D (
        nx2821), .CLK (CLK)) ;
    nand03 ix6191 (.Y (nx6190), .A0 (nx8078), .A1 (WindowDout_4__4__1), .A2 (
           nx7942)) ;
    oai21 ix2832 (.Y (nx2831), .A0 (nx6194), .A1 (nx7942), .B0 (nx6196)) ;
    dff L0_3_L1_4_Wij_reg_Dout_2 (.Q (WindowDout_3__4__2), .QB (nx6194), .D (
        nx2831), .CLK (CLK)) ;
    nand03 ix6197 (.Y (nx6196), .A0 (nx8078), .A1 (WindowDout_4__4__2), .A2 (
           nx7942)) ;
    oai21 ix2842 (.Y (nx2841), .A0 (nx6200), .A1 (nx7942), .B0 (nx6202)) ;
    dff L0_3_L1_4_Wij_reg_Dout_3 (.Q (WindowDout_3__4__3), .QB (nx6200), .D (
        nx2841), .CLK (CLK)) ;
    nand03 ix6203 (.Y (nx6202), .A0 (nx8080), .A1 (WindowDout_4__4__3), .A2 (
           nx7944)) ;
    oai21 ix2852 (.Y (nx2851), .A0 (nx6206), .A1 (nx7944), .B0 (nx6208)) ;
    dff L0_3_L1_4_Wij_reg_Dout_4 (.Q (WindowDout_3__4__4), .QB (nx6206), .D (
        nx2851), .CLK (CLK)) ;
    nand03 ix6209 (.Y (nx6208), .A0 (nx8080), .A1 (WindowDout_4__4__4), .A2 (
           nx7944)) ;
    oai21 ix2862 (.Y (nx2861), .A0 (nx6212), .A1 (nx7944), .B0 (nx6214)) ;
    dff L0_3_L1_4_Wij_reg_Dout_5 (.Q (WindowDout_3__4__5), .QB (nx6212), .D (
        nx2861), .CLK (CLK)) ;
    nand03 ix6215 (.Y (nx6214), .A0 (nx8080), .A1 (WindowDout_4__4__5), .A2 (
           nx7944)) ;
    oai21 ix2872 (.Y (nx2871), .A0 (nx6218), .A1 (nx7944), .B0 (nx6220)) ;
    dff L0_3_L1_4_Wij_reg_Dout_6 (.Q (WindowDout_3__4__6), .QB (nx6218), .D (
        nx2871), .CLK (CLK)) ;
    nand03 ix6221 (.Y (nx6220), .A0 (nx8080), .A1 (WindowDout_4__4__6), .A2 (
           nx7944)) ;
    oai21 ix2882 (.Y (nx2881), .A0 (nx6224), .A1 (nx7946), .B0 (nx6226)) ;
    dff L0_3_L1_4_Wij_reg_Dout_7 (.Q (WindowDout_3__4__7), .QB (nx6224), .D (
        nx2881), .CLK (CLK)) ;
    nand03 ix6227 (.Y (nx6226), .A0 (nx8080), .A1 (WindowDout_4__4__7), .A2 (
           nx7946)) ;
    oai21 ix2972 (.Y (nx2971), .A0 (nx6230), .A1 (nx7946), .B0 (nx6232)) ;
    dff L0_3_L1_3_Wij_reg_Dout_0 (.Q (WindowDout_3__3__0), .QB (nx6230), .D (
        nx2971), .CLK (CLK)) ;
    nand03 ix6233 (.Y (nx6232), .A0 (nx8080), .A1 (WindowDout_4__3__0), .A2 (
           nx7946)) ;
    oai21 ix2982 (.Y (nx2981), .A0 (nx6236), .A1 (nx7946), .B0 (nx6238)) ;
    dff L0_3_L1_3_Wij_reg_Dout_1 (.Q (WindowDout_3__3__1), .QB (nx6236), .D (
        nx2981), .CLK (CLK)) ;
    nand03 ix6239 (.Y (nx6238), .A0 (nx8080), .A1 (WindowDout_4__3__1), .A2 (
           nx7946)) ;
    oai21 ix2992 (.Y (nx2991), .A0 (nx6242), .A1 (nx7946), .B0 (nx6244)) ;
    dff L0_3_L1_3_Wij_reg_Dout_2 (.Q (WindowDout_3__3__2), .QB (nx6242), .D (
        nx2991), .CLK (CLK)) ;
    nand03 ix6245 (.Y (nx6244), .A0 (nx8082), .A1 (WindowDout_4__3__2), .A2 (
           nx7948)) ;
    oai21 ix3002 (.Y (nx3001), .A0 (nx6248), .A1 (nx7948), .B0 (nx6250)) ;
    dff L0_3_L1_3_Wij_reg_Dout_3 (.Q (WindowDout_3__3__3), .QB (nx6248), .D (
        nx3001), .CLK (CLK)) ;
    nand03 ix6251 (.Y (nx6250), .A0 (nx8082), .A1 (WindowDout_4__3__3), .A2 (
           nx7948)) ;
    oai21 ix3012 (.Y (nx3011), .A0 (nx6254), .A1 (nx7948), .B0 (nx6256)) ;
    dff L0_3_L1_3_Wij_reg_Dout_4 (.Q (WindowDout_3__3__4), .QB (nx6254), .D (
        nx3011), .CLK (CLK)) ;
    nand03 ix6257 (.Y (nx6256), .A0 (nx8082), .A1 (WindowDout_4__3__4), .A2 (
           nx7948)) ;
    oai21 ix3022 (.Y (nx3021), .A0 (nx6260), .A1 (nx7948), .B0 (nx6262)) ;
    dff L0_3_L1_3_Wij_reg_Dout_5 (.Q (WindowDout_3__3__5), .QB (nx6260), .D (
        nx3021), .CLK (CLK)) ;
    nand03 ix6263 (.Y (nx6262), .A0 (nx8082), .A1 (WindowDout_4__3__5), .A2 (
           nx7948)) ;
    oai21 ix3032 (.Y (nx3031), .A0 (nx6266), .A1 (nx7950), .B0 (nx6268)) ;
    dff L0_3_L1_3_Wij_reg_Dout_6 (.Q (WindowDout_3__3__6), .QB (nx6266), .D (
        nx3031), .CLK (CLK)) ;
    nand03 ix6269 (.Y (nx6268), .A0 (nx8082), .A1 (WindowDout_4__3__6), .A2 (
           nx7950)) ;
    oai21 ix3042 (.Y (nx3041), .A0 (nx6272), .A1 (nx7950), .B0 (nx6274)) ;
    dff L0_3_L1_3_Wij_reg_Dout_7 (.Q (WindowDout_3__3__7), .QB (nx6272), .D (
        nx3041), .CLK (CLK)) ;
    nand03 ix6275 (.Y (nx6274), .A0 (nx8082), .A1 (WindowDout_4__3__7), .A2 (
           nx7950)) ;
    dff L0_3_L1_2_Wij_reg_Dout_0 (.Q (WindowDout_3__2__0), .QB (\$dummy [48]), .D (
        nx3131), .CLK (CLK)) ;
    ao32 ix3132 (.Y (nx3131), .A0 (nx8082), .A1 (WindowDout_4__2__0), .A2 (
         WindowWR), .B0 (WindowDout_3__2__0), .B1 (nx8200)) ;
    dff L0_3_L1_2_Wij_reg_Dout_1 (.Q (WindowDout_3__2__1), .QB (\$dummy [49]), .D (
        nx3141), .CLK (CLK)) ;
    ao32 ix3142 (.Y (nx3141), .A0 (nx8084), .A1 (WindowDout_4__2__1), .A2 (
         WindowWR), .B0 (WindowDout_3__2__1), .B1 (nx8200)) ;
    dff L0_3_L1_2_Wij_reg_Dout_2 (.Q (WindowDout_3__2__2), .QB (\$dummy [50]), .D (
        nx3151), .CLK (CLK)) ;
    ao32 ix3152 (.Y (nx3151), .A0 (nx8084), .A1 (WindowDout_4__2__2), .A2 (
         WindowWR), .B0 (WindowDout_3__2__2), .B1 (nx8200)) ;
    dff L0_3_L1_2_Wij_reg_Dout_3 (.Q (WindowDout_3__2__3), .QB (\$dummy [51]), .D (
        nx3161), .CLK (CLK)) ;
    ao32 ix3162 (.Y (nx3161), .A0 (nx8084), .A1 (WindowDout_4__2__3), .A2 (
         WindowWR), .B0 (WindowDout_3__2__3), .B1 (nx8200)) ;
    dff L0_3_L1_2_Wij_reg_Dout_4 (.Q (WindowDout_3__2__4), .QB (\$dummy [52]), .D (
        nx3171), .CLK (CLK)) ;
    ao32 ix3172 (.Y (nx3171), .A0 (nx8084), .A1 (WindowDout_4__2__4), .A2 (
         WindowWR), .B0 (WindowDout_3__2__4), .B1 (nx8202)) ;
    dff L0_3_L1_2_Wij_reg_Dout_5 (.Q (WindowDout_3__2__5), .QB (\$dummy [53]), .D (
        nx3181), .CLK (CLK)) ;
    ao32 ix3182 (.Y (nx3181), .A0 (nx8084), .A1 (WindowDout_4__2__5), .A2 (
         WindowWR), .B0 (WindowDout_3__2__5), .B1 (nx8202)) ;
    dff L0_3_L1_2_Wij_reg_Dout_6 (.Q (WindowDout_3__2__6), .QB (\$dummy [54]), .D (
        nx3191), .CLK (CLK)) ;
    ao32 ix3192 (.Y (nx3191), .A0 (nx8084), .A1 (WindowDout_4__2__6), .A2 (
         WindowWR), .B0 (WindowDout_3__2__6), .B1 (nx8202)) ;
    dff L0_3_L1_2_Wij_reg_Dout_7 (.Q (WindowDout_3__2__7), .QB (\$dummy [55]), .D (
        nx3201), .CLK (CLK)) ;
    ao32 ix3202 (.Y (nx3201), .A0 (nx8084), .A1 (WindowDout_4__2__7), .A2 (
         WindowWR), .B0 (WindowDout_3__2__7), .B1 (nx8202)) ;
    dff L0_3_L1_1_Wij_reg_Dout_0 (.Q (WindowDout_3__1__0), .QB (\$dummy [56]), .D (
        nx3291), .CLK (CLK)) ;
    ao32 ix3292 (.Y (nx3291), .A0 (nx8086), .A1 (WindowDout_4__1__0), .A2 (
         WindowWR), .B0 (WindowDout_3__1__0), .B1 (nx8202)) ;
    dff L0_3_L1_1_Wij_reg_Dout_1 (.Q (WindowDout_3__1__1), .QB (\$dummy [57]), .D (
        nx3301), .CLK (CLK)) ;
    ao32 ix3302 (.Y (nx3301), .A0 (nx8086), .A1 (WindowDout_4__1__1), .A2 (
         WindowWR), .B0 (WindowDout_3__1__1), .B1 (nx8202)) ;
    dff L0_3_L1_1_Wij_reg_Dout_2 (.Q (WindowDout_3__1__2), .QB (\$dummy [58]), .D (
        nx3311), .CLK (CLK)) ;
    ao32 ix3312 (.Y (nx3311), .A0 (nx8086), .A1 (WindowDout_4__1__2), .A2 (
         WindowWR), .B0 (WindowDout_3__1__2), .B1 (nx8202)) ;
    dff L0_3_L1_1_Wij_reg_Dout_3 (.Q (WindowDout_3__1__3), .QB (\$dummy [59]), .D (
        nx3321), .CLK (CLK)) ;
    ao32 ix3322 (.Y (nx3321), .A0 (nx8086), .A1 (WindowDout_4__1__3), .A2 (
         WindowWR), .B0 (WindowDout_3__1__3), .B1 (nx8204)) ;
    dff L0_3_L1_1_Wij_reg_Dout_4 (.Q (WindowDout_3__1__4), .QB (\$dummy [60]), .D (
        nx3331), .CLK (CLK)) ;
    ao32 ix3332 (.Y (nx3331), .A0 (nx8086), .A1 (WindowDout_4__1__4), .A2 (
         WindowWR), .B0 (WindowDout_3__1__4), .B1 (nx8204)) ;
    dff L0_3_L1_1_Wij_reg_Dout_5 (.Q (WindowDout_3__1__5), .QB (\$dummy [61]), .D (
        nx3341), .CLK (CLK)) ;
    ao32 ix3342 (.Y (nx3341), .A0 (nx8086), .A1 (WindowDout_4__1__5), .A2 (
         WindowWR), .B0 (WindowDout_3__1__5), .B1 (nx8204)) ;
    dff L0_3_L1_1_Wij_reg_Dout_6 (.Q (WindowDout_3__1__6), .QB (\$dummy [62]), .D (
        nx3351), .CLK (CLK)) ;
    ao32 ix3352 (.Y (nx3351), .A0 (nx8086), .A1 (WindowDout_4__1__6), .A2 (
         WindowWR), .B0 (WindowDout_3__1__6), .B1 (nx8204)) ;
    dff L0_3_L1_1_Wij_reg_Dout_7 (.Q (WindowDout_3__1__7), .QB (\$dummy [63]), .D (
        nx3361), .CLK (CLK)) ;
    ao32 ix3362 (.Y (nx3361), .A0 (nx8088), .A1 (WindowDout_4__1__7), .A2 (
         WindowWR), .B0 (WindowDout_3__1__7), .B1 (nx8204)) ;
    dff L0_3_L1_0_Wij_reg_Dout_0 (.Q (WindowDout_3__0__0), .QB (\$dummy [64]), .D (
        nx3451), .CLK (CLK)) ;
    ao32 ix3452 (.Y (nx3451), .A0 (nx8088), .A1 (WindowDout_4__0__0), .A2 (
         WindowWR), .B0 (WindowDout_3__0__0), .B1 (nx8204)) ;
    dff L0_3_L1_0_Wij_reg_Dout_1 (.Q (WindowDout_3__0__1), .QB (\$dummy [65]), .D (
        nx3461), .CLK (CLK)) ;
    ao32 ix3462 (.Y (nx3461), .A0 (nx8088), .A1 (WindowDout_4__0__1), .A2 (
         WindowWR), .B0 (WindowDout_3__0__1), .B1 (nx8204)) ;
    dff L0_3_L1_0_Wij_reg_Dout_2 (.Q (WindowDout_3__0__2), .QB (\$dummy [66]), .D (
        nx3471), .CLK (CLK)) ;
    ao32 ix3472 (.Y (nx3471), .A0 (nx8088), .A1 (WindowDout_4__0__2), .A2 (
         WindowWR), .B0 (WindowDout_3__0__2), .B1 (nx8206)) ;
    dff L0_3_L1_0_Wij_reg_Dout_3 (.Q (WindowDout_3__0__3), .QB (\$dummy [67]), .D (
        nx3481), .CLK (CLK)) ;
    ao32 ix3482 (.Y (nx3481), .A0 (nx8088), .A1 (WindowDout_4__0__3), .A2 (
         WindowWR), .B0 (WindowDout_3__0__3), .B1 (nx8206)) ;
    dff L0_3_L1_0_Wij_reg_Dout_4 (.Q (WindowDout_3__0__4), .QB (\$dummy [68]), .D (
        nx3491), .CLK (CLK)) ;
    ao32 ix3492 (.Y (nx3491), .A0 (nx8088), .A1 (WindowDout_4__0__4), .A2 (
         WindowWR), .B0 (WindowDout_3__0__4), .B1 (nx8206)) ;
    dff L0_3_L1_0_Wij_reg_Dout_5 (.Q (WindowDout_3__0__5), .QB (\$dummy [69]), .D (
        nx3501), .CLK (CLK)) ;
    ao32 ix3502 (.Y (nx3501), .A0 (nx8088), .A1 (WindowDout_4__0__5), .A2 (
         WindowWR), .B0 (WindowDout_3__0__5), .B1 (nx8206)) ;
    dff L0_3_L1_0_Wij_reg_Dout_6 (.Q (WindowDout_3__0__6), .QB (\$dummy [70]), .D (
        nx3511), .CLK (CLK)) ;
    ao32 ix3512 (.Y (nx3511), .A0 (nx8090), .A1 (WindowDout_4__0__6), .A2 (
         WindowWR), .B0 (WindowDout_3__0__6), .B1 (nx8206)) ;
    dff L0_3_L1_0_Wij_reg_Dout_7 (.Q (WindowDout_3__0__7), .QB (\$dummy [71]), .D (
        nx3521), .CLK (CLK)) ;
    ao32 ix3522 (.Y (nx3521), .A0 (nx8090), .A1 (WindowDout_4__0__7), .A2 (
         WindowWR), .B0 (WindowDout_3__0__7), .B1 (nx8206)) ;
    oai21 ix3612 (.Y (nx3611), .A0 (nx6350), .A1 (nx7950), .B0 (nx6352)) ;
    dff L0_2_L1_4_Wij_reg_Dout_0 (.Q (WindowDout_2__4__0), .QB (nx6350), .D (
        nx3611), .CLK (CLK)) ;
    oai21 ix3622 (.Y (nx3621), .A0 (nx6356), .A1 (nx7950), .B0 (nx6358)) ;
    dff L0_2_L1_4_Wij_reg_Dout_1 (.Q (WindowDout_2__4__1), .QB (nx6356), .D (
        nx3621), .CLK (CLK)) ;
    oai21 ix3632 (.Y (nx3631), .A0 (nx6362), .A1 (nx7952), .B0 (nx6364)) ;
    dff L0_2_L1_4_Wij_reg_Dout_2 (.Q (WindowDout_2__4__2), .QB (nx6362), .D (
        nx3631), .CLK (CLK)) ;
    oai21 ix3642 (.Y (nx3641), .A0 (nx6368), .A1 (nx7952), .B0 (nx6370)) ;
    dff L0_2_L1_4_Wij_reg_Dout_3 (.Q (WindowDout_2__4__3), .QB (nx6368), .D (
        nx3641), .CLK (CLK)) ;
    oai21 ix3652 (.Y (nx3651), .A0 (nx6374), .A1 (nx7952), .B0 (nx6376)) ;
    dff L0_2_L1_4_Wij_reg_Dout_4 (.Q (WindowDout_2__4__4), .QB (nx6374), .D (
        nx3651), .CLK (CLK)) ;
    oai21 ix3662 (.Y (nx3661), .A0 (nx6380), .A1 (nx7954), .B0 (nx6382)) ;
    dff L0_2_L1_4_Wij_reg_Dout_5 (.Q (WindowDout_2__4__5), .QB (nx6380), .D (
        nx3661), .CLK (CLK)) ;
    oai21 ix3672 (.Y (nx3671), .A0 (nx6386), .A1 (nx7954), .B0 (nx6388)) ;
    dff L0_2_L1_4_Wij_reg_Dout_6 (.Q (WindowDout_2__4__6), .QB (nx6386), .D (
        nx3671), .CLK (CLK)) ;
    oai21 ix3682 (.Y (nx3681), .A0 (nx6392), .A1 (nx7954), .B0 (nx6394)) ;
    dff L0_2_L1_4_Wij_reg_Dout_7 (.Q (WindowDout_2__4__7), .QB (nx6392), .D (
        nx3681), .CLK (CLK)) ;
    oai21 ix3772 (.Y (nx3771), .A0 (nx6398), .A1 (nx7954), .B0 (nx6400)) ;
    dff L0_2_L1_3_Wij_reg_Dout_0 (.Q (WindowDout_2__3__0), .QB (nx6398), .D (
        nx3771), .CLK (CLK)) ;
    oai21 ix3782 (.Y (nx3781), .A0 (nx6404), .A1 (nx7956), .B0 (nx6406)) ;
    dff L0_2_L1_3_Wij_reg_Dout_1 (.Q (WindowDout_2__3__1), .QB (nx6404), .D (
        nx3781), .CLK (CLK)) ;
    oai21 ix3792 (.Y (nx3791), .A0 (nx6410), .A1 (nx7956), .B0 (nx6412)) ;
    dff L0_2_L1_3_Wij_reg_Dout_2 (.Q (WindowDout_2__3__2), .QB (nx6410), .D (
        nx3791), .CLK (CLK)) ;
    oai21 ix3802 (.Y (nx3801), .A0 (nx6416), .A1 (nx7956), .B0 (nx6418)) ;
    dff L0_2_L1_3_Wij_reg_Dout_3 (.Q (WindowDout_2__3__3), .QB (nx6416), .D (
        nx3801), .CLK (CLK)) ;
    oai21 ix3812 (.Y (nx3811), .A0 (nx6422), .A1 (nx7958), .B0 (nx6424)) ;
    dff L0_2_L1_3_Wij_reg_Dout_4 (.Q (WindowDout_2__3__4), .QB (nx6422), .D (
        nx3811), .CLK (CLK)) ;
    oai21 ix3822 (.Y (nx3821), .A0 (nx6428), .A1 (nx7958), .B0 (nx6430)) ;
    dff L0_2_L1_3_Wij_reg_Dout_5 (.Q (WindowDout_2__3__5), .QB (nx6428), .D (
        nx3821), .CLK (CLK)) ;
    oai21 ix3832 (.Y (nx3831), .A0 (nx6434), .A1 (nx7958), .B0 (nx6436)) ;
    dff L0_2_L1_3_Wij_reg_Dout_6 (.Q (WindowDout_2__3__6), .QB (nx6434), .D (
        nx3831), .CLK (CLK)) ;
    oai21 ix3842 (.Y (nx3841), .A0 (nx6440), .A1 (nx7958), .B0 (nx6442)) ;
    dff L0_2_L1_3_Wij_reg_Dout_7 (.Q (WindowDout_2__3__7), .QB (nx6440), .D (
        nx3841), .CLK (CLK)) ;
    dff L0_2_L1_2_Wij_reg_Dout_0 (.Q (WindowDout_2__2__0), .QB (\$dummy [72]), .D (
        nx3931), .CLK (CLK)) ;
    ao32 ix3932 (.Y (nx3931), .A0 (nx8094), .A1 (WindowDout_3__2__0), .A2 (
         WindowWR), .B0 (WindowDout_2__2__0), .B1 (nx8206)) ;
    dff L0_2_L1_2_Wij_reg_Dout_1 (.Q (WindowDout_2__2__1), .QB (\$dummy [73]), .D (
        nx3941), .CLK (CLK)) ;
    ao32 ix3942 (.Y (nx3941), .A0 (nx8094), .A1 (WindowDout_3__2__1), .A2 (
         WindowWR), .B0 (WindowDout_2__2__1), .B1 (nx8208)) ;
    dff L0_2_L1_2_Wij_reg_Dout_2 (.Q (WindowDout_2__2__2), .QB (\$dummy [74]), .D (
        nx3951), .CLK (CLK)) ;
    ao32 ix3952 (.Y (nx3951), .A0 (nx8094), .A1 (WindowDout_3__2__2), .A2 (
         WindowWR), .B0 (WindowDout_2__2__2), .B1 (nx8208)) ;
    dff L0_2_L1_2_Wij_reg_Dout_3 (.Q (WindowDout_2__2__3), .QB (\$dummy [75]), .D (
        nx3961), .CLK (CLK)) ;
    ao32 ix3962 (.Y (nx3961), .A0 (nx8096), .A1 (WindowDout_3__2__3), .A2 (
         WindowWR), .B0 (WindowDout_2__2__3), .B1 (nx8208)) ;
    dff L0_2_L1_2_Wij_reg_Dout_4 (.Q (WindowDout_2__2__4), .QB (\$dummy [76]), .D (
        nx3971), .CLK (CLK)) ;
    ao32 ix3972 (.Y (nx3971), .A0 (nx8096), .A1 (WindowDout_3__2__4), .A2 (
         WindowWR), .B0 (WindowDout_2__2__4), .B1 (nx8208)) ;
    dff L0_2_L1_2_Wij_reg_Dout_5 (.Q (WindowDout_2__2__5), .QB (\$dummy [77]), .D (
        nx3981), .CLK (CLK)) ;
    ao32 ix3982 (.Y (nx3981), .A0 (nx8096), .A1 (WindowDout_3__2__5), .A2 (
         WindowWR), .B0 (WindowDout_2__2__5), .B1 (nx8208)) ;
    dff L0_2_L1_2_Wij_reg_Dout_6 (.Q (WindowDout_2__2__6), .QB (\$dummy [78]), .D (
        nx3991), .CLK (CLK)) ;
    ao32 ix3992 (.Y (nx3991), .A0 (nx8096), .A1 (WindowDout_3__2__6), .A2 (
         WindowWR), .B0 (WindowDout_2__2__6), .B1 (nx8208)) ;
    dff L0_2_L1_2_Wij_reg_Dout_7 (.Q (WindowDout_2__2__7), .QB (\$dummy [79]), .D (
        nx4001), .CLK (CLK)) ;
    ao32 ix4002 (.Y (nx4001), .A0 (nx8096), .A1 (WindowDout_3__2__7), .A2 (
         WindowWR), .B0 (WindowDout_2__2__7), .B1 (nx8208)) ;
    dff L0_2_L1_1_Wij_reg_Dout_0 (.Q (WindowDout_2__1__0), .QB (\$dummy [80]), .D (
        nx4091), .CLK (CLK)) ;
    ao32 ix4092 (.Y (nx4091), .A0 (nx8096), .A1 (WindowDout_3__1__0), .A2 (
         WindowWR), .B0 (WindowDout_2__1__0), .B1 (nx8210)) ;
    dff L0_2_L1_1_Wij_reg_Dout_1 (.Q (WindowDout_2__1__1), .QB (\$dummy [81]), .D (
        nx4101), .CLK (CLK)) ;
    ao32 ix4102 (.Y (nx4101), .A0 (nx8096), .A1 (WindowDout_3__1__1), .A2 (
         WindowWR), .B0 (WindowDout_2__1__1), .B1 (nx8210)) ;
    dff L0_2_L1_1_Wij_reg_Dout_2 (.Q (WindowDout_2__1__2), .QB (\$dummy [82]), .D (
        nx4111), .CLK (CLK)) ;
    ao32 ix4112 (.Y (nx4111), .A0 (nx8098), .A1 (WindowDout_3__1__2), .A2 (
         WindowWR), .B0 (WindowDout_2__1__2), .B1 (nx8210)) ;
    dff L0_2_L1_1_Wij_reg_Dout_3 (.Q (WindowDout_2__1__3), .QB (\$dummy [83]), .D (
        nx4121), .CLK (CLK)) ;
    ao32 ix4122 (.Y (nx4121), .A0 (nx8098), .A1 (WindowDout_3__1__3), .A2 (
         WindowWR), .B0 (WindowDout_2__1__3), .B1 (nx8210)) ;
    dff L0_2_L1_1_Wij_reg_Dout_4 (.Q (WindowDout_2__1__4), .QB (\$dummy [84]), .D (
        nx4131), .CLK (CLK)) ;
    ao32 ix4132 (.Y (nx4131), .A0 (nx8098), .A1 (WindowDout_3__1__4), .A2 (
         WindowWR), .B0 (WindowDout_2__1__4), .B1 (nx8210)) ;
    dff L0_2_L1_1_Wij_reg_Dout_5 (.Q (WindowDout_2__1__5), .QB (\$dummy [85]), .D (
        nx4141), .CLK (CLK)) ;
    ao32 ix4142 (.Y (nx4141), .A0 (nx8098), .A1 (WindowDout_3__1__5), .A2 (
         WindowWR), .B0 (WindowDout_2__1__5), .B1 (nx8210)) ;
    dff L0_2_L1_1_Wij_reg_Dout_6 (.Q (WindowDout_2__1__6), .QB (\$dummy [86]), .D (
        nx4151), .CLK (CLK)) ;
    ao32 ix4152 (.Y (nx4151), .A0 (nx8098), .A1 (WindowDout_3__1__6), .A2 (
         WindowWR), .B0 (WindowDout_2__1__6), .B1 (nx8210)) ;
    dff L0_2_L1_1_Wij_reg_Dout_7 (.Q (WindowDout_2__1__7), .QB (\$dummy [87]), .D (
        nx4161), .CLK (CLK)) ;
    ao32 ix4162 (.Y (nx4161), .A0 (nx8098), .A1 (WindowDout_3__1__7), .A2 (
         WindowWR), .B0 (WindowDout_2__1__7), .B1 (nx8212)) ;
    dff L0_2_L1_0_Wij_reg_Dout_0 (.Q (WindowDout_2__0__0), .QB (\$dummy [88]), .D (
        nx4251), .CLK (CLK)) ;
    ao32 ix4252 (.Y (nx4251), .A0 (nx8098), .A1 (WindowDout_3__0__0), .A2 (
         WindowWR), .B0 (WindowDout_2__0__0), .B1 (nx8212)) ;
    dff L0_2_L1_0_Wij_reg_Dout_1 (.Q (WindowDout_2__0__1), .QB (\$dummy [89]), .D (
        nx4261), .CLK (CLK)) ;
    ao32 ix4262 (.Y (nx4261), .A0 (nx8100), .A1 (WindowDout_3__0__1), .A2 (
         WindowWR), .B0 (WindowDout_2__0__1), .B1 (nx8212)) ;
    dff L0_2_L1_0_Wij_reg_Dout_2 (.Q (WindowDout_2__0__2), .QB (\$dummy [90]), .D (
        nx4271), .CLK (CLK)) ;
    ao32 ix4272 (.Y (nx4271), .A0 (nx8100), .A1 (WindowDout_3__0__2), .A2 (
         WindowWR), .B0 (WindowDout_2__0__2), .B1 (nx8212)) ;
    dff L0_2_L1_0_Wij_reg_Dout_3 (.Q (WindowDout_2__0__3), .QB (\$dummy [91]), .D (
        nx4281), .CLK (CLK)) ;
    ao32 ix4282 (.Y (nx4281), .A0 (nx8100), .A1 (WindowDout_3__0__3), .A2 (
         WindowWR), .B0 (WindowDout_2__0__3), .B1 (nx8212)) ;
    dff L0_2_L1_0_Wij_reg_Dout_4 (.Q (WindowDout_2__0__4), .QB (\$dummy [92]), .D (
        nx4291), .CLK (CLK)) ;
    ao32 ix4292 (.Y (nx4291), .A0 (nx8100), .A1 (WindowDout_3__0__4), .A2 (
         WindowWR), .B0 (WindowDout_2__0__4), .B1 (nx8212)) ;
    dff L0_2_L1_0_Wij_reg_Dout_5 (.Q (WindowDout_2__0__5), .QB (\$dummy [93]), .D (
        nx4301), .CLK (CLK)) ;
    ao32 ix4302 (.Y (nx4301), .A0 (nx8100), .A1 (WindowDout_3__0__5), .A2 (
         WindowWR), .B0 (WindowDout_2__0__5), .B1 (nx8212)) ;
    dff L0_2_L1_0_Wij_reg_Dout_6 (.Q (WindowDout_2__0__6), .QB (\$dummy [94]), .D (
        nx4311), .CLK (CLK)) ;
    ao32 ix4312 (.Y (nx4311), .A0 (nx8100), .A1 (WindowDout_3__0__6), .A2 (
         WindowWR), .B0 (WindowDout_2__0__6), .B1 (nx8214)) ;
    dff L0_2_L1_0_Wij_reg_Dout_7 (.Q (WindowDout_2__0__7), .QB (\$dummy [95]), .D (
        nx4321), .CLK (CLK)) ;
    ao32 ix4322 (.Y (nx4321), .A0 (nx8100), .A1 (WindowDout_3__0__7), .A2 (
         WindowWR), .B0 (WindowDout_2__0__7), .B1 (nx8214)) ;
    oai21 ix4412 (.Y (nx4411), .A0 (nx6518), .A1 (nx7960), .B0 (nx6520)) ;
    dff L0_1_L1_4_Wij_reg_Dout_0 (.Q (WindowDout_1__4__0), .QB (nx6518), .D (
        nx4411), .CLK (CLK)) ;
    oai21 ix4422 (.Y (nx4421), .A0 (nx6524), .A1 (nx7960), .B0 (nx6526)) ;
    dff L0_1_L1_4_Wij_reg_Dout_1 (.Q (WindowDout_1__4__1), .QB (nx6524), .D (
        nx4421), .CLK (CLK)) ;
    oai21 ix4432 (.Y (nx4431), .A0 (nx6530), .A1 (nx7960), .B0 (nx6532)) ;
    dff L0_1_L1_4_Wij_reg_Dout_2 (.Q (WindowDout_1__4__2), .QB (nx6530), .D (
        nx4431), .CLK (CLK)) ;
    oai21 ix4442 (.Y (nx4441), .A0 (nx6536), .A1 (nx7962), .B0 (nx6538)) ;
    dff L0_1_L1_4_Wij_reg_Dout_3 (.Q (WindowDout_1__4__3), .QB (nx6536), .D (
        nx4441), .CLK (CLK)) ;
    oai21 ix4452 (.Y (nx4451), .A0 (nx6542), .A1 (nx7962), .B0 (nx6544)) ;
    dff L0_1_L1_4_Wij_reg_Dout_4 (.Q (WindowDout_1__4__4), .QB (nx6542), .D (
        nx4451), .CLK (CLK)) ;
    oai21 ix4462 (.Y (nx4461), .A0 (nx6548), .A1 (nx7962), .B0 (nx6550)) ;
    dff L0_1_L1_4_Wij_reg_Dout_5 (.Q (WindowDout_1__4__5), .QB (nx6548), .D (
        nx4461), .CLK (CLK)) ;
    oai21 ix4472 (.Y (nx4471), .A0 (nx6554), .A1 (nx7962), .B0 (nx6556)) ;
    dff L0_1_L1_4_Wij_reg_Dout_6 (.Q (WindowDout_1__4__6), .QB (nx6554), .D (
        nx4471), .CLK (CLK)) ;
    oai21 ix4482 (.Y (nx4481), .A0 (nx6560), .A1 (nx7964), .B0 (nx6562)) ;
    dff L0_1_L1_4_Wij_reg_Dout_7 (.Q (WindowDout_1__4__7), .QB (nx6560), .D (
        nx4481), .CLK (CLK)) ;
    oai21 ix4732 (.Y (nx4731), .A0 (nx6566), .A1 (nx7964), .B0 (nx6568)) ;
    dff L0_1_L1_3_Wij_reg_Dout_0 (.Q (WindowDout_1__3__0), .QB (nx6566), .D (
        nx4731), .CLK (CLK)) ;
    oai21 ix4742 (.Y (nx4741), .A0 (nx6572), .A1 (nx7964), .B0 (nx6574)) ;
    dff L0_1_L1_3_Wij_reg_Dout_1 (.Q (WindowDout_1__3__1), .QB (nx6572), .D (
        nx4741), .CLK (CLK)) ;
    oai21 ix4752 (.Y (nx4751), .A0 (nx6578), .A1 (nx7966), .B0 (nx6580)) ;
    dff L0_1_L1_3_Wij_reg_Dout_2 (.Q (WindowDout_1__3__2), .QB (nx6578), .D (
        nx4751), .CLK (CLK)) ;
    oai21 ix4762 (.Y (nx4761), .A0 (nx6584), .A1 (nx7966), .B0 (nx6586)) ;
    dff L0_1_L1_3_Wij_reg_Dout_3 (.Q (WindowDout_1__3__3), .QB (nx6584), .D (
        nx4761), .CLK (CLK)) ;
    oai21 ix4772 (.Y (nx4771), .A0 (nx6590), .A1 (nx7966), .B0 (nx6592)) ;
    dff L0_1_L1_3_Wij_reg_Dout_4 (.Q (WindowDout_1__3__4), .QB (nx6590), .D (
        nx4771), .CLK (CLK)) ;
    oai21 ix4782 (.Y (nx4781), .A0 (nx6596), .A1 (nx7966), .B0 (nx6598)) ;
    dff L0_1_L1_3_Wij_reg_Dout_5 (.Q (WindowDout_1__3__5), .QB (nx6596), .D (
        nx4781), .CLK (CLK)) ;
    oai21 ix4792 (.Y (nx4791), .A0 (nx6602), .A1 (nx7968), .B0 (nx6604)) ;
    dff L0_1_L1_3_Wij_reg_Dout_6 (.Q (WindowDout_1__3__6), .QB (nx6602), .D (
        nx4791), .CLK (CLK)) ;
    oai21 ix4802 (.Y (nx4801), .A0 (nx6608), .A1 (nx7968), .B0 (nx6610)) ;
    dff L0_1_L1_3_Wij_reg_Dout_7 (.Q (WindowDout_1__3__7), .QB (nx6608), .D (
        nx4801), .CLK (CLK)) ;
    oai21 ix5052 (.Y (nx5051), .A0 (nx6614), .A1 (nx7968), .B0 (nx6616)) ;
    dff L0_1_L1_2_Wij_reg_Dout_0 (.Q (WindowDout_1__2__0), .QB (nx6614), .D (
        nx5051), .CLK (CLK)) ;
    nand03 ix6617 (.Y (nx6616), .A0 (nx8106), .A1 (WindowDout_2__2__0), .A2 (
           nx7968)) ;
    oai21 ix5062 (.Y (nx5061), .A0 (nx6620), .A1 (nx7970), .B0 (nx6622)) ;
    dff L0_1_L1_2_Wij_reg_Dout_1 (.Q (WindowDout_1__2__1), .QB (nx6620), .D (
        nx5061), .CLK (CLK)) ;
    nand03 ix6623 (.Y (nx6622), .A0 (nx8106), .A1 (WindowDout_2__2__1), .A2 (
           nx7970)) ;
    oai21 ix5072 (.Y (nx5071), .A0 (nx6626), .A1 (nx7970), .B0 (nx6628)) ;
    dff L0_1_L1_2_Wij_reg_Dout_2 (.Q (WindowDout_1__2__2), .QB (nx6626), .D (
        nx5071), .CLK (CLK)) ;
    nand03 ix6629 (.Y (nx6628), .A0 (nx8106), .A1 (WindowDout_2__2__2), .A2 (
           nx7970)) ;
    oai21 ix5082 (.Y (nx5081), .A0 (nx6632), .A1 (nx7970), .B0 (nx6634)) ;
    dff L0_1_L1_2_Wij_reg_Dout_3 (.Q (WindowDout_1__2__3), .QB (nx6632), .D (
        nx5081), .CLK (CLK)) ;
    nand03 ix6635 (.Y (nx6634), .A0 (nx8106), .A1 (WindowDout_2__2__3), .A2 (
           nx7970)) ;
    oai21 ix5092 (.Y (nx5091), .A0 (nx6638), .A1 (nx7970), .B0 (nx6640)) ;
    dff L0_1_L1_2_Wij_reg_Dout_4 (.Q (WindowDout_1__2__4), .QB (nx6638), .D (
        nx5091), .CLK (CLK)) ;
    nand03 ix6641 (.Y (nx6640), .A0 (nx8106), .A1 (WindowDout_2__2__4), .A2 (
           nx7972)) ;
    oai21 ix5102 (.Y (nx5101), .A0 (nx6644), .A1 (nx7972), .B0 (nx6646)) ;
    dff L0_1_L1_2_Wij_reg_Dout_5 (.Q (WindowDout_1__2__5), .QB (nx6644), .D (
        nx5101), .CLK (CLK)) ;
    nand03 ix6647 (.Y (nx6646), .A0 (nx8108), .A1 (WindowDout_2__2__5), .A2 (
           nx7972)) ;
    oai21 ix5112 (.Y (nx5111), .A0 (nx6650), .A1 (nx7972), .B0 (nx6652)) ;
    dff L0_1_L1_2_Wij_reg_Dout_6 (.Q (WindowDout_1__2__6), .QB (nx6650), .D (
        nx5111), .CLK (CLK)) ;
    nand03 ix6653 (.Y (nx6652), .A0 (nx8108), .A1 (WindowDout_2__2__6), .A2 (
           nx7972)) ;
    oai21 ix5122 (.Y (nx5121), .A0 (nx6656), .A1 (nx7972), .B0 (nx6658)) ;
    dff L0_1_L1_2_Wij_reg_Dout_7 (.Q (WindowDout_1__2__7), .QB (nx6656), .D (
        nx5121), .CLK (CLK)) ;
    nand03 ix6659 (.Y (nx6658), .A0 (nx8108), .A1 (WindowDout_2__2__7), .A2 (
           nx7972)) ;
    oai21 ix5372 (.Y (nx5371), .A0 (nx6662), .A1 (nx7974), .B0 (nx6664)) ;
    dff L0_1_L1_1_Wij_reg_Dout_0 (.Q (WindowDout_1__1__0), .QB (nx6662), .D (
        nx5371), .CLK (CLK)) ;
    nand03 ix6665 (.Y (nx6664), .A0 (nx8108), .A1 (WindowDout_2__1__0), .A2 (
           nx7974)) ;
    oai21 ix5382 (.Y (nx5381), .A0 (nx6668), .A1 (nx7974), .B0 (nx6670)) ;
    dff L0_1_L1_1_Wij_reg_Dout_1 (.Q (WindowDout_1__1__1), .QB (nx6668), .D (
        nx5381), .CLK (CLK)) ;
    nand03 ix6671 (.Y (nx6670), .A0 (nx8108), .A1 (WindowDout_2__1__1), .A2 (
           nx7974)) ;
    oai21 ix5392 (.Y (nx5391), .A0 (nx6674), .A1 (nx7974), .B0 (nx6676)) ;
    dff L0_1_L1_1_Wij_reg_Dout_2 (.Q (WindowDout_1__1__2), .QB (nx6674), .D (
        nx5391), .CLK (CLK)) ;
    nand03 ix6677 (.Y (nx6676), .A0 (nx8108), .A1 (WindowDout_2__1__2), .A2 (
           nx7974)) ;
    oai21 ix5402 (.Y (nx5401), .A0 (nx6680), .A1 (nx7974), .B0 (nx6682)) ;
    dff L0_1_L1_1_Wij_reg_Dout_3 (.Q (WindowDout_1__1__3), .QB (nx6680), .D (
        nx5401), .CLK (CLK)) ;
    nand03 ix6683 (.Y (nx6682), .A0 (nx8108), .A1 (WindowDout_2__1__3), .A2 (
           nx7976)) ;
    oai21 ix5412 (.Y (nx5411), .A0 (nx6686), .A1 (nx7976), .B0 (nx6688)) ;
    dff L0_1_L1_1_Wij_reg_Dout_4 (.Q (WindowDout_1__1__4), .QB (nx6686), .D (
        nx5411), .CLK (CLK)) ;
    nand03 ix6689 (.Y (nx6688), .A0 (nx8110), .A1 (WindowDout_2__1__4), .A2 (
           nx7976)) ;
    oai21 ix5422 (.Y (nx5421), .A0 (nx6692), .A1 (nx7976), .B0 (nx6694)) ;
    dff L0_1_L1_1_Wij_reg_Dout_5 (.Q (WindowDout_1__1__5), .QB (nx6692), .D (
        nx5421), .CLK (CLK)) ;
    nand03 ix6695 (.Y (nx6694), .A0 (nx8110), .A1 (WindowDout_2__1__5), .A2 (
           nx7976)) ;
    oai21 ix5432 (.Y (nx5431), .A0 (nx6698), .A1 (nx7976), .B0 (nx6700)) ;
    dff L0_1_L1_1_Wij_reg_Dout_6 (.Q (WindowDout_1__1__6), .QB (nx6698), .D (
        nx5431), .CLK (CLK)) ;
    nand03 ix6701 (.Y (nx6700), .A0 (nx8110), .A1 (WindowDout_2__1__6), .A2 (
           nx7976)) ;
    oai21 ix5442 (.Y (nx5441), .A0 (nx6704), .A1 (nx7978), .B0 (nx6706)) ;
    dff L0_1_L1_1_Wij_reg_Dout_7 (.Q (WindowDout_1__1__7), .QB (nx6704), .D (
        nx5441), .CLK (CLK)) ;
    nand03 ix6707 (.Y (nx6706), .A0 (nx8110), .A1 (WindowDout_2__1__7), .A2 (
           nx7978)) ;
    oai21 ix5692 (.Y (nx5691), .A0 (nx6710), .A1 (nx7978), .B0 (nx6712)) ;
    dff L0_1_L1_0_Wij_reg_Dout_0 (.Q (WindowDout_1__0__0), .QB (nx6710), .D (
        nx5691), .CLK (CLK)) ;
    nand03 ix6713 (.Y (nx6712), .A0 (nx8110), .A1 (WindowDout_2__0__0), .A2 (
           nx7978)) ;
    oai21 ix5702 (.Y (nx5701), .A0 (nx6716), .A1 (nx7978), .B0 (nx6718)) ;
    dff L0_1_L1_0_Wij_reg_Dout_1 (.Q (WindowDout_1__0__1), .QB (nx6716), .D (
        nx5701), .CLK (CLK)) ;
    nand03 ix6719 (.Y (nx6718), .A0 (nx8110), .A1 (WindowDout_2__0__1), .A2 (
           nx7978)) ;
    oai21 ix5712 (.Y (nx5711), .A0 (nx6722), .A1 (nx7978), .B0 (nx6724)) ;
    dff L0_1_L1_0_Wij_reg_Dout_2 (.Q (WindowDout_1__0__2), .QB (nx6722), .D (
        nx5711), .CLK (CLK)) ;
    nand03 ix6725 (.Y (nx6724), .A0 (nx8110), .A1 (WindowDout_2__0__2), .A2 (
           nx7980)) ;
    oai21 ix5722 (.Y (nx5721), .A0 (nx6728), .A1 (nx7980), .B0 (nx6730)) ;
    dff L0_1_L1_0_Wij_reg_Dout_3 (.Q (WindowDout_1__0__3), .QB (nx6728), .D (
        nx5721), .CLK (CLK)) ;
    nand03 ix6731 (.Y (nx6730), .A0 (nx8112), .A1 (WindowDout_2__0__3), .A2 (
           nx7980)) ;
    oai21 ix5732 (.Y (nx5731), .A0 (nx6734), .A1 (nx7980), .B0 (nx6736)) ;
    dff L0_1_L1_0_Wij_reg_Dout_4 (.Q (WindowDout_1__0__4), .QB (nx6734), .D (
        nx5731), .CLK (CLK)) ;
    nand03 ix6737 (.Y (nx6736), .A0 (nx8112), .A1 (WindowDout_2__0__4), .A2 (
           nx7980)) ;
    oai21 ix5742 (.Y (nx5741), .A0 (nx6740), .A1 (nx7980), .B0 (nx6742)) ;
    dff L0_1_L1_0_Wij_reg_Dout_5 (.Q (WindowDout_1__0__5), .QB (nx6740), .D (
        nx5741), .CLK (CLK)) ;
    nand03 ix6743 (.Y (nx6742), .A0 (nx8112), .A1 (WindowDout_2__0__5), .A2 (
           nx7980)) ;
    oai21 ix5752 (.Y (nx5751), .A0 (nx6746), .A1 (nx7982), .B0 (nx6748)) ;
    dff L0_1_L1_0_Wij_reg_Dout_6 (.Q (WindowDout_1__0__6), .QB (nx6746), .D (
        nx5751), .CLK (CLK)) ;
    nand03 ix6749 (.Y (nx6748), .A0 (nx8112), .A1 (WindowDout_2__0__6), .A2 (
           nx7982)) ;
    oai21 ix5762 (.Y (nx5761), .A0 (nx6752), .A1 (nx7982), .B0 (nx6754)) ;
    dff L0_1_L1_0_Wij_reg_Dout_7 (.Q (WindowDout_1__0__7), .QB (nx6752), .D (
        nx5761), .CLK (CLK)) ;
    nand03 ix6755 (.Y (nx6754), .A0 (nx8112), .A1 (WindowDout_2__0__7), .A2 (
           nx7982)) ;
    oai21 ix4492 (.Y (nx4491), .A0 (nx6758), .A1 (nx7982), .B0 (nx6760)) ;
    dff L0_0_L1_4_Wij_reg_Dout_0 (.Q (WindowDout_0__4__0), .QB (nx6758), .D (
        nx4491), .CLK (CLK)) ;
    oai21 ix4502 (.Y (nx4501), .A0 (nx6764), .A1 (nx7982), .B0 (nx6766)) ;
    dff L0_0_L1_4_Wij_reg_Dout_1 (.Q (WindowDout_0__4__1), .QB (nx6764), .D (
        nx4501), .CLK (CLK)) ;
    oai21 ix4512 (.Y (nx4511), .A0 (nx6770), .A1 (nx7984), .B0 (nx6772)) ;
    dff L0_0_L1_4_Wij_reg_Dout_2 (.Q (WindowDout_0__4__2), .QB (nx6770), .D (
        nx4511), .CLK (CLK)) ;
    oai21 ix4522 (.Y (nx4521), .A0 (nx6776), .A1 (nx7984), .B0 (nx6778)) ;
    dff L0_0_L1_4_Wij_reg_Dout_3 (.Q (WindowDout_0__4__3), .QB (nx6776), .D (
        nx4521), .CLK (CLK)) ;
    oai21 ix4532 (.Y (nx4531), .A0 (nx6782), .A1 (nx7984), .B0 (nx6784)) ;
    dff L0_0_L1_4_Wij_reg_Dout_4 (.Q (WindowDout_0__4__4), .QB (nx6782), .D (
        nx4531), .CLK (CLK)) ;
    oai21 ix4542 (.Y (nx4541), .A0 (nx6788), .A1 (nx7986), .B0 (nx6790)) ;
    dff L0_0_L1_4_Wij_reg_Dout_5 (.Q (WindowDout_0__4__5), .QB (nx6788), .D (
        nx4541), .CLK (CLK)) ;
    oai21 ix4552 (.Y (nx4551), .A0 (nx6794), .A1 (nx7986), .B0 (nx6796)) ;
    dff L0_0_L1_4_Wij_reg_Dout_6 (.Q (WindowDout_0__4__6), .QB (nx6794), .D (
        nx4551), .CLK (CLK)) ;
    oai21 ix4562 (.Y (nx4561), .A0 (nx6800), .A1 (nx7986), .B0 (nx6802)) ;
    dff L0_0_L1_4_Wij_reg_Dout_7 (.Q (WindowDout_0__4__7), .QB (nx6800), .D (
        nx4561), .CLK (CLK)) ;
    oai21 ix4812 (.Y (nx4811), .A0 (nx6806), .A1 (nx7986), .B0 (nx6808)) ;
    dff L0_0_L1_3_Wij_reg_Dout_0 (.Q (WindowDout_0__3__0), .QB (nx6806), .D (
        nx4811), .CLK (CLK)) ;
    oai21 ix4822 (.Y (nx4821), .A0 (nx6812), .A1 (nx7988), .B0 (nx6814)) ;
    dff L0_0_L1_3_Wij_reg_Dout_1 (.Q (WindowDout_0__3__1), .QB (nx6812), .D (
        nx4821), .CLK (CLK)) ;
    oai21 ix4832 (.Y (nx4831), .A0 (nx6818), .A1 (nx7988), .B0 (nx6820)) ;
    dff L0_0_L1_3_Wij_reg_Dout_2 (.Q (WindowDout_0__3__2), .QB (nx6818), .D (
        nx4831), .CLK (CLK)) ;
    oai21 ix4842 (.Y (nx4841), .A0 (nx6824), .A1 (nx7988), .B0 (nx6826)) ;
    dff L0_0_L1_3_Wij_reg_Dout_3 (.Q (WindowDout_0__3__3), .QB (nx6824), .D (
        nx4841), .CLK (CLK)) ;
    oai21 ix4852 (.Y (nx4851), .A0 (nx6830), .A1 (nx7990), .B0 (nx6832)) ;
    dff L0_0_L1_3_Wij_reg_Dout_4 (.Q (WindowDout_0__3__4), .QB (nx6830), .D (
        nx4851), .CLK (CLK)) ;
    oai21 ix4862 (.Y (nx4861), .A0 (nx6836), .A1 (nx7990), .B0 (nx6838)) ;
    dff L0_0_L1_3_Wij_reg_Dout_5 (.Q (WindowDout_0__3__5), .QB (nx6836), .D (
        nx4861), .CLK (CLK)) ;
    oai21 ix4872 (.Y (nx4871), .A0 (nx6842), .A1 (nx7990), .B0 (nx6844)) ;
    dff L0_0_L1_3_Wij_reg_Dout_6 (.Q (WindowDout_0__3__6), .QB (nx6842), .D (
        nx4871), .CLK (CLK)) ;
    oai21 ix4882 (.Y (nx4881), .A0 (nx6848), .A1 (nx7990), .B0 (nx6850)) ;
    dff L0_0_L1_3_Wij_reg_Dout_7 (.Q (WindowDout_0__3__7), .QB (nx6848), .D (
        nx4881), .CLK (CLK)) ;
    oai21 ix5132 (.Y (nx5131), .A0 (nx6854), .A1 (nx7992), .B0 (nx6856)) ;
    dff L0_0_L1_2_Wij_reg_Dout_0 (.Q (WindowDout_0__2__0), .QB (nx6854), .D (
        nx5131), .CLK (CLK)) ;
    oai21 ix5142 (.Y (nx5141), .A0 (nx6860), .A1 (nx7992), .B0 (nx6862)) ;
    dff L0_0_L1_2_Wij_reg_Dout_1 (.Q (WindowDout_0__2__1), .QB (nx6860), .D (
        nx5141), .CLK (CLK)) ;
    oai21 ix5152 (.Y (nx5151), .A0 (nx6866), .A1 (nx7992), .B0 (nx6868)) ;
    dff L0_0_L1_2_Wij_reg_Dout_2 (.Q (WindowDout_0__2__2), .QB (nx6866), .D (
        nx5151), .CLK (CLK)) ;
    oai21 ix5162 (.Y (nx5161), .A0 (nx6872), .A1 (nx7994), .B0 (nx6874)) ;
    dff L0_0_L1_2_Wij_reg_Dout_3 (.Q (WindowDout_0__2__3), .QB (nx6872), .D (
        nx5161), .CLK (CLK)) ;
    oai21 ix5172 (.Y (nx5171), .A0 (nx6878), .A1 (nx7994), .B0 (nx6880)) ;
    dff L0_0_L1_2_Wij_reg_Dout_4 (.Q (WindowDout_0__2__4), .QB (nx6878), .D (
        nx5171), .CLK (CLK)) ;
    oai21 ix5182 (.Y (nx5181), .A0 (nx6884), .A1 (nx7994), .B0 (nx6886)) ;
    dff L0_0_L1_2_Wij_reg_Dout_5 (.Q (WindowDout_0__2__5), .QB (nx6884), .D (
        nx5181), .CLK (CLK)) ;
    oai21 ix5192 (.Y (nx5191), .A0 (nx6890), .A1 (nx7994), .B0 (nx6892)) ;
    dff L0_0_L1_2_Wij_reg_Dout_6 (.Q (WindowDout_0__2__6), .QB (nx6890), .D (
        nx5191), .CLK (CLK)) ;
    oai21 ix5202 (.Y (nx5201), .A0 (nx6896), .A1 (nx7996), .B0 (nx6898)) ;
    dff L0_0_L1_2_Wij_reg_Dout_7 (.Q (WindowDout_0__2__7), .QB (nx6896), .D (
        nx5201), .CLK (CLK)) ;
    oai21 ix5452 (.Y (nx5451), .A0 (nx6902), .A1 (nx7996), .B0 (nx6904)) ;
    dff L0_0_L1_1_Wij_reg_Dout_0 (.Q (WindowDout_0__1__0), .QB (nx6902), .D (
        nx5451), .CLK (CLK)) ;
    oai21 ix5462 (.Y (nx5461), .A0 (nx6908), .A1 (nx7996), .B0 (nx6910)) ;
    dff L0_0_L1_1_Wij_reg_Dout_1 (.Q (WindowDout_0__1__1), .QB (nx6908), .D (
        nx5461), .CLK (CLK)) ;
    oai21 ix5472 (.Y (nx5471), .A0 (nx6914), .A1 (nx7998), .B0 (nx6916)) ;
    dff L0_0_L1_1_Wij_reg_Dout_2 (.Q (WindowDout_0__1__2), .QB (nx6914), .D (
        nx5471), .CLK (CLK)) ;
    oai21 ix5482 (.Y (nx5481), .A0 (nx6920), .A1 (nx7998), .B0 (nx6922)) ;
    dff L0_0_L1_1_Wij_reg_Dout_3 (.Q (WindowDout_0__1__3), .QB (nx6920), .D (
        nx5481), .CLK (CLK)) ;
    oai21 ix5492 (.Y (nx5491), .A0 (nx6926), .A1 (nx7998), .B0 (nx6928)) ;
    dff L0_0_L1_1_Wij_reg_Dout_4 (.Q (WindowDout_0__1__4), .QB (nx6926), .D (
        nx5491), .CLK (CLK)) ;
    oai21 ix5502 (.Y (nx5501), .A0 (nx6932), .A1 (nx7998), .B0 (nx6934)) ;
    dff L0_0_L1_1_Wij_reg_Dout_5 (.Q (WindowDout_0__1__5), .QB (nx6932), .D (
        nx5501), .CLK (CLK)) ;
    oai21 ix5512 (.Y (nx5511), .A0 (nx6938), .A1 (nx8000), .B0 (nx6940)) ;
    dff L0_0_L1_1_Wij_reg_Dout_6 (.Q (WindowDout_0__1__6), .QB (nx6938), .D (
        nx5511), .CLK (CLK)) ;
    oai21 ix5522 (.Y (nx5521), .A0 (nx6944), .A1 (nx8000), .B0 (nx6946)) ;
    dff L0_0_L1_1_Wij_reg_Dout_7 (.Q (WindowDout_0__1__7), .QB (nx6944), .D (
        nx5521), .CLK (CLK)) ;
    oai21 ix5772 (.Y (nx5771), .A0 (nx6950), .A1 (nx8000), .B0 (nx6952)) ;
    dff L0_0_L1_0_Wij_reg_Dout_0 (.Q (WindowDout_0__0__0), .QB (nx6950), .D (
        nx5771), .CLK (CLK)) ;
    oai21 ix5782 (.Y (nx5781), .A0 (nx6956), .A1 (nx8002), .B0 (nx6958)) ;
    dff L0_0_L1_0_Wij_reg_Dout_1 (.Q (WindowDout_0__0__1), .QB (nx6956), .D (
        nx5781), .CLK (CLK)) ;
    oai21 ix5792 (.Y (nx5791), .A0 (nx6962), .A1 (nx8002), .B0 (nx6964)) ;
    dff L0_0_L1_0_Wij_reg_Dout_2 (.Q (WindowDout_0__0__2), .QB (nx6962), .D (
        nx5791), .CLK (CLK)) ;
    oai21 ix5802 (.Y (nx5801), .A0 (nx6968), .A1 (nx8002), .B0 (nx6970)) ;
    dff L0_0_L1_0_Wij_reg_Dout_3 (.Q (WindowDout_0__0__3), .QB (nx6968), .D (
        nx5801), .CLK (CLK)) ;
    oai21 ix5812 (.Y (nx5811), .A0 (nx6974), .A1 (nx8002), .B0 (nx6976)) ;
    dff L0_0_L1_0_Wij_reg_Dout_4 (.Q (WindowDout_0__0__4), .QB (nx6974), .D (
        nx5811), .CLK (CLK)) ;
    oai21 ix5822 (.Y (nx5821), .A0 (nx6980), .A1 (nx8004), .B0 (nx6982)) ;
    dff L0_0_L1_0_Wij_reg_Dout_5 (.Q (WindowDout_0__0__5), .QB (nx6980), .D (
        nx5821), .CLK (CLK)) ;
    oai21 ix5832 (.Y (nx5831), .A0 (nx6986), .A1 (nx8004), .B0 (nx6988)) ;
    dff L0_0_L1_0_Wij_reg_Dout_6 (.Q (WindowDout_0__0__6), .QB (nx6986), .D (
        nx5831), .CLK (CLK)) ;
    oai21 ix5842 (.Y (nx5841), .A0 (nx6992), .A1 (nx8004), .B0 (nx6994)) ;
    dff L0_0_L1_0_Wij_reg_Dout_7 (.Q (WindowDout_0__0__7), .QB (nx6992), .D (
        nx5841), .CLK (CLK)) ;
    dff L0_4_L1_4_Fij_reg_Dout_0 (.Q (FilterDout_4__4__0), .QB (\$dummy [96]), .D (
        nx2091), .CLK (CLK)) ;
    aoi21 ix6999 (.Y (nx6998), .A0 (FilterSize), .A1 (FilterWR), .B0 (RST)) ;
    dff L0_4_L1_4_Fij_reg_Dout_1 (.Q (FilterDout_4__4__1), .QB (\$dummy [97]), .D (
        nx2101), .CLK (CLK)) ;
    dff L0_4_L1_4_Fij_reg_Dout_2 (.Q (FilterDout_4__4__2), .QB (\$dummy [98]), .D (
        nx2111), .CLK (CLK)) ;
    dff L0_4_L1_4_Fij_reg_Dout_3 (.Q (FilterDout_4__4__3), .QB (\$dummy [99]), .D (
        nx2121), .CLK (CLK)) ;
    dff L0_4_L1_4_Fij_reg_Dout_4 (.Q (FilterDout_4__4__4), .QB (\$dummy [100]), 
        .D (nx2131), .CLK (CLK)) ;
    dff L0_4_L1_4_Fij_reg_Dout_5 (.Q (FilterDout_4__4__5), .QB (\$dummy [101]), 
        .D (nx2141), .CLK (CLK)) ;
    dff L0_4_L1_4_Fij_reg_Dout_6 (.Q (FilterDout_4__4__6), .QB (\$dummy [102]), 
        .D (nx2151), .CLK (CLK)) ;
    dff L0_4_L1_4_Fij_reg_Dout_7 (.Q (FilterDout_4__4__7), .QB (\$dummy [103]), 
        .D (nx2161), .CLK (CLK)) ;
    dff L0_4_L1_3_Fij_reg_Dout_0 (.Q (FilterDout_4__3__0), .QB (\$dummy [104]), 
        .D (nx2251), .CLK (CLK)) ;
    dff L0_4_L1_3_Fij_reg_Dout_1 (.Q (FilterDout_4__3__1), .QB (\$dummy [105]), 
        .D (nx2261), .CLK (CLK)) ;
    dff L0_4_L1_3_Fij_reg_Dout_2 (.Q (FilterDout_4__3__2), .QB (\$dummy [106]), 
        .D (nx2271), .CLK (CLK)) ;
    dff L0_4_L1_3_Fij_reg_Dout_3 (.Q (FilterDout_4__3__3), .QB (\$dummy [107]), 
        .D (nx2281), .CLK (CLK)) ;
    dff L0_4_L1_3_Fij_reg_Dout_4 (.Q (FilterDout_4__3__4), .QB (\$dummy [108]), 
        .D (nx2291), .CLK (CLK)) ;
    dff L0_4_L1_3_Fij_reg_Dout_5 (.Q (FilterDout_4__3__5), .QB (\$dummy [109]), 
        .D (nx2301), .CLK (CLK)) ;
    dff L0_4_L1_3_Fij_reg_Dout_6 (.Q (FilterDout_4__3__6), .QB (\$dummy [110]), 
        .D (nx2311), .CLK (CLK)) ;
    dff L0_4_L1_3_Fij_reg_Dout_7 (.Q (FilterDout_4__3__7), .QB (\$dummy [111]), 
        .D (nx2321), .CLK (CLK)) ;
    dff L0_4_L1_2_Fij_reg_Dout_0 (.Q (FilterDout_4__2__0), .QB (\$dummy [112]), 
        .D (nx2411), .CLK (CLK)) ;
    ao32 ix2412 (.Y (nx2411), .A0 (Din[16]), .A1 (nx8124), .A2 (FilterWR), .B0 (
         FilterDout_4__2__0), .B1 (nx8232)) ;
    nor02_2x ix7049 (.Y (nx7048), .A0 (FilterWR), .A1 (RST)) ;
    dff L0_4_L1_2_Fij_reg_Dout_1 (.Q (FilterDout_4__2__1), .QB (\$dummy [113]), 
        .D (nx2421), .CLK (CLK)) ;
    ao32 ix2422 (.Y (nx2421), .A0 (Din[17]), .A1 (nx8124), .A2 (FilterWR), .B0 (
         FilterDout_4__2__1), .B1 (nx8232)) ;
    dff L0_4_L1_2_Fij_reg_Dout_2 (.Q (FilterDout_4__2__2), .QB (\$dummy [114]), 
        .D (nx2431), .CLK (CLK)) ;
    ao32 ix2432 (.Y (nx2431), .A0 (Din[18]), .A1 (nx8124), .A2 (FilterWR), .B0 (
         FilterDout_4__2__2), .B1 (nx8232)) ;
    dff L0_4_L1_2_Fij_reg_Dout_3 (.Q (FilterDout_4__2__3), .QB (\$dummy [115]), 
        .D (nx2441), .CLK (CLK)) ;
    ao32 ix2442 (.Y (nx2441), .A0 (Din[19]), .A1 (nx8124), .A2 (FilterWR), .B0 (
         FilterDout_4__2__3), .B1 (nx8232)) ;
    dff L0_4_L1_2_Fij_reg_Dout_4 (.Q (FilterDout_4__2__4), .QB (\$dummy [116]), 
        .D (nx2451), .CLK (CLK)) ;
    ao32 ix2452 (.Y (nx2451), .A0 (Din[20]), .A1 (nx8126), .A2 (FilterWR), .B0 (
         FilterDout_4__2__4), .B1 (nx8232)) ;
    dff L0_4_L1_2_Fij_reg_Dout_5 (.Q (FilterDout_4__2__5), .QB (\$dummy [117]), 
        .D (nx2461), .CLK (CLK)) ;
    ao32 ix2462 (.Y (nx2461), .A0 (Din[21]), .A1 (nx8126), .A2 (FilterWR), .B0 (
         FilterDout_4__2__5), .B1 (nx8232)) ;
    dff L0_4_L1_2_Fij_reg_Dout_6 (.Q (FilterDout_4__2__6), .QB (\$dummy [118]), 
        .D (nx2471), .CLK (CLK)) ;
    ao32 ix2472 (.Y (nx2471), .A0 (Din[22]), .A1 (nx8126), .A2 (FilterWR), .B0 (
         FilterDout_4__2__6), .B1 (nx8232)) ;
    dff L0_4_L1_2_Fij_reg_Dout_7 (.Q (FilterDout_4__2__7), .QB (\$dummy [119]), 
        .D (nx2481), .CLK (CLK)) ;
    ao32 ix2482 (.Y (nx2481), .A0 (Din[23]), .A1 (nx8126), .A2 (FilterWR), .B0 (
         FilterDout_4__2__7), .B1 (nx8234)) ;
    dff L0_4_L1_1_Fij_reg_Dout_0 (.Q (FilterDout_4__1__0), .QB (\$dummy [120]), 
        .D (nx2571), .CLK (CLK)) ;
    ao32 ix2572 (.Y (nx2571), .A0 (Din[8]), .A1 (nx8126), .A2 (FilterWR), .B0 (
         FilterDout_4__1__0), .B1 (nx8234)) ;
    dff L0_4_L1_1_Fij_reg_Dout_1 (.Q (FilterDout_4__1__1), .QB (\$dummy [121]), 
        .D (nx2581), .CLK (CLK)) ;
    ao32 ix2582 (.Y (nx2581), .A0 (Din[9]), .A1 (nx8126), .A2 (FilterWR), .B0 (
         FilterDout_4__1__1), .B1 (nx8234)) ;
    dff L0_4_L1_1_Fij_reg_Dout_2 (.Q (FilterDout_4__1__2), .QB (\$dummy [122]), 
        .D (nx2591), .CLK (CLK)) ;
    ao32 ix2592 (.Y (nx2591), .A0 (Din[10]), .A1 (nx8126), .A2 (FilterWR), .B0 (
         FilterDout_4__1__2), .B1 (nx8234)) ;
    dff L0_4_L1_1_Fij_reg_Dout_3 (.Q (FilterDout_4__1__3), .QB (\$dummy [123]), 
        .D (nx2601), .CLK (CLK)) ;
    ao32 ix2602 (.Y (nx2601), .A0 (Din[11]), .A1 (nx8128), .A2 (FilterWR), .B0 (
         FilterDout_4__1__3), .B1 (nx8234)) ;
    dff L0_4_L1_1_Fij_reg_Dout_4 (.Q (FilterDout_4__1__4), .QB (\$dummy [124]), 
        .D (nx2611), .CLK (CLK)) ;
    ao32 ix2612 (.Y (nx2611), .A0 (Din[12]), .A1 (nx8128), .A2 (FilterWR), .B0 (
         FilterDout_4__1__4), .B1 (nx8234)) ;
    dff L0_4_L1_1_Fij_reg_Dout_5 (.Q (FilterDout_4__1__5), .QB (\$dummy [125]), 
        .D (nx2621), .CLK (CLK)) ;
    ao32 ix2622 (.Y (nx2621), .A0 (Din[13]), .A1 (nx8128), .A2 (FilterWR), .B0 (
         FilterDout_4__1__5), .B1 (nx8234)) ;
    dff L0_4_L1_1_Fij_reg_Dout_6 (.Q (FilterDout_4__1__6), .QB (\$dummy [126]), 
        .D (nx2631), .CLK (CLK)) ;
    ao32 ix2632 (.Y (nx2631), .A0 (Din[14]), .A1 (nx8128), .A2 (FilterWR), .B0 (
         FilterDout_4__1__6), .B1 (nx8236)) ;
    dff L0_4_L1_1_Fij_reg_Dout_7 (.Q (FilterDout_4__1__7), .QB (\$dummy [127]), 
        .D (nx2641), .CLK (CLK)) ;
    ao32 ix2642 (.Y (nx2641), .A0 (Din[15]), .A1 (nx8128), .A2 (FilterWR), .B0 (
         FilterDout_4__1__7), .B1 (nx8236)) ;
    dff L0_4_L1_0_Fij_reg_Dout_0 (.Q (FilterDout_4__0__0), .QB (\$dummy [128]), 
        .D (nx2731), .CLK (CLK)) ;
    ao32 ix2732 (.Y (nx2731), .A0 (Din[0]), .A1 (nx8128), .A2 (FilterWR), .B0 (
         FilterDout_4__0__0), .B1 (nx8236)) ;
    dff L0_4_L1_0_Fij_reg_Dout_1 (.Q (FilterDout_4__0__1), .QB (\$dummy [129]), 
        .D (nx2741), .CLK (CLK)) ;
    ao32 ix2742 (.Y (nx2741), .A0 (Din[1]), .A1 (nx8128), .A2 (FilterWR), .B0 (
         FilterDout_4__0__1), .B1 (nx8236)) ;
    dff L0_4_L1_0_Fij_reg_Dout_2 (.Q (FilterDout_4__0__2), .QB (\$dummy [130]), 
        .D (nx2751), .CLK (CLK)) ;
    ao32 ix2752 (.Y (nx2751), .A0 (Din[2]), .A1 (nx8130), .A2 (FilterWR), .B0 (
         FilterDout_4__0__2), .B1 (nx8236)) ;
    dff L0_4_L1_0_Fij_reg_Dout_3 (.Q (FilterDout_4__0__3), .QB (\$dummy [131]), 
        .D (nx2761), .CLK (CLK)) ;
    ao32 ix2762 (.Y (nx2761), .A0 (Din[3]), .A1 (nx8130), .A2 (FilterWR), .B0 (
         FilterDout_4__0__3), .B1 (nx8236)) ;
    dff L0_4_L1_0_Fij_reg_Dout_4 (.Q (FilterDout_4__0__4), .QB (\$dummy [132]), 
        .D (nx2771), .CLK (CLK)) ;
    ao32 ix2772 (.Y (nx2771), .A0 (Din[4]), .A1 (nx8130), .A2 (FilterWR), .B0 (
         FilterDout_4__0__4), .B1 (nx8236)) ;
    dff L0_4_L1_0_Fij_reg_Dout_5 (.Q (FilterDout_4__0__5), .QB (\$dummy [133]), 
        .D (nx2781), .CLK (CLK)) ;
    ao32 ix2782 (.Y (nx2781), .A0 (Din[5]), .A1 (nx8130), .A2 (FilterWR), .B0 (
         FilterDout_4__0__5), .B1 (nx8238)) ;
    dff L0_4_L1_0_Fij_reg_Dout_6 (.Q (FilterDout_4__0__6), .QB (\$dummy [134]), 
        .D (nx2791), .CLK (CLK)) ;
    ao32 ix2792 (.Y (nx2791), .A0 (Din[6]), .A1 (nx8130), .A2 (FilterWR), .B0 (
         FilterDout_4__0__6), .B1 (nx8238)) ;
    dff L0_4_L1_0_Fij_reg_Dout_7 (.Q (FilterDout_4__0__7), .QB (\$dummy [135]), 
        .D (nx2801), .CLK (CLK)) ;
    ao32 ix2802 (.Y (nx2801), .A0 (Din[7]), .A1 (nx8130), .A2 (FilterWR), .B0 (
         FilterDout_4__0__7), .B1 (nx8238)) ;
    oai21 ix2892 (.Y (nx2891), .A0 (nx7122), .A1 (nx8006), .B0 (nx7125)) ;
    dff L0_3_L1_4_Fij_reg_Dout_0 (.Q (FilterDout_3__4__0), .QB (nx7122), .D (
        nx2891), .CLK (CLK)) ;
    nand03 ix7126 (.Y (nx7125), .A0 (nx8130), .A1 (FilterDout_4__4__0), .A2 (
           nx8006)) ;
    oai21 ix2902 (.Y (nx2901), .A0 (nx7129), .A1 (nx8006), .B0 (nx7131)) ;
    dff L0_3_L1_4_Fij_reg_Dout_1 (.Q (FilterDout_3__4__1), .QB (nx7129), .D (
        nx2901), .CLK (CLK)) ;
    nand03 ix7132 (.Y (nx7131), .A0 (nx8132), .A1 (FilterDout_4__4__1), .A2 (
           nx8006)) ;
    oai21 ix2912 (.Y (nx2911), .A0 (nx7135), .A1 (nx8006), .B0 (nx7137)) ;
    dff L0_3_L1_4_Fij_reg_Dout_2 (.Q (FilterDout_3__4__2), .QB (nx7135), .D (
        nx2911), .CLK (CLK)) ;
    nand03 ix7138 (.Y (nx7137), .A0 (nx8132), .A1 (FilterDout_4__4__2), .A2 (
           nx8006)) ;
    oai21 ix2922 (.Y (nx2921), .A0 (nx7141), .A1 (nx8006), .B0 (nx7143)) ;
    dff L0_3_L1_4_Fij_reg_Dout_3 (.Q (FilterDout_3__4__3), .QB (nx7141), .D (
        nx2921), .CLK (CLK)) ;
    nand03 ix7144 (.Y (nx7143), .A0 (nx8132), .A1 (FilterDout_4__4__3), .A2 (
           nx8008)) ;
    oai21 ix2932 (.Y (nx2931), .A0 (nx7147), .A1 (nx8008), .B0 (nx7149)) ;
    dff L0_3_L1_4_Fij_reg_Dout_4 (.Q (FilterDout_3__4__4), .QB (nx7147), .D (
        nx2931), .CLK (CLK)) ;
    nand03 ix7150 (.Y (nx7149), .A0 (nx8132), .A1 (FilterDout_4__4__4), .A2 (
           nx8008)) ;
    oai21 ix2942 (.Y (nx2941), .A0 (nx7153), .A1 (nx8008), .B0 (nx7155)) ;
    dff L0_3_L1_4_Fij_reg_Dout_5 (.Q (FilterDout_3__4__5), .QB (nx7153), .D (
        nx2941), .CLK (CLK)) ;
    nand03 ix7156 (.Y (nx7155), .A0 (nx8132), .A1 (FilterDout_4__4__5), .A2 (
           nx8008)) ;
    oai21 ix2952 (.Y (nx2951), .A0 (nx7159), .A1 (nx8008), .B0 (nx7161)) ;
    dff L0_3_L1_4_Fij_reg_Dout_6 (.Q (FilterDout_3__4__6), .QB (nx7159), .D (
        nx2951), .CLK (CLK)) ;
    nand03 ix7162 (.Y (nx7161), .A0 (nx8132), .A1 (FilterDout_4__4__6), .A2 (
           nx8008)) ;
    oai21 ix2962 (.Y (nx2961), .A0 (nx7165), .A1 (nx8010), .B0 (nx7167)) ;
    dff L0_3_L1_4_Fij_reg_Dout_7 (.Q (FilterDout_3__4__7), .QB (nx7165), .D (
        nx2961), .CLK (CLK)) ;
    nand03 ix7168 (.Y (nx7167), .A0 (nx8132), .A1 (FilterDout_4__4__7), .A2 (
           nx8010)) ;
    oai21 ix3052 (.Y (nx3051), .A0 (nx7171), .A1 (nx8010), .B0 (nx7173)) ;
    dff L0_3_L1_3_Fij_reg_Dout_0 (.Q (FilterDout_3__3__0), .QB (nx7171), .D (
        nx3051), .CLK (CLK)) ;
    nand03 ix7174 (.Y (nx7173), .A0 (nx8134), .A1 (FilterDout_4__3__0), .A2 (
           nx8010)) ;
    oai21 ix3062 (.Y (nx3061), .A0 (nx7177), .A1 (nx8010), .B0 (nx7179)) ;
    dff L0_3_L1_3_Fij_reg_Dout_1 (.Q (FilterDout_3__3__1), .QB (nx7177), .D (
        nx3061), .CLK (CLK)) ;
    nand03 ix7180 (.Y (nx7179), .A0 (nx8134), .A1 (FilterDout_4__3__1), .A2 (
           nx8010)) ;
    oai21 ix3072 (.Y (nx3071), .A0 (nx7183), .A1 (nx8010), .B0 (nx7185)) ;
    dff L0_3_L1_3_Fij_reg_Dout_2 (.Q (FilterDout_3__3__2), .QB (nx7183), .D (
        nx3071), .CLK (CLK)) ;
    nand03 ix7186 (.Y (nx7185), .A0 (nx8134), .A1 (FilterDout_4__3__2), .A2 (
           nx8012)) ;
    oai21 ix3082 (.Y (nx3081), .A0 (nx7189), .A1 (nx8012), .B0 (nx7191)) ;
    dff L0_3_L1_3_Fij_reg_Dout_3 (.Q (FilterDout_3__3__3), .QB (nx7189), .D (
        nx3081), .CLK (CLK)) ;
    nand03 ix7192 (.Y (nx7191), .A0 (nx8134), .A1 (FilterDout_4__3__3), .A2 (
           nx8012)) ;
    oai21 ix3092 (.Y (nx3091), .A0 (nx7195), .A1 (nx8012), .B0 (nx7197)) ;
    dff L0_3_L1_3_Fij_reg_Dout_4 (.Q (FilterDout_3__3__4), .QB (nx7195), .D (
        nx3091), .CLK (CLK)) ;
    nand03 ix7198 (.Y (nx7197), .A0 (nx8134), .A1 (FilterDout_4__3__4), .A2 (
           nx8012)) ;
    oai21 ix3102 (.Y (nx3101), .A0 (nx7201), .A1 (nx8012), .B0 (nx7203)) ;
    dff L0_3_L1_3_Fij_reg_Dout_5 (.Q (FilterDout_3__3__5), .QB (nx7201), .D (
        nx3101), .CLK (CLK)) ;
    nand03 ix7204 (.Y (nx7203), .A0 (nx8134), .A1 (FilterDout_4__3__5), .A2 (
           nx8012)) ;
    oai21 ix3112 (.Y (nx3111), .A0 (nx7207), .A1 (nx8014), .B0 (nx7209)) ;
    dff L0_3_L1_3_Fij_reg_Dout_6 (.Q (FilterDout_3__3__6), .QB (nx7207), .D (
        nx3111), .CLK (CLK)) ;
    nand03 ix7210 (.Y (nx7209), .A0 (nx8134), .A1 (FilterDout_4__3__6), .A2 (
           nx8014)) ;
    oai21 ix3122 (.Y (nx3121), .A0 (nx7213), .A1 (nx8014), .B0 (nx7215)) ;
    dff L0_3_L1_3_Fij_reg_Dout_7 (.Q (FilterDout_3__3__7), .QB (nx7213), .D (
        nx3121), .CLK (CLK)) ;
    nand03 ix7216 (.Y (nx7215), .A0 (nx8136), .A1 (FilterDout_4__3__7), .A2 (
           nx8014)) ;
    dff L0_3_L1_2_Fij_reg_Dout_0 (.Q (FilterDout_3__2__0), .QB (\$dummy [136]), 
        .D (nx3211), .CLK (CLK)) ;
    ao32 ix3212 (.Y (nx3211), .A0 (nx8136), .A1 (FilterDout_4__2__0), .A2 (
         FilterWR), .B0 (FilterDout_3__2__0), .B1 (nx8238)) ;
    dff L0_3_L1_2_Fij_reg_Dout_1 (.Q (FilterDout_3__2__1), .QB (\$dummy [137]), 
        .D (nx3221), .CLK (CLK)) ;
    ao32 ix3222 (.Y (nx3221), .A0 (nx8136), .A1 (FilterDout_4__2__1), .A2 (
         FilterWR), .B0 (FilterDout_3__2__1), .B1 (nx8238)) ;
    dff L0_3_L1_2_Fij_reg_Dout_2 (.Q (FilterDout_3__2__2), .QB (\$dummy [138]), 
        .D (nx3231), .CLK (CLK)) ;
    ao32 ix3232 (.Y (nx3231), .A0 (nx8136), .A1 (FilterDout_4__2__2), .A2 (
         FilterWR), .B0 (FilterDout_3__2__2), .B1 (nx8238)) ;
    dff L0_3_L1_2_Fij_reg_Dout_3 (.Q (FilterDout_3__2__3), .QB (\$dummy [139]), 
        .D (nx3241), .CLK (CLK)) ;
    ao32 ix3242 (.Y (nx3241), .A0 (nx8136), .A1 (FilterDout_4__2__3), .A2 (
         FilterWR), .B0 (FilterDout_3__2__3), .B1 (nx8238)) ;
    dff L0_3_L1_2_Fij_reg_Dout_4 (.Q (FilterDout_3__2__4), .QB (\$dummy [140]), 
        .D (nx3251), .CLK (CLK)) ;
    ao32 ix3252 (.Y (nx3251), .A0 (nx8136), .A1 (FilterDout_4__2__4), .A2 (
         FilterWR), .B0 (FilterDout_3__2__4), .B1 (nx8240)) ;
    dff L0_3_L1_2_Fij_reg_Dout_5 (.Q (FilterDout_3__2__5), .QB (\$dummy [141]), 
        .D (nx3261), .CLK (CLK)) ;
    ao32 ix3262 (.Y (nx3261), .A0 (nx8136), .A1 (FilterDout_4__2__5), .A2 (
         FilterWR), .B0 (FilterDout_3__2__5), .B1 (nx8240)) ;
    dff L0_3_L1_2_Fij_reg_Dout_6 (.Q (FilterDout_3__2__6), .QB (\$dummy [142]), 
        .D (nx3271), .CLK (CLK)) ;
    ao32 ix3272 (.Y (nx3271), .A0 (nx8138), .A1 (FilterDout_4__2__6), .A2 (
         FilterWR), .B0 (FilterDout_3__2__6), .B1 (nx8240)) ;
    dff L0_3_L1_2_Fij_reg_Dout_7 (.Q (FilterDout_3__2__7), .QB (\$dummy [143]), 
        .D (nx3281), .CLK (CLK)) ;
    ao32 ix3282 (.Y (nx3281), .A0 (nx8138), .A1 (FilterDout_4__2__7), .A2 (
         FilterWR), .B0 (FilterDout_3__2__7), .B1 (nx8240)) ;
    dff L0_3_L1_1_Fij_reg_Dout_0 (.Q (FilterDout_3__1__0), .QB (\$dummy [144]), 
        .D (nx3371), .CLK (CLK)) ;
    ao32 ix3372 (.Y (nx3371), .A0 (nx8138), .A1 (FilterDout_4__1__0), .A2 (
         FilterWR), .B0 (FilterDout_3__1__0), .B1 (nx8240)) ;
    dff L0_3_L1_1_Fij_reg_Dout_1 (.Q (FilterDout_3__1__1), .QB (\$dummy [145]), 
        .D (nx3381), .CLK (CLK)) ;
    ao32 ix3382 (.Y (nx3381), .A0 (nx8138), .A1 (FilterDout_4__1__1), .A2 (
         FilterWR), .B0 (FilterDout_3__1__1), .B1 (nx8240)) ;
    dff L0_3_L1_1_Fij_reg_Dout_2 (.Q (FilterDout_3__1__2), .QB (\$dummy [146]), 
        .D (nx3391), .CLK (CLK)) ;
    ao32 ix3392 (.Y (nx3391), .A0 (nx8138), .A1 (FilterDout_4__1__2), .A2 (
         FilterWR), .B0 (FilterDout_3__1__2), .B1 (nx8240)) ;
    dff L0_3_L1_1_Fij_reg_Dout_3 (.Q (FilterDout_3__1__3), .QB (\$dummy [147]), 
        .D (nx3401), .CLK (CLK)) ;
    ao32 ix3402 (.Y (nx3401), .A0 (nx8138), .A1 (FilterDout_4__1__3), .A2 (
         FilterWR), .B0 (FilterDout_3__1__3), .B1 (nx8242)) ;
    dff L0_3_L1_1_Fij_reg_Dout_4 (.Q (FilterDout_3__1__4), .QB (\$dummy [148]), 
        .D (nx3411), .CLK (CLK)) ;
    ao32 ix3412 (.Y (nx3411), .A0 (nx8138), .A1 (FilterDout_4__1__4), .A2 (
         FilterWR), .B0 (FilterDout_3__1__4), .B1 (nx8242)) ;
    dff L0_3_L1_1_Fij_reg_Dout_5 (.Q (FilterDout_3__1__5), .QB (\$dummy [149]), 
        .D (nx3421), .CLK (CLK)) ;
    ao32 ix3422 (.Y (nx3421), .A0 (nx8140), .A1 (FilterDout_4__1__5), .A2 (
         FilterWR), .B0 (FilterDout_3__1__5), .B1 (nx8242)) ;
    dff L0_3_L1_1_Fij_reg_Dout_6 (.Q (FilterDout_3__1__6), .QB (\$dummy [150]), 
        .D (nx3431), .CLK (CLK)) ;
    ao32 ix3432 (.Y (nx3431), .A0 (nx8140), .A1 (FilterDout_4__1__6), .A2 (
         FilterWR), .B0 (FilterDout_3__1__6), .B1 (nx8242)) ;
    dff L0_3_L1_1_Fij_reg_Dout_7 (.Q (FilterDout_3__1__7), .QB (\$dummy [151]), 
        .D (nx3441), .CLK (CLK)) ;
    ao32 ix3442 (.Y (nx3441), .A0 (nx8140), .A1 (FilterDout_4__1__7), .A2 (
         FilterWR), .B0 (FilterDout_3__1__7), .B1 (nx8242)) ;
    dff L0_3_L1_0_Fij_reg_Dout_0 (.Q (FilterDout_3__0__0), .QB (\$dummy [152]), 
        .D (nx3531), .CLK (CLK)) ;
    ao32 ix3532 (.Y (nx3531), .A0 (nx8140), .A1 (FilterDout_4__0__0), .A2 (
         FilterWR), .B0 (FilterDout_3__0__0), .B1 (nx8242)) ;
    dff L0_3_L1_0_Fij_reg_Dout_1 (.Q (FilterDout_3__0__1), .QB (\$dummy [153]), 
        .D (nx3541), .CLK (CLK)) ;
    ao32 ix3542 (.Y (nx3541), .A0 (nx8140), .A1 (FilterDout_4__0__1), .A2 (
         FilterWR), .B0 (FilterDout_3__0__1), .B1 (nx8242)) ;
    dff L0_3_L1_0_Fij_reg_Dout_2 (.Q (FilterDout_3__0__2), .QB (\$dummy [154]), 
        .D (nx3551), .CLK (CLK)) ;
    ao32 ix3552 (.Y (nx3551), .A0 (nx8140), .A1 (FilterDout_4__0__2), .A2 (
         FilterWR), .B0 (FilterDout_3__0__2), .B1 (nx8244)) ;
    dff L0_3_L1_0_Fij_reg_Dout_3 (.Q (FilterDout_3__0__3), .QB (\$dummy [155]), 
        .D (nx3561), .CLK (CLK)) ;
    ao32 ix3562 (.Y (nx3561), .A0 (nx8140), .A1 (FilterDout_4__0__3), .A2 (
         FilterWR), .B0 (FilterDout_3__0__3), .B1 (nx8244)) ;
    dff L0_3_L1_0_Fij_reg_Dout_4 (.Q (FilterDout_3__0__4), .QB (\$dummy [156]), 
        .D (nx3571), .CLK (CLK)) ;
    ao32 ix3572 (.Y (nx3571), .A0 (nx8142), .A1 (FilterDout_4__0__4), .A2 (
         FilterWR), .B0 (FilterDout_3__0__4), .B1 (nx8244)) ;
    dff L0_3_L1_0_Fij_reg_Dout_5 (.Q (FilterDout_3__0__5), .QB (\$dummy [157]), 
        .D (nx3581), .CLK (CLK)) ;
    ao32 ix3582 (.Y (nx3581), .A0 (nx8142), .A1 (FilterDout_4__0__5), .A2 (
         FilterWR), .B0 (FilterDout_3__0__5), .B1 (nx8244)) ;
    dff L0_3_L1_0_Fij_reg_Dout_6 (.Q (FilterDout_3__0__6), .QB (\$dummy [158]), 
        .D (nx3591), .CLK (CLK)) ;
    ao32 ix3592 (.Y (nx3591), .A0 (nx8142), .A1 (FilterDout_4__0__6), .A2 (
         FilterWR), .B0 (FilterDout_3__0__6), .B1 (nx8244)) ;
    dff L0_3_L1_0_Fij_reg_Dout_7 (.Q (FilterDout_3__0__7), .QB (\$dummy [159]), 
        .D (nx3601), .CLK (CLK)) ;
    ao32 ix3602 (.Y (nx3601), .A0 (nx8142), .A1 (FilterDout_4__0__7), .A2 (
         FilterWR), .B0 (FilterDout_3__0__7), .B1 (nx8244)) ;
    oai21 ix3692 (.Y (nx3691), .A0 (nx7291), .A1 (nx8014), .B0 (nx7293)) ;
    dff L0_2_L1_4_Fij_reg_Dout_0 (.Q (FilterDout_2__4__0), .QB (nx7291), .D (
        nx3691), .CLK (CLK)) ;
    oai21 ix3702 (.Y (nx3701), .A0 (nx7297), .A1 (nx8014), .B0 (nx7299)) ;
    dff L0_2_L1_4_Fij_reg_Dout_1 (.Q (FilterDout_2__4__1), .QB (nx7297), .D (
        nx3701), .CLK (CLK)) ;
    oai21 ix3712 (.Y (nx3711), .A0 (nx7303), .A1 (nx8016), .B0 (nx7305)) ;
    dff L0_2_L1_4_Fij_reg_Dout_2 (.Q (FilterDout_2__4__2), .QB (nx7303), .D (
        nx3711), .CLK (CLK)) ;
    oai21 ix3722 (.Y (nx3721), .A0 (nx7309), .A1 (nx8016), .B0 (nx7311)) ;
    dff L0_2_L1_4_Fij_reg_Dout_3 (.Q (FilterDout_2__4__3), .QB (nx7309), .D (
        nx3721), .CLK (CLK)) ;
    oai21 ix3732 (.Y (nx3731), .A0 (nx7315), .A1 (nx8016), .B0 (nx7317)) ;
    dff L0_2_L1_4_Fij_reg_Dout_4 (.Q (FilterDout_2__4__4), .QB (nx7315), .D (
        nx3731), .CLK (CLK)) ;
    oai21 ix3742 (.Y (nx3741), .A0 (nx7321), .A1 (nx8018), .B0 (nx7323)) ;
    dff L0_2_L1_4_Fij_reg_Dout_5 (.Q (FilterDout_2__4__5), .QB (nx7321), .D (
        nx3741), .CLK (CLK)) ;
    oai21 ix3752 (.Y (nx3751), .A0 (nx7327), .A1 (nx8018), .B0 (nx7329)) ;
    dff L0_2_L1_4_Fij_reg_Dout_6 (.Q (FilterDout_2__4__6), .QB (nx7327), .D (
        nx3751), .CLK (CLK)) ;
    oai21 ix3762 (.Y (nx3761), .A0 (nx7333), .A1 (nx8018), .B0 (nx7335)) ;
    dff L0_2_L1_4_Fij_reg_Dout_7 (.Q (FilterDout_2__4__7), .QB (nx7333), .D (
        nx3761), .CLK (CLK)) ;
    oai21 ix3852 (.Y (nx3851), .A0 (nx7339), .A1 (nx8018), .B0 (nx7341)) ;
    dff L0_2_L1_3_Fij_reg_Dout_0 (.Q (FilterDout_2__3__0), .QB (nx7339), .D (
        nx3851), .CLK (CLK)) ;
    oai21 ix3862 (.Y (nx3861), .A0 (nx7345), .A1 (nx8020), .B0 (nx7347)) ;
    dff L0_2_L1_3_Fij_reg_Dout_1 (.Q (FilterDout_2__3__1), .QB (nx7345), .D (
        nx3861), .CLK (CLK)) ;
    oai21 ix3872 (.Y (nx3871), .A0 (nx7351), .A1 (nx8020), .B0 (nx7353)) ;
    dff L0_2_L1_3_Fij_reg_Dout_2 (.Q (FilterDout_2__3__2), .QB (nx7351), .D (
        nx3871), .CLK (CLK)) ;
    oai21 ix3882 (.Y (nx3881), .A0 (nx7357), .A1 (nx8020), .B0 (nx7359)) ;
    dff L0_2_L1_3_Fij_reg_Dout_3 (.Q (FilterDout_2__3__3), .QB (nx7357), .D (
        nx3881), .CLK (CLK)) ;
    oai21 ix3892 (.Y (nx3891), .A0 (nx7363), .A1 (nx8022), .B0 (nx7365)) ;
    dff L0_2_L1_3_Fij_reg_Dout_4 (.Q (FilterDout_2__3__4), .QB (nx7363), .D (
        nx3891), .CLK (CLK)) ;
    oai21 ix3902 (.Y (nx3901), .A0 (nx7369), .A1 (nx8022), .B0 (nx7371)) ;
    dff L0_2_L1_3_Fij_reg_Dout_5 (.Q (FilterDout_2__3__5), .QB (nx7369), .D (
        nx3901), .CLK (CLK)) ;
    oai21 ix3912 (.Y (nx3911), .A0 (nx7375), .A1 (nx8022), .B0 (nx7377)) ;
    dff L0_2_L1_3_Fij_reg_Dout_6 (.Q (FilterDout_2__3__6), .QB (nx7375), .D (
        nx3911), .CLK (CLK)) ;
    oai21 ix3922 (.Y (nx3921), .A0 (nx7381), .A1 (nx8022), .B0 (nx7383)) ;
    dff L0_2_L1_3_Fij_reg_Dout_7 (.Q (FilterDout_2__3__7), .QB (nx7381), .D (
        nx3921), .CLK (CLK)) ;
    dff L0_2_L1_2_Fij_reg_Dout_0 (.Q (FilterDout_2__2__0), .QB (\$dummy [160]), 
        .D (nx4011), .CLK (CLK)) ;
    ao32 ix4012 (.Y (nx4011), .A0 (nx8146), .A1 (FilterDout_3__2__0), .A2 (
         FilterWR), .B0 (FilterDout_2__2__0), .B1 (nx8244)) ;
    dff L0_2_L1_2_Fij_reg_Dout_1 (.Q (FilterDout_2__2__1), .QB (\$dummy [161]), 
        .D (nx4021), .CLK (CLK)) ;
    ao32 ix4022 (.Y (nx4021), .A0 (nx8148), .A1 (FilterDout_3__2__1), .A2 (
         FilterWR), .B0 (FilterDout_2__2__1), .B1 (nx8246)) ;
    dff L0_2_L1_2_Fij_reg_Dout_2 (.Q (FilterDout_2__2__2), .QB (\$dummy [162]), 
        .D (nx4031), .CLK (CLK)) ;
    ao32 ix4032 (.Y (nx4031), .A0 (nx8148), .A1 (FilterDout_3__2__2), .A2 (
         FilterWR), .B0 (FilterDout_2__2__2), .B1 (nx8246)) ;
    dff L0_2_L1_2_Fij_reg_Dout_3 (.Q (FilterDout_2__2__3), .QB (\$dummy [163]), 
        .D (nx4041), .CLK (CLK)) ;
    ao32 ix4042 (.Y (nx4041), .A0 (nx8148), .A1 (FilterDout_3__2__3), .A2 (
         FilterWR), .B0 (FilterDout_2__2__3), .B1 (nx8246)) ;
    dff L0_2_L1_2_Fij_reg_Dout_4 (.Q (FilterDout_2__2__4), .QB (\$dummy [164]), 
        .D (nx4051), .CLK (CLK)) ;
    ao32 ix4052 (.Y (nx4051), .A0 (nx8148), .A1 (FilterDout_3__2__4), .A2 (
         FilterWR), .B0 (FilterDout_2__2__4), .B1 (nx8246)) ;
    dff L0_2_L1_2_Fij_reg_Dout_5 (.Q (FilterDout_2__2__5), .QB (\$dummy [165]), 
        .D (nx4061), .CLK (CLK)) ;
    ao32 ix4062 (.Y (nx4061), .A0 (nx8148), .A1 (FilterDout_3__2__5), .A2 (
         FilterWR), .B0 (FilterDout_2__2__5), .B1 (nx8246)) ;
    dff L0_2_L1_2_Fij_reg_Dout_6 (.Q (FilterDout_2__2__6), .QB (\$dummy [166]), 
        .D (nx4071), .CLK (CLK)) ;
    ao32 ix4072 (.Y (nx4071), .A0 (nx8148), .A1 (FilterDout_3__2__6), .A2 (
         FilterWR), .B0 (FilterDout_2__2__6), .B1 (nx8246)) ;
    dff L0_2_L1_2_Fij_reg_Dout_7 (.Q (FilterDout_2__2__7), .QB (\$dummy [167]), 
        .D (nx4081), .CLK (CLK)) ;
    ao32 ix4082 (.Y (nx4081), .A0 (nx8148), .A1 (FilterDout_3__2__7), .A2 (
         FilterWR), .B0 (FilterDout_2__2__7), .B1 (nx8246)) ;
    dff L0_2_L1_1_Fij_reg_Dout_0 (.Q (FilterDout_2__1__0), .QB (\$dummy [168]), 
        .D (nx4171), .CLK (CLK)) ;
    ao32 ix4172 (.Y (nx4171), .A0 (nx8150), .A1 (FilterDout_3__1__0), .A2 (
         FilterWR), .B0 (FilterDout_2__1__0), .B1 (nx8248)) ;
    dff L0_2_L1_1_Fij_reg_Dout_1 (.Q (FilterDout_2__1__1), .QB (\$dummy [169]), 
        .D (nx4181), .CLK (CLK)) ;
    ao32 ix4182 (.Y (nx4181), .A0 (nx8150), .A1 (FilterDout_3__1__1), .A2 (
         FilterWR), .B0 (FilterDout_2__1__1), .B1 (nx8248)) ;
    dff L0_2_L1_1_Fij_reg_Dout_2 (.Q (FilterDout_2__1__2), .QB (\$dummy [170]), 
        .D (nx4191), .CLK (CLK)) ;
    ao32 ix4192 (.Y (nx4191), .A0 (nx8150), .A1 (FilterDout_3__1__2), .A2 (
         FilterWR), .B0 (FilterDout_2__1__2), .B1 (nx8248)) ;
    dff L0_2_L1_1_Fij_reg_Dout_3 (.Q (FilterDout_2__1__3), .QB (\$dummy [171]), 
        .D (nx4201), .CLK (CLK)) ;
    ao32 ix4202 (.Y (nx4201), .A0 (nx8150), .A1 (FilterDout_3__1__3), .A2 (
         FilterWR), .B0 (FilterDout_2__1__3), .B1 (nx8248)) ;
    dff L0_2_L1_1_Fij_reg_Dout_4 (.Q (FilterDout_2__1__4), .QB (\$dummy [172]), 
        .D (nx4211), .CLK (CLK)) ;
    ao32 ix4212 (.Y (nx4211), .A0 (nx8150), .A1 (FilterDout_3__1__4), .A2 (
         FilterWR), .B0 (FilterDout_2__1__4), .B1 (nx8248)) ;
    dff L0_2_L1_1_Fij_reg_Dout_5 (.Q (FilterDout_2__1__5), .QB (\$dummy [173]), 
        .D (nx4221), .CLK (CLK)) ;
    ao32 ix4222 (.Y (nx4221), .A0 (nx8150), .A1 (FilterDout_3__1__5), .A2 (
         FilterWR), .B0 (FilterDout_2__1__5), .B1 (nx8248)) ;
    dff L0_2_L1_1_Fij_reg_Dout_6 (.Q (FilterDout_2__1__6), .QB (\$dummy [174]), 
        .D (nx4231), .CLK (CLK)) ;
    ao32 ix4232 (.Y (nx4231), .A0 (nx8150), .A1 (FilterDout_3__1__6), .A2 (
         FilterWR), .B0 (FilterDout_2__1__6), .B1 (nx8248)) ;
    dff L0_2_L1_1_Fij_reg_Dout_7 (.Q (FilterDout_2__1__7), .QB (\$dummy [175]), 
        .D (nx4241), .CLK (CLK)) ;
    ao32 ix4242 (.Y (nx4241), .A0 (nx8152), .A1 (FilterDout_3__1__7), .A2 (
         FilterWR), .B0 (FilterDout_2__1__7), .B1 (nx8250)) ;
    dff L0_2_L1_0_Fij_reg_Dout_0 (.Q (FilterDout_2__0__0), .QB (\$dummy [176]), 
        .D (nx4331), .CLK (CLK)) ;
    ao32 ix4332 (.Y (nx4331), .A0 (nx8152), .A1 (FilterDout_3__0__0), .A2 (
         FilterWR), .B0 (FilterDout_2__0__0), .B1 (nx8250)) ;
    dff L0_2_L1_0_Fij_reg_Dout_1 (.Q (FilterDout_2__0__1), .QB (\$dummy [177]), 
        .D (nx4341), .CLK (CLK)) ;
    ao32 ix4342 (.Y (nx4341), .A0 (nx8152), .A1 (FilterDout_3__0__1), .A2 (
         FilterWR), .B0 (FilterDout_2__0__1), .B1 (nx8250)) ;
    dff L0_2_L1_0_Fij_reg_Dout_2 (.Q (FilterDout_2__0__2), .QB (\$dummy [178]), 
        .D (nx4351), .CLK (CLK)) ;
    ao32 ix4352 (.Y (nx4351), .A0 (nx8152), .A1 (FilterDout_3__0__2), .A2 (
         FilterWR), .B0 (FilterDout_2__0__2), .B1 (nx8250)) ;
    dff L0_2_L1_0_Fij_reg_Dout_3 (.Q (FilterDout_2__0__3), .QB (\$dummy [179]), 
        .D (nx4361), .CLK (CLK)) ;
    ao32 ix4362 (.Y (nx4361), .A0 (nx8152), .A1 (FilterDout_3__0__3), .A2 (
         FilterWR), .B0 (FilterDout_2__0__3), .B1 (nx8250)) ;
    dff L0_2_L1_0_Fij_reg_Dout_4 (.Q (FilterDout_2__0__4), .QB (\$dummy [180]), 
        .D (nx4371), .CLK (CLK)) ;
    ao32 ix4372 (.Y (nx4371), .A0 (nx8152), .A1 (FilterDout_3__0__4), .A2 (
         FilterWR), .B0 (FilterDout_2__0__4), .B1 (nx8250)) ;
    dff L0_2_L1_0_Fij_reg_Dout_5 (.Q (FilterDout_2__0__5), .QB (\$dummy [181]), 
        .D (nx4381), .CLK (CLK)) ;
    ao32 ix4382 (.Y (nx4381), .A0 (nx8152), .A1 (FilterDout_3__0__5), .A2 (
         FilterWR), .B0 (FilterDout_2__0__5), .B1 (nx8250)) ;
    dff L0_2_L1_0_Fij_reg_Dout_6 (.Q (FilterDout_2__0__6), .QB (\$dummy [182]), 
        .D (nx4391), .CLK (CLK)) ;
    ao32 ix4392 (.Y (nx4391), .A0 (nx8154), .A1 (FilterDout_3__0__6), .A2 (
         FilterWR), .B0 (FilterDout_2__0__6), .B1 (nx8252)) ;
    dff L0_2_L1_0_Fij_reg_Dout_7 (.Q (FilterDout_2__0__7), .QB (\$dummy [183]), 
        .D (nx4401), .CLK (CLK)) ;
    ao32 ix4402 (.Y (nx4401), .A0 (nx8154), .A1 (FilterDout_3__0__7), .A2 (
         FilterWR), .B0 (FilterDout_2__0__7), .B1 (nx8252)) ;
    oai21 ix4572 (.Y (nx4571), .A0 (nx7459), .A1 (nx8024), .B0 (nx7461)) ;
    dff L0_1_L1_4_Fij_reg_Dout_0 (.Q (FilterDout_1__4__0), .QB (nx7459), .D (
        nx4571), .CLK (CLK)) ;
    oai21 ix4582 (.Y (nx4581), .A0 (nx7465), .A1 (nx8024), .B0 (nx7467)) ;
    dff L0_1_L1_4_Fij_reg_Dout_1 (.Q (FilterDout_1__4__1), .QB (nx7465), .D (
        nx4581), .CLK (CLK)) ;
    oai21 ix4592 (.Y (nx4591), .A0 (nx7471), .A1 (nx8024), .B0 (nx7473)) ;
    dff L0_1_L1_4_Fij_reg_Dout_2 (.Q (FilterDout_1__4__2), .QB (nx7471), .D (
        nx4591), .CLK (CLK)) ;
    oai21 ix4602 (.Y (nx4601), .A0 (nx7477), .A1 (nx8026), .B0 (nx7479)) ;
    dff L0_1_L1_4_Fij_reg_Dout_3 (.Q (FilterDout_1__4__3), .QB (nx7477), .D (
        nx4601), .CLK (CLK)) ;
    oai21 ix4612 (.Y (nx4611), .A0 (nx7483), .A1 (nx8026), .B0 (nx7485)) ;
    dff L0_1_L1_4_Fij_reg_Dout_4 (.Q (FilterDout_1__4__4), .QB (nx7483), .D (
        nx4611), .CLK (CLK)) ;
    oai21 ix4622 (.Y (nx4621), .A0 (nx7489), .A1 (nx8026), .B0 (nx7491)) ;
    dff L0_1_L1_4_Fij_reg_Dout_5 (.Q (FilterDout_1__4__5), .QB (nx7489), .D (
        nx4621), .CLK (CLK)) ;
    oai21 ix4632 (.Y (nx4631), .A0 (nx7495), .A1 (nx8026), .B0 (nx7497)) ;
    dff L0_1_L1_4_Fij_reg_Dout_6 (.Q (FilterDout_1__4__6), .QB (nx7495), .D (
        nx4631), .CLK (CLK)) ;
    oai21 ix4642 (.Y (nx4641), .A0 (nx7501), .A1 (nx8028), .B0 (nx7503)) ;
    dff L0_1_L1_4_Fij_reg_Dout_7 (.Q (FilterDout_1__4__7), .QB (nx7501), .D (
        nx4641), .CLK (CLK)) ;
    oai21 ix4892 (.Y (nx4891), .A0 (nx7507), .A1 (nx8028), .B0 (nx7509)) ;
    dff L0_1_L1_3_Fij_reg_Dout_0 (.Q (FilterDout_1__3__0), .QB (nx7507), .D (
        nx4891), .CLK (CLK)) ;
    oai21 ix4902 (.Y (nx4901), .A0 (nx7513), .A1 (nx8028), .B0 (nx7515)) ;
    dff L0_1_L1_3_Fij_reg_Dout_1 (.Q (FilterDout_1__3__1), .QB (nx7513), .D (
        nx4901), .CLK (CLK)) ;
    oai21 ix4912 (.Y (nx4911), .A0 (nx7519), .A1 (nx8030), .B0 (nx7521)) ;
    dff L0_1_L1_3_Fij_reg_Dout_2 (.Q (FilterDout_1__3__2), .QB (nx7519), .D (
        nx4911), .CLK (CLK)) ;
    oai21 ix4922 (.Y (nx4921), .A0 (nx7525), .A1 (nx8030), .B0 (nx7527)) ;
    dff L0_1_L1_3_Fij_reg_Dout_3 (.Q (FilterDout_1__3__3), .QB (nx7525), .D (
        nx4921), .CLK (CLK)) ;
    oai21 ix4932 (.Y (nx4931), .A0 (nx7531), .A1 (nx8030), .B0 (nx7533)) ;
    dff L0_1_L1_3_Fij_reg_Dout_4 (.Q (FilterDout_1__3__4), .QB (nx7531), .D (
        nx4931), .CLK (CLK)) ;
    oai21 ix4942 (.Y (nx4941), .A0 (nx7537), .A1 (nx8030), .B0 (nx7539)) ;
    dff L0_1_L1_3_Fij_reg_Dout_5 (.Q (FilterDout_1__3__5), .QB (nx7537), .D (
        nx4941), .CLK (CLK)) ;
    oai21 ix4952 (.Y (nx4951), .A0 (nx7543), .A1 (nx8032), .B0 (nx7545)) ;
    dff L0_1_L1_3_Fij_reg_Dout_6 (.Q (FilterDout_1__3__6), .QB (nx7543), .D (
        nx4951), .CLK (CLK)) ;
    oai21 ix4962 (.Y (nx4961), .A0 (nx7549), .A1 (nx8032), .B0 (nx7551)) ;
    dff L0_1_L1_3_Fij_reg_Dout_7 (.Q (FilterDout_1__3__7), .QB (nx7549), .D (
        nx4961), .CLK (CLK)) ;
    oai21 ix5212 (.Y (nx5211), .A0 (nx7555), .A1 (nx8032), .B0 (nx7557)) ;
    dff L0_1_L1_2_Fij_reg_Dout_0 (.Q (FilterDout_1__2__0), .QB (nx7555), .D (
        nx5211), .CLK (CLK)) ;
    nand03 ix7558 (.Y (nx7557), .A0 (nx8158), .A1 (FilterDout_2__2__0), .A2 (
           nx8032)) ;
    oai21 ix5222 (.Y (nx5221), .A0 (nx7561), .A1 (nx8034), .B0 (nx7563)) ;
    dff L0_1_L1_2_Fij_reg_Dout_1 (.Q (FilterDout_1__2__1), .QB (nx7561), .D (
        nx5221), .CLK (CLK)) ;
    nand03 ix7564 (.Y (nx7563), .A0 (nx8158), .A1 (FilterDout_2__2__1), .A2 (
           nx8034)) ;
    oai21 ix5232 (.Y (nx5231), .A0 (nx7567), .A1 (nx8034), .B0 (nx7569)) ;
    dff L0_1_L1_2_Fij_reg_Dout_2 (.Q (FilterDout_1__2__2), .QB (nx7567), .D (
        nx5231), .CLK (CLK)) ;
    nand03 ix7570 (.Y (nx7569), .A0 (nx8158), .A1 (FilterDout_2__2__2), .A2 (
           nx8034)) ;
    oai21 ix5242 (.Y (nx5241), .A0 (nx7573), .A1 (nx8034), .B0 (nx7575)) ;
    dff L0_1_L1_2_Fij_reg_Dout_3 (.Q (FilterDout_1__2__3), .QB (nx7573), .D (
        nx5241), .CLK (CLK)) ;
    nand03 ix7576 (.Y (nx7575), .A0 (nx8160), .A1 (FilterDout_2__2__3), .A2 (
           nx8034)) ;
    oai21 ix5252 (.Y (nx5251), .A0 (nx7579), .A1 (nx8034), .B0 (nx7581)) ;
    dff L0_1_L1_2_Fij_reg_Dout_4 (.Q (FilterDout_1__2__4), .QB (nx7579), .D (
        nx5251), .CLK (CLK)) ;
    nand03 ix7582 (.Y (nx7581), .A0 (nx8160), .A1 (FilterDout_2__2__4), .A2 (
           nx8036)) ;
    oai21 ix5262 (.Y (nx5261), .A0 (nx7585), .A1 (nx8036), .B0 (nx7587)) ;
    dff L0_1_L1_2_Fij_reg_Dout_5 (.Q (FilterDout_1__2__5), .QB (nx7585), .D (
        nx5261), .CLK (CLK)) ;
    nand03 ix7588 (.Y (nx7587), .A0 (nx8160), .A1 (FilterDout_2__2__5), .A2 (
           nx8036)) ;
    oai21 ix5272 (.Y (nx5271), .A0 (nx7591), .A1 (nx8036), .B0 (nx7593)) ;
    dff L0_1_L1_2_Fij_reg_Dout_6 (.Q (FilterDout_1__2__6), .QB (nx7591), .D (
        nx5271), .CLK (CLK)) ;
    nand03 ix7594 (.Y (nx7593), .A0 (nx8160), .A1 (FilterDout_2__2__6), .A2 (
           nx8036)) ;
    oai21 ix5282 (.Y (nx5281), .A0 (nx7597), .A1 (nx8036), .B0 (nx7599)) ;
    dff L0_1_L1_2_Fij_reg_Dout_7 (.Q (FilterDout_1__2__7), .QB (nx7597), .D (
        nx5281), .CLK (CLK)) ;
    nand03 ix7600 (.Y (nx7599), .A0 (nx8160), .A1 (FilterDout_2__2__7), .A2 (
           nx8036)) ;
    oai21 ix5532 (.Y (nx5531), .A0 (nx7603), .A1 (nx8038), .B0 (nx7605)) ;
    dff L0_1_L1_1_Fij_reg_Dout_0 (.Q (FilterDout_1__1__0), .QB (nx7603), .D (
        nx5531), .CLK (CLK)) ;
    nand03 ix7606 (.Y (nx7605), .A0 (nx8160), .A1 (FilterDout_2__1__0), .A2 (
           nx8038)) ;
    oai21 ix5542 (.Y (nx5541), .A0 (nx7609), .A1 (nx8038), .B0 (nx7611)) ;
    dff L0_1_L1_1_Fij_reg_Dout_1 (.Q (FilterDout_1__1__1), .QB (nx7609), .D (
        nx5541), .CLK (CLK)) ;
    nand03 ix7612 (.Y (nx7611), .A0 (nx8160), .A1 (FilterDout_2__1__1), .A2 (
           nx8038)) ;
    oai21 ix5552 (.Y (nx5551), .A0 (nx7615), .A1 (nx8038), .B0 (nx7617)) ;
    dff L0_1_L1_1_Fij_reg_Dout_2 (.Q (FilterDout_1__1__2), .QB (nx7615), .D (
        nx5551), .CLK (CLK)) ;
    nand03 ix7618 (.Y (nx7617), .A0 (nx8162), .A1 (FilterDout_2__1__2), .A2 (
           nx8038)) ;
    oai21 ix5562 (.Y (nx5561), .A0 (nx7621), .A1 (nx8038), .B0 (nx7623)) ;
    dff L0_1_L1_1_Fij_reg_Dout_3 (.Q (FilterDout_1__1__3), .QB (nx7621), .D (
        nx5561), .CLK (CLK)) ;
    nand03 ix7624 (.Y (nx7623), .A0 (nx8162), .A1 (FilterDout_2__1__3), .A2 (
           nx8040)) ;
    oai21 ix5572 (.Y (nx5571), .A0 (nx7627), .A1 (nx8040), .B0 (nx7629)) ;
    dff L0_1_L1_1_Fij_reg_Dout_4 (.Q (FilterDout_1__1__4), .QB (nx7627), .D (
        nx5571), .CLK (CLK)) ;
    nand03 ix7630 (.Y (nx7629), .A0 (nx8162), .A1 (FilterDout_2__1__4), .A2 (
           nx8040)) ;
    oai21 ix5582 (.Y (nx5581), .A0 (nx7633), .A1 (nx8040), .B0 (nx7635)) ;
    dff L0_1_L1_1_Fij_reg_Dout_5 (.Q (FilterDout_1__1__5), .QB (nx7633), .D (
        nx5581), .CLK (CLK)) ;
    nand03 ix7636 (.Y (nx7635), .A0 (nx8162), .A1 (FilterDout_2__1__5), .A2 (
           nx8040)) ;
    oai21 ix5592 (.Y (nx5591), .A0 (nx7639), .A1 (nx8040), .B0 (nx7641)) ;
    dff L0_1_L1_1_Fij_reg_Dout_6 (.Q (FilterDout_1__1__6), .QB (nx7639), .D (
        nx5591), .CLK (CLK)) ;
    nand03 ix7642 (.Y (nx7641), .A0 (nx8162), .A1 (FilterDout_2__1__6), .A2 (
           nx8040)) ;
    oai21 ix5602 (.Y (nx5601), .A0 (nx7645), .A1 (nx8042), .B0 (nx7647)) ;
    dff L0_1_L1_1_Fij_reg_Dout_7 (.Q (FilterDout_1__1__7), .QB (nx7645), .D (
        nx5601), .CLK (CLK)) ;
    nand03 ix7648 (.Y (nx7647), .A0 (nx8162), .A1 (FilterDout_2__1__7), .A2 (
           nx8042)) ;
    oai21 ix5852 (.Y (nx5851), .A0 (nx7651), .A1 (nx8042), .B0 (nx7653)) ;
    dff L0_1_L1_0_Fij_reg_Dout_0 (.Q (FilterDout_1__0__0), .QB (nx7651), .D (
        nx5851), .CLK (CLK)) ;
    nand03 ix7654 (.Y (nx7653), .A0 (nx8162), .A1 (FilterDout_2__0__0), .A2 (
           nx8042)) ;
    oai21 ix5862 (.Y (nx5861), .A0 (nx7657), .A1 (nx8042), .B0 (nx7659)) ;
    dff L0_1_L1_0_Fij_reg_Dout_1 (.Q (FilterDout_1__0__1), .QB (nx7657), .D (
        nx5861), .CLK (CLK)) ;
    nand03 ix7660 (.Y (nx7659), .A0 (nx8164), .A1 (FilterDout_2__0__1), .A2 (
           nx8042)) ;
    oai21 ix5872 (.Y (nx5871), .A0 (nx7663), .A1 (nx8042), .B0 (nx7665)) ;
    dff L0_1_L1_0_Fij_reg_Dout_2 (.Q (FilterDout_1__0__2), .QB (nx7663), .D (
        nx5871), .CLK (CLK)) ;
    nand03 ix7666 (.Y (nx7665), .A0 (nx8164), .A1 (FilterDout_2__0__2), .A2 (
           nx8044)) ;
    oai21 ix5882 (.Y (nx5881), .A0 (nx7669), .A1 (nx8044), .B0 (nx7671)) ;
    dff L0_1_L1_0_Fij_reg_Dout_3 (.Q (FilterDout_1__0__3), .QB (nx7669), .D (
        nx5881), .CLK (CLK)) ;
    nand03 ix7672 (.Y (nx7671), .A0 (nx8164), .A1 (FilterDout_2__0__3), .A2 (
           nx8044)) ;
    oai21 ix5892 (.Y (nx5891), .A0 (nx7675), .A1 (nx8044), .B0 (nx7677)) ;
    dff L0_1_L1_0_Fij_reg_Dout_4 (.Q (FilterDout_1__0__4), .QB (nx7675), .D (
        nx5891), .CLK (CLK)) ;
    nand03 ix7678 (.Y (nx7677), .A0 (nx8164), .A1 (FilterDout_2__0__4), .A2 (
           nx8044)) ;
    oai21 ix5902 (.Y (nx5901), .A0 (nx7681), .A1 (nx8044), .B0 (nx7683)) ;
    dff L0_1_L1_0_Fij_reg_Dout_5 (.Q (FilterDout_1__0__5), .QB (nx7681), .D (
        nx5901), .CLK (CLK)) ;
    nand03 ix7684 (.Y (nx7683), .A0 (nx8164), .A1 (FilterDout_2__0__5), .A2 (
           nx8044)) ;
    oai21 ix5912 (.Y (nx5911), .A0 (nx7687), .A1 (nx8046), .B0 (nx7689)) ;
    dff L0_1_L1_0_Fij_reg_Dout_6 (.Q (FilterDout_1__0__6), .QB (nx7687), .D (
        nx5911), .CLK (CLK)) ;
    nand03 ix7690 (.Y (nx7689), .A0 (nx8164), .A1 (FilterDout_2__0__6), .A2 (
           nx8046)) ;
    oai21 ix5922 (.Y (nx5921), .A0 (nx7693), .A1 (nx8046), .B0 (nx7695)) ;
    dff L0_1_L1_0_Fij_reg_Dout_7 (.Q (FilterDout_1__0__7), .QB (nx7693), .D (
        nx5921), .CLK (CLK)) ;
    nand03 ix7696 (.Y (nx7695), .A0 (nx8164), .A1 (FilterDout_2__0__7), .A2 (
           nx8046)) ;
    oai21 ix4652 (.Y (nx4651), .A0 (nx7699), .A1 (nx8046), .B0 (nx7701)) ;
    dff L0_0_L1_4_Fij_reg_Dout_0 (.Q (FilterDout_0__4__0), .QB (nx7699), .D (
        nx4651), .CLK (CLK)) ;
    oai21 ix4662 (.Y (nx4661), .A0 (nx7705), .A1 (nx8046), .B0 (nx7707)) ;
    dff L0_0_L1_4_Fij_reg_Dout_1 (.Q (FilterDout_0__4__1), .QB (nx7705), .D (
        nx4661), .CLK (CLK)) ;
    oai21 ix4672 (.Y (nx4671), .A0 (nx7711), .A1 (nx8048), .B0 (nx7713)) ;
    dff L0_0_L1_4_Fij_reg_Dout_2 (.Q (FilterDout_0__4__2), .QB (nx7711), .D (
        nx4671), .CLK (CLK)) ;
    oai21 ix4682 (.Y (nx4681), .A0 (nx7717), .A1 (nx8048), .B0 (nx7719)) ;
    dff L0_0_L1_4_Fij_reg_Dout_3 (.Q (FilterDout_0__4__3), .QB (nx7717), .D (
        nx4681), .CLK (CLK)) ;
    oai21 ix4692 (.Y (nx4691), .A0 (nx7723), .A1 (nx8048), .B0 (nx7725)) ;
    dff L0_0_L1_4_Fij_reg_Dout_4 (.Q (FilterDout_0__4__4), .QB (nx7723), .D (
        nx4691), .CLK (CLK)) ;
    oai21 ix4702 (.Y (nx4701), .A0 (nx7729), .A1 (nx8050), .B0 (nx7731)) ;
    dff L0_0_L1_4_Fij_reg_Dout_5 (.Q (FilterDout_0__4__5), .QB (nx7729), .D (
        nx4701), .CLK (CLK)) ;
    oai21 ix4712 (.Y (nx4711), .A0 (nx7735), .A1 (nx8050), .B0 (nx7737)) ;
    dff L0_0_L1_4_Fij_reg_Dout_6 (.Q (FilterDout_0__4__6), .QB (nx7735), .D (
        nx4711), .CLK (CLK)) ;
    oai21 ix4722 (.Y (nx4721), .A0 (nx7741), .A1 (nx8050), .B0 (nx7743)) ;
    dff L0_0_L1_4_Fij_reg_Dout_7 (.Q (FilterDout_0__4__7), .QB (nx7741), .D (
        nx4721), .CLK (CLK)) ;
    oai21 ix4972 (.Y (nx4971), .A0 (nx7747), .A1 (nx8050), .B0 (nx7749)) ;
    dff L0_0_L1_3_Fij_reg_Dout_0 (.Q (FilterDout_0__3__0), .QB (nx7747), .D (
        nx4971), .CLK (CLK)) ;
    oai21 ix4982 (.Y (nx4981), .A0 (nx7753), .A1 (nx8052), .B0 (nx7755)) ;
    dff L0_0_L1_3_Fij_reg_Dout_1 (.Q (FilterDout_0__3__1), .QB (nx7753), .D (
        nx4981), .CLK (CLK)) ;
    oai21 ix4992 (.Y (nx4991), .A0 (nx7759), .A1 (nx8052), .B0 (nx7761)) ;
    dff L0_0_L1_3_Fij_reg_Dout_2 (.Q (FilterDout_0__3__2), .QB (nx7759), .D (
        nx4991), .CLK (CLK)) ;
    oai21 ix5002 (.Y (nx5001), .A0 (nx7765), .A1 (nx8052), .B0 (nx7767)) ;
    dff L0_0_L1_3_Fij_reg_Dout_3 (.Q (FilterDout_0__3__3), .QB (nx7765), .D (
        nx5001), .CLK (CLK)) ;
    oai21 ix5012 (.Y (nx5011), .A0 (nx7771), .A1 (nx8054), .B0 (nx7773)) ;
    dff L0_0_L1_3_Fij_reg_Dout_4 (.Q (FilterDout_0__3__4), .QB (nx7771), .D (
        nx5011), .CLK (CLK)) ;
    oai21 ix5022 (.Y (nx5021), .A0 (nx7777), .A1 (nx8054), .B0 (nx7779)) ;
    dff L0_0_L1_3_Fij_reg_Dout_5 (.Q (FilterDout_0__3__5), .QB (nx7777), .D (
        nx5021), .CLK (CLK)) ;
    oai21 ix5032 (.Y (nx5031), .A0 (nx7783), .A1 (nx8054), .B0 (nx7785)) ;
    dff L0_0_L1_3_Fij_reg_Dout_6 (.Q (FilterDout_0__3__6), .QB (nx7783), .D (
        nx5031), .CLK (CLK)) ;
    oai21 ix5042 (.Y (nx5041), .A0 (nx7789), .A1 (nx8054), .B0 (nx7791)) ;
    dff L0_0_L1_3_Fij_reg_Dout_7 (.Q (FilterDout_0__3__7), .QB (nx7789), .D (
        nx5041), .CLK (CLK)) ;
    oai21 ix5292 (.Y (nx5291), .A0 (nx7795), .A1 (nx8056), .B0 (nx7797)) ;
    dff L0_0_L1_2_Fij_reg_Dout_0 (.Q (FilterDout_0__2__0), .QB (nx7795), .D (
        nx5291), .CLK (CLK)) ;
    oai21 ix5302 (.Y (nx5301), .A0 (nx7801), .A1 (nx8056), .B0 (nx7803)) ;
    dff L0_0_L1_2_Fij_reg_Dout_1 (.Q (FilterDout_0__2__1), .QB (nx7801), .D (
        nx5301), .CLK (CLK)) ;
    oai21 ix5312 (.Y (nx5311), .A0 (nx7807), .A1 (nx8056), .B0 (nx7809)) ;
    dff L0_0_L1_2_Fij_reg_Dout_2 (.Q (FilterDout_0__2__2), .QB (nx7807), .D (
        nx5311), .CLK (CLK)) ;
    oai21 ix5322 (.Y (nx5321), .A0 (nx7813), .A1 (nx8058), .B0 (nx7815)) ;
    dff L0_0_L1_2_Fij_reg_Dout_3 (.Q (FilterDout_0__2__3), .QB (nx7813), .D (
        nx5321), .CLK (CLK)) ;
    oai21 ix5332 (.Y (nx5331), .A0 (nx7819), .A1 (nx8058), .B0 (nx7821)) ;
    dff L0_0_L1_2_Fij_reg_Dout_4 (.Q (FilterDout_0__2__4), .QB (nx7819), .D (
        nx5331), .CLK (CLK)) ;
    oai21 ix5342 (.Y (nx5341), .A0 (nx7825), .A1 (nx8058), .B0 (nx7827)) ;
    dff L0_0_L1_2_Fij_reg_Dout_5 (.Q (FilterDout_0__2__5), .QB (nx7825), .D (
        nx5341), .CLK (CLK)) ;
    oai21 ix5352 (.Y (nx5351), .A0 (nx7831), .A1 (nx8058), .B0 (nx7833)) ;
    dff L0_0_L1_2_Fij_reg_Dout_6 (.Q (FilterDout_0__2__6), .QB (nx7831), .D (
        nx5351), .CLK (CLK)) ;
    oai21 ix5362 (.Y (nx5361), .A0 (nx7837), .A1 (nx8060), .B0 (nx7839)) ;
    dff L0_0_L1_2_Fij_reg_Dout_7 (.Q (FilterDout_0__2__7), .QB (nx7837), .D (
        nx5361), .CLK (CLK)) ;
    oai21 ix5612 (.Y (nx5611), .A0 (nx7843), .A1 (nx8060), .B0 (nx7845)) ;
    dff L0_0_L1_1_Fij_reg_Dout_0 (.Q (FilterDout_0__1__0), .QB (nx7843), .D (
        nx5611), .CLK (CLK)) ;
    oai21 ix5622 (.Y (nx5621), .A0 (nx7849), .A1 (nx8060), .B0 (nx7851)) ;
    dff L0_0_L1_1_Fij_reg_Dout_1 (.Q (FilterDout_0__1__1), .QB (nx7849), .D (
        nx5621), .CLK (CLK)) ;
    oai21 ix5632 (.Y (nx5631), .A0 (nx7855), .A1 (nx8062), .B0 (nx7857)) ;
    dff L0_0_L1_1_Fij_reg_Dout_2 (.Q (FilterDout_0__1__2), .QB (nx7855), .D (
        nx5631), .CLK (CLK)) ;
    oai21 ix5642 (.Y (nx5641), .A0 (nx7861), .A1 (nx8062), .B0 (nx7863)) ;
    dff L0_0_L1_1_Fij_reg_Dout_3 (.Q (FilterDout_0__1__3), .QB (nx7861), .D (
        nx5641), .CLK (CLK)) ;
    oai21 ix5652 (.Y (nx5651), .A0 (nx7867), .A1 (nx8062), .B0 (nx7869)) ;
    dff L0_0_L1_1_Fij_reg_Dout_4 (.Q (FilterDout_0__1__4), .QB (nx7867), .D (
        nx5651), .CLK (CLK)) ;
    oai21 ix5662 (.Y (nx5661), .A0 (nx7873), .A1 (nx8062), .B0 (nx7875)) ;
    dff L0_0_L1_1_Fij_reg_Dout_5 (.Q (FilterDout_0__1__5), .QB (nx7873), .D (
        nx5661), .CLK (CLK)) ;
    oai21 ix5672 (.Y (nx5671), .A0 (nx7879), .A1 (nx8064), .B0 (nx7881)) ;
    dff L0_0_L1_1_Fij_reg_Dout_6 (.Q (FilterDout_0__1__6), .QB (nx7879), .D (
        nx5671), .CLK (CLK)) ;
    oai21 ix5682 (.Y (nx5681), .A0 (nx7885), .A1 (nx8064), .B0 (nx7887)) ;
    dff L0_0_L1_1_Fij_reg_Dout_7 (.Q (FilterDout_0__1__7), .QB (nx7885), .D (
        nx5681), .CLK (CLK)) ;
    oai21 ix5932 (.Y (nx5931), .A0 (nx7891), .A1 (nx8064), .B0 (nx7893)) ;
    dff L0_0_L1_0_Fij_reg_Dout_0 (.Q (FilterDout_0__0__0), .QB (nx7891), .D (
        nx5931), .CLK (CLK)) ;
    oai21 ix5942 (.Y (nx5941), .A0 (nx7897), .A1 (nx8066), .B0 (nx7899)) ;
    dff L0_0_L1_0_Fij_reg_Dout_1 (.Q (FilterDout_0__0__1), .QB (nx7897), .D (
        nx5941), .CLK (CLK)) ;
    oai21 ix5952 (.Y (nx5951), .A0 (nx7903), .A1 (nx8066), .B0 (nx7905)) ;
    dff L0_0_L1_0_Fij_reg_Dout_2 (.Q (FilterDout_0__0__2), .QB (nx7903), .D (
        nx5951), .CLK (CLK)) ;
    oai21 ix5962 (.Y (nx5961), .A0 (nx7909), .A1 (nx8066), .B0 (nx7911)) ;
    dff L0_0_L1_0_Fij_reg_Dout_3 (.Q (FilterDout_0__0__3), .QB (nx7909), .D (
        nx5961), .CLK (CLK)) ;
    oai21 ix5972 (.Y (nx5971), .A0 (nx7915), .A1 (nx8066), .B0 (nx7917)) ;
    dff L0_0_L1_0_Fij_reg_Dout_4 (.Q (FilterDout_0__0__4), .QB (nx7915), .D (
        nx5971), .CLK (CLK)) ;
    oai21 ix5982 (.Y (nx5981), .A0 (nx7921), .A1 (nx8068), .B0 (nx7923)) ;
    dff L0_0_L1_0_Fij_reg_Dout_5 (.Q (FilterDout_0__0__5), .QB (nx7921), .D (
        nx5981), .CLK (CLK)) ;
    oai21 ix5992 (.Y (nx5991), .A0 (nx7927), .A1 (nx8068), .B0 (nx7929)) ;
    dff L0_0_L1_0_Fij_reg_Dout_6 (.Q (FilterDout_0__0__6), .QB (nx7927), .D (
        nx5991), .CLK (CLK)) ;
    oai21 ix6002 (.Y (nx6001), .A0 (nx7933), .A1 (nx8068), .B0 (nx7935)) ;
    dff L0_0_L1_0_Fij_reg_Dout_7 (.Q (FilterDout_0__0__7), .QB (nx7933), .D (
        nx6001), .CLK (CLK)) ;
    inv02 ix169 (.Y (nx168), .A (nx6998)) ;
    inv02 ix85 (.Y (nx84), .A (nx6042)) ;
    inv02 ix7941 (.Y (nx7942), .A (nx8182)) ;
    inv02 ix7943 (.Y (nx7944), .A (nx8182)) ;
    inv02 ix7945 (.Y (nx7946), .A (nx8182)) ;
    inv02 ix7947 (.Y (nx7948), .A (nx8182)) ;
    inv02 ix7949 (.Y (nx7950), .A (nx8182)) ;
    inv02 ix7951 (.Y (nx7952), .A (nx8278)) ;
    inv02 ix7953 (.Y (nx7954), .A (nx8278)) ;
    inv02 ix7955 (.Y (nx7956), .A (nx8278)) ;
    inv02 ix7957 (.Y (nx7958), .A (nx8278)) ;
    inv02 ix7959 (.Y (nx7960), .A (nx8278)) ;
    inv02 ix7961 (.Y (nx7962), .A (nx8278)) ;
    inv02 ix7963 (.Y (nx7964), .A (nx8278)) ;
    inv02 ix7965 (.Y (nx7966), .A (nx8286)) ;
    inv02 ix7967 (.Y (nx7968), .A (nx8286)) ;
    inv02 ix7969 (.Y (nx7970), .A (nx8286)) ;
    inv02 ix7971 (.Y (nx7972), .A (nx8286)) ;
    inv02 ix7973 (.Y (nx7974), .A (nx8286)) ;
    inv02 ix7975 (.Y (nx7976), .A (nx8286)) ;
    inv02 ix7977 (.Y (nx7978), .A (nx8286)) ;
    inv02 ix7979 (.Y (nx7980), .A (nx8288)) ;
    inv02 ix7981 (.Y (nx7982), .A (nx8288)) ;
    inv02 ix7983 (.Y (nx7984), .A (nx8288)) ;
    inv02 ix7985 (.Y (nx7986), .A (nx8288)) ;
    inv02 ix7987 (.Y (nx7988), .A (nx8288)) ;
    inv02 ix7989 (.Y (nx7990), .A (nx8288)) ;
    inv02 ix7991 (.Y (nx7992), .A (nx8288)) ;
    inv02 ix7993 (.Y (nx7994), .A (nx8294)) ;
    inv02 ix7995 (.Y (nx7996), .A (nx8294)) ;
    inv02 ix7997 (.Y (nx7998), .A (nx8294)) ;
    inv02 ix7999 (.Y (nx8000), .A (nx8294)) ;
    inv02 ix8001 (.Y (nx8002), .A (nx8294)) ;
    inv02 ix8003 (.Y (nx8004), .A (nx8294)) ;
    inv02 ix8005 (.Y (nx8006), .A (nx8220)) ;
    inv02 ix8007 (.Y (nx8008), .A (nx8220)) ;
    inv02 ix8009 (.Y (nx8010), .A (nx8220)) ;
    inv02 ix8011 (.Y (nx8012), .A (nx8220)) ;
    inv02 ix8013 (.Y (nx8014), .A (nx8220)) ;
    inv02 ix8015 (.Y (nx8016), .A (nx8300)) ;
    inv02 ix8017 (.Y (nx8018), .A (nx8300)) ;
    inv02 ix8019 (.Y (nx8020), .A (nx8300)) ;
    inv02 ix8021 (.Y (nx8022), .A (nx8300)) ;
    inv02 ix8023 (.Y (nx8024), .A (nx8300)) ;
    inv02 ix8025 (.Y (nx8026), .A (nx8300)) ;
    inv02 ix8027 (.Y (nx8028), .A (nx8300)) ;
    inv02 ix8029 (.Y (nx8030), .A (nx8308)) ;
    inv02 ix8031 (.Y (nx8032), .A (nx8308)) ;
    inv02 ix8033 (.Y (nx8034), .A (nx8308)) ;
    inv02 ix8035 (.Y (nx8036), .A (nx8308)) ;
    inv02 ix8037 (.Y (nx8038), .A (nx8308)) ;
    inv02 ix8039 (.Y (nx8040), .A (nx8308)) ;
    inv02 ix8041 (.Y (nx8042), .A (nx8308)) ;
    inv02 ix8043 (.Y (nx8044), .A (nx8310)) ;
    inv02 ix8045 (.Y (nx8046), .A (nx8310)) ;
    inv02 ix8047 (.Y (nx8048), .A (nx8310)) ;
    inv02 ix8049 (.Y (nx8050), .A (nx8310)) ;
    inv02 ix8051 (.Y (nx8052), .A (nx8310)) ;
    inv02 ix8053 (.Y (nx8054), .A (nx8310)) ;
    inv02 ix8055 (.Y (nx8056), .A (nx8310)) ;
    inv02 ix8057 (.Y (nx8058), .A (nx8316)) ;
    inv02 ix8059 (.Y (nx8060), .A (nx8316)) ;
    inv02 ix8061 (.Y (nx8062), .A (nx8316)) ;
    inv02 ix8063 (.Y (nx8064), .A (nx8316)) ;
    inv02 ix8065 (.Y (nx8066), .A (nx8316)) ;
    inv02 ix8067 (.Y (nx8068), .A (nx8316)) ;
    inv02 ix8069 (.Y (nx8070), .A (RST)) ;
    inv02 ix8071 (.Y (nx8072), .A (RST)) ;
    inv02 ix8073 (.Y (nx8074), .A (RST)) ;
    inv02 ix8075 (.Y (nx8076), .A (RST)) ;
    inv02 ix8077 (.Y (nx8078), .A (RST)) ;
    inv02 ix8079 (.Y (nx8080), .A (RST)) ;
    inv02 ix8081 (.Y (nx8082), .A (RST)) ;
    inv02 ix8083 (.Y (nx8084), .A (RST)) ;
    inv02 ix8085 (.Y (nx8086), .A (RST)) ;
    inv02 ix8087 (.Y (nx8088), .A (RST)) ;
    inv02 ix8089 (.Y (nx8090), .A (RST)) ;
    inv02 ix8093 (.Y (nx8094), .A (RST)) ;
    inv02 ix8095 (.Y (nx8096), .A (RST)) ;
    inv02 ix8097 (.Y (nx8098), .A (RST)) ;
    inv02 ix8099 (.Y (nx8100), .A (RST)) ;
    inv02 ix8105 (.Y (nx8106), .A (RST)) ;
    inv02 ix8107 (.Y (nx8108), .A (RST)) ;
    inv02 ix8109 (.Y (nx8110), .A (RST)) ;
    inv02 ix8111 (.Y (nx8112), .A (RST)) ;
    inv02 ix8123 (.Y (nx8124), .A (RST)) ;
    inv02 ix8125 (.Y (nx8126), .A (RST)) ;
    inv02 ix8127 (.Y (nx8128), .A (RST)) ;
    inv02 ix8129 (.Y (nx8130), .A (RST)) ;
    inv02 ix8131 (.Y (nx8132), .A (RST)) ;
    inv02 ix8133 (.Y (nx8134), .A (RST)) ;
    inv02 ix8135 (.Y (nx8136), .A (RST)) ;
    inv02 ix8137 (.Y (nx8138), .A (RST)) ;
    inv02 ix8139 (.Y (nx8140), .A (RST)) ;
    inv02 ix8141 (.Y (nx8142), .A (RST)) ;
    inv02 ix8145 (.Y (nx8146), .A (RST)) ;
    inv02 ix8147 (.Y (nx8148), .A (RST)) ;
    inv02 ix8149 (.Y (nx8150), .A (RST)) ;
    inv02 ix8151 (.Y (nx8152), .A (RST)) ;
    inv02 ix8153 (.Y (nx8154), .A (RST)) ;
    inv02 ix8157 (.Y (nx8158), .A (RST)) ;
    inv02 ix8159 (.Y (nx8160), .A (RST)) ;
    inv02 ix8161 (.Y (nx8162), .A (RST)) ;
    inv02 ix8163 (.Y (nx8164), .A (RST)) ;
    inv02 ix8181 (.Y (nx8182), .A (nx8322)) ;
    inv02 ix8183 (.Y (nx8184), .A (nx8322)) ;
    inv02 ix8185 (.Y (nx8186), .A (nx8322)) ;
    inv02 ix8187 (.Y (nx8188), .A (nx8322)) ;
    inv02 ix8189 (.Y (nx8190), .A (nx8322)) ;
    inv02 ix8193 (.Y (nx8194), .A (nx8254)) ;
    inv02 ix8195 (.Y (nx8196), .A (nx8254)) ;
    inv02 ix8197 (.Y (nx8198), .A (nx8254)) ;
    inv02 ix8199 (.Y (nx8200), .A (nx8254)) ;
    inv02 ix8201 (.Y (nx8202), .A (nx8254)) ;
    inv02 ix8203 (.Y (nx8204), .A (nx8254)) ;
    inv02 ix8205 (.Y (nx8206), .A (nx8254)) ;
    inv02 ix8207 (.Y (nx8208), .A (nx8256)) ;
    inv02 ix8209 (.Y (nx8210), .A (nx8256)) ;
    inv02 ix8211 (.Y (nx8212), .A (nx8256)) ;
    inv02 ix8213 (.Y (nx8214), .A (nx8256)) ;
    inv02 ix8219 (.Y (nx8220), .A (nx8326)) ;
    inv02 ix8221 (.Y (nx8222), .A (nx8326)) ;
    inv02 ix8223 (.Y (nx8224), .A (nx8326)) ;
    inv02 ix8225 (.Y (nx8226), .A (nx8326)) ;
    inv02 ix8227 (.Y (nx8228), .A (nx8326)) ;
    inv02 ix8231 (.Y (nx8232), .A (nx8258)) ;
    inv02 ix8233 (.Y (nx8234), .A (nx8258)) ;
    inv02 ix8235 (.Y (nx8236), .A (nx8258)) ;
    inv02 ix8237 (.Y (nx8238), .A (nx8258)) ;
    inv02 ix8239 (.Y (nx8240), .A (nx8258)) ;
    inv02 ix8241 (.Y (nx8242), .A (nx8258)) ;
    inv02 ix8243 (.Y (nx8244), .A (nx8258)) ;
    inv02 ix8245 (.Y (nx8246), .A (nx8260)) ;
    inv02 ix8247 (.Y (nx8248), .A (nx8260)) ;
    inv02 ix8249 (.Y (nx8250), .A (nx8260)) ;
    inv02 ix8251 (.Y (nx8252), .A (nx8260)) ;
    inv02 ix8253 (.Y (nx8254), .A (nx6107)) ;
    inv02 ix8255 (.Y (nx8256), .A (nx6107)) ;
    inv02 ix8257 (.Y (nx8258), .A (nx7048)) ;
    inv02 ix8259 (.Y (nx8260), .A (nx7048)) ;
    mux21_ni ix2012 (.Y (nx2011), .A0 (WindowDout_4__4__0), .A1 (nx88), .S0 (
             nx8322)) ;
    mux21_ni ix2022 (.Y (nx2021), .A0 (WindowDout_4__4__1), .A1 (nx98), .S0 (
             nx8322)) ;
    mux21_ni ix2032 (.Y (nx2031), .A0 (WindowDout_4__4__2), .A1 (nx108), .S0 (
             nx8272)) ;
    mux21_ni ix2042 (.Y (nx2041), .A0 (WindowDout_4__4__3), .A1 (nx118), .S0 (
             nx8272)) ;
    mux21_ni ix2052 (.Y (nx2051), .A0 (WindowDout_4__4__4), .A1 (nx128), .S0 (
             nx8272)) ;
    mux21_ni ix2062 (.Y (nx2061), .A0 (WindowDout_4__4__5), .A1 (nx138), .S0 (
             nx8272)) ;
    mux21_ni ix2072 (.Y (nx2071), .A0 (WindowDout_4__4__6), .A1 (nx148), .S0 (
             nx8272)) ;
    mux21_ni ix2082 (.Y (nx2081), .A0 (WindowDout_4__4__7), .A1 (nx158), .S0 (
             nx8272)) ;
    mux21_ni ix2172 (.Y (nx2171), .A0 (WindowDout_4__3__0), .A1 (nx220), .S0 (
             nx8272)) ;
    mux21_ni ix2182 (.Y (nx2181), .A0 (WindowDout_4__3__1), .A1 (nx230), .S0 (
             nx84)) ;
    mux21_ni ix2192 (.Y (nx2191), .A0 (WindowDout_4__3__2), .A1 (nx240), .S0 (
             nx84)) ;
    mux21_ni ix2202 (.Y (nx2201), .A0 (WindowDout_4__3__3), .A1 (nx250), .S0 (
             nx84)) ;
    mux21_ni ix2212 (.Y (nx2211), .A0 (WindowDout_4__3__4), .A1 (nx260), .S0 (
             nx84)) ;
    mux21_ni ix2222 (.Y (nx2221), .A0 (WindowDout_4__3__5), .A1 (nx270), .S0 (
             nx84)) ;
    mux21_ni ix2232 (.Y (nx2231), .A0 (WindowDout_4__3__6), .A1 (nx280), .S0 (
             nx84)) ;
    mux21_ni ix2242 (.Y (nx2241), .A0 (WindowDout_4__3__7), .A1 (nx290), .S0 (
             nx84)) ;
    or03 ix6353 (.Y (nx6352), .A0 (RST), .A1 (nx6181), .A2 (nx8182)) ;
    or03 ix6359 (.Y (nx6358), .A0 (RST), .A1 (nx6188), .A2 (nx8280)) ;
    or03 ix6365 (.Y (nx6364), .A0 (RST), .A1 (nx6194), .A2 (nx8280)) ;
    or03 ix6371 (.Y (nx6370), .A0 (RST), .A1 (nx6200), .A2 (nx8280)) ;
    or03 ix6377 (.Y (nx6376), .A0 (RST), .A1 (nx6206), .A2 (nx8280)) ;
    or03 ix6383 (.Y (nx6382), .A0 (RST), .A1 (nx6212), .A2 (nx8280)) ;
    or03 ix6389 (.Y (nx6388), .A0 (RST), .A1 (nx6218), .A2 (nx8280)) ;
    or03 ix6395 (.Y (nx6394), .A0 (RST), .A1 (nx6224), .A2 (nx8280)) ;
    or03 ix6401 (.Y (nx6400), .A0 (RST), .A1 (nx6230), .A2 (nx8282)) ;
    or03 ix6407 (.Y (nx6406), .A0 (RST), .A1 (nx6236), .A2 (nx8282)) ;
    or03 ix6413 (.Y (nx6412), .A0 (RST), .A1 (nx6242), .A2 (nx8282)) ;
    or03 ix6419 (.Y (nx6418), .A0 (RST), .A1 (nx6248), .A2 (nx8282)) ;
    or03 ix6425 (.Y (nx6424), .A0 (RST), .A1 (nx6254), .A2 (nx8282)) ;
    or03 ix6431 (.Y (nx6430), .A0 (RST), .A1 (nx6260), .A2 (nx8282)) ;
    or03 ix6437 (.Y (nx6436), .A0 (RST), .A1 (nx6266), .A2 (nx8282)) ;
    or03 ix6443 (.Y (nx6442), .A0 (RST), .A1 (nx6272), .A2 (nx8284)) ;
    or03 ix6521 (.Y (nx6520), .A0 (RST), .A1 (nx6350), .A2 (nx8284)) ;
    or03 ix6527 (.Y (nx6526), .A0 (RST), .A1 (nx6356), .A2 (nx8284)) ;
    or03 ix6533 (.Y (nx6532), .A0 (RST), .A1 (nx6362), .A2 (nx8284)) ;
    or03 ix6539 (.Y (nx6538), .A0 (RST), .A1 (nx6368), .A2 (nx8284)) ;
    or03 ix6545 (.Y (nx6544), .A0 (RST), .A1 (nx6374), .A2 (nx8284)) ;
    or03 ix6551 (.Y (nx6550), .A0 (RST), .A1 (nx6380), .A2 (nx8284)) ;
    or03 ix6557 (.Y (nx6556), .A0 (RST), .A1 (nx6386), .A2 (nx8184)) ;
    or03 ix6563 (.Y (nx6562), .A0 (RST), .A1 (nx6392), .A2 (nx8184)) ;
    or03 ix6569 (.Y (nx6568), .A0 (RST), .A1 (nx6398), .A2 (nx8184)) ;
    or03 ix6575 (.Y (nx6574), .A0 (RST), .A1 (nx6404), .A2 (nx8184)) ;
    or03 ix6581 (.Y (nx6580), .A0 (RST), .A1 (nx6410), .A2 (nx8186)) ;
    or03 ix6587 (.Y (nx6586), .A0 (RST), .A1 (nx6416), .A2 (nx8186)) ;
    or03 ix6593 (.Y (nx6592), .A0 (RST), .A1 (nx6422), .A2 (nx8186)) ;
    or03 ix6599 (.Y (nx6598), .A0 (RST), .A1 (nx6428), .A2 (nx8186)) ;
    or03 ix6605 (.Y (nx6604), .A0 (RST), .A1 (nx6434), .A2 (nx8186)) ;
    or03 ix6611 (.Y (nx6610), .A0 (RST), .A1 (nx6440), .A2 (nx8186)) ;
    or03 ix6761 (.Y (nx6760), .A0 (RST), .A1 (nx6518), .A2 (nx8290)) ;
    or03 ix6767 (.Y (nx6766), .A0 (RST), .A1 (nx6524), .A2 (nx8290)) ;
    or03 ix6773 (.Y (nx6772), .A0 (RST), .A1 (nx6530), .A2 (nx8290)) ;
    or03 ix6779 (.Y (nx6778), .A0 (RST), .A1 (nx6536), .A2 (nx8290)) ;
    or03 ix6785 (.Y (nx6784), .A0 (RST), .A1 (nx6542), .A2 (nx8290)) ;
    or03 ix6791 (.Y (nx6790), .A0 (RST), .A1 (nx6548), .A2 (nx8290)) ;
    or03 ix6797 (.Y (nx6796), .A0 (RST), .A1 (nx6554), .A2 (nx8290)) ;
    or03 ix6803 (.Y (nx6802), .A0 (RST), .A1 (nx6560), .A2 (nx8292)) ;
    or03 ix6809 (.Y (nx6808), .A0 (RST), .A1 (nx6566), .A2 (nx8292)) ;
    or03 ix6815 (.Y (nx6814), .A0 (RST), .A1 (nx6572), .A2 (nx8292)) ;
    or03 ix6821 (.Y (nx6820), .A0 (RST), .A1 (nx6578), .A2 (nx8292)) ;
    or03 ix6827 (.Y (nx6826), .A0 (RST), .A1 (nx6584), .A2 (nx8292)) ;
    or03 ix6833 (.Y (nx6832), .A0 (RST), .A1 (nx6590), .A2 (nx8292)) ;
    or03 ix6839 (.Y (nx6838), .A0 (RST), .A1 (nx6596), .A2 (nx8292)) ;
    or03 ix6845 (.Y (nx6844), .A0 (RST), .A1 (nx6602), .A2 (nx8188)) ;
    or03 ix6851 (.Y (nx6850), .A0 (RST), .A1 (nx6608), .A2 (nx8188)) ;
    or03 ix6857 (.Y (nx6856), .A0 (RST), .A1 (nx6614), .A2 (nx8188)) ;
    or03 ix6863 (.Y (nx6862), .A0 (RST), .A1 (nx6620), .A2 (nx8188)) ;
    or03 ix6869 (.Y (nx6868), .A0 (RST), .A1 (nx6626), .A2 (nx8188)) ;
    or03 ix6875 (.Y (nx6874), .A0 (RST), .A1 (nx6632), .A2 (nx8294)) ;
    or03 ix6881 (.Y (nx6880), .A0 (RST), .A1 (nx6638), .A2 (nx8296)) ;
    or03 ix6887 (.Y (nx6886), .A0 (RST), .A1 (nx6644), .A2 (nx8296)) ;
    or03 ix6893 (.Y (nx6892), .A0 (RST), .A1 (nx6650), .A2 (nx8296)) ;
    or03 ix6899 (.Y (nx6898), .A0 (RST), .A1 (nx6656), .A2 (nx8296)) ;
    or03 ix6905 (.Y (nx6904), .A0 (RST), .A1 (nx6662), .A2 (nx8296)) ;
    or03 ix6911 (.Y (nx6910), .A0 (RST), .A1 (nx6668), .A2 (nx8296)) ;
    or03 ix6917 (.Y (nx6916), .A0 (RST), .A1 (nx6674), .A2 (nx8296)) ;
    or03 ix6923 (.Y (nx6922), .A0 (RST), .A1 (nx6680), .A2 (nx8298)) ;
    or03 ix6929 (.Y (nx6928), .A0 (RST), .A1 (nx6686), .A2 (nx8298)) ;
    or03 ix6935 (.Y (nx6934), .A0 (RST), .A1 (nx6692), .A2 (nx8298)) ;
    or03 ix6941 (.Y (nx6940), .A0 (RST), .A1 (nx6698), .A2 (nx8298)) ;
    or03 ix6947 (.Y (nx6946), .A0 (RST), .A1 (nx6704), .A2 (nx8298)) ;
    or03 ix6953 (.Y (nx6952), .A0 (RST), .A1 (nx6710), .A2 (nx8298)) ;
    or03 ix6959 (.Y (nx6958), .A0 (RST), .A1 (nx6716), .A2 (nx8298)) ;
    or03 ix6965 (.Y (nx6964), .A0 (RST), .A1 (nx6722), .A2 (nx8190)) ;
    or03 ix6971 (.Y (nx6970), .A0 (RST), .A1 (nx6728), .A2 (nx8190)) ;
    or03 ix6977 (.Y (nx6976), .A0 (RST), .A1 (nx6734), .A2 (nx8190)) ;
    or03 ix6983 (.Y (nx6982), .A0 (RST), .A1 (nx6740), .A2 (nx8190)) ;
    or03 ix6989 (.Y (nx6988), .A0 (RST), .A1 (nx6746), .A2 (nx8190)) ;
    or03 ix6995 (.Y (nx6994), .A0 (RST), .A1 (nx6752), .A2 (nx8190)) ;
    mux21_ni ix2092 (.Y (nx2091), .A0 (FilterDout_4__4__0), .A1 (nx88), .S0 (
             nx8326)) ;
    mux21_ni ix2102 (.Y (nx2101), .A0 (FilterDout_4__4__1), .A1 (nx98), .S0 (
             nx8326)) ;
    mux21_ni ix2112 (.Y (nx2111), .A0 (FilterDout_4__4__2), .A1 (nx108), .S0 (
             nx8276)) ;
    mux21_ni ix2122 (.Y (nx2121), .A0 (FilterDout_4__4__3), .A1 (nx118), .S0 (
             nx8276)) ;
    mux21_ni ix2132 (.Y (nx2131), .A0 (FilterDout_4__4__4), .A1 (nx128), .S0 (
             nx8276)) ;
    mux21_ni ix2142 (.Y (nx2141), .A0 (FilterDout_4__4__5), .A1 (nx138), .S0 (
             nx8276)) ;
    mux21_ni ix2152 (.Y (nx2151), .A0 (FilterDout_4__4__6), .A1 (nx148), .S0 (
             nx8276)) ;
    mux21_ni ix2162 (.Y (nx2161), .A0 (FilterDout_4__4__7), .A1 (nx158), .S0 (
             nx8276)) ;
    mux21_ni ix2252 (.Y (nx2251), .A0 (FilterDout_4__3__0), .A1 (nx220), .S0 (
             nx8276)) ;
    mux21_ni ix2262 (.Y (nx2261), .A0 (FilterDout_4__3__1), .A1 (nx230), .S0 (
             nx168)) ;
    mux21_ni ix2272 (.Y (nx2271), .A0 (FilterDout_4__3__2), .A1 (nx240), .S0 (
             nx168)) ;
    mux21_ni ix2282 (.Y (nx2281), .A0 (FilterDout_4__3__3), .A1 (nx250), .S0 (
             nx168)) ;
    mux21_ni ix2292 (.Y (nx2291), .A0 (FilterDout_4__3__4), .A1 (nx260), .S0 (
             nx168)) ;
    mux21_ni ix2302 (.Y (nx2301), .A0 (FilterDout_4__3__5), .A1 (nx270), .S0 (
             nx168)) ;
    mux21_ni ix2312 (.Y (nx2311), .A0 (FilterDout_4__3__6), .A1 (nx280), .S0 (
             nx168)) ;
    mux21_ni ix2322 (.Y (nx2321), .A0 (FilterDout_4__3__7), .A1 (nx290), .S0 (
             nx168)) ;
    or03 ix7294 (.Y (nx7293), .A0 (RST), .A1 (nx7122), .A2 (nx8220)) ;
    or03 ix7300 (.Y (nx7299), .A0 (RST), .A1 (nx7129), .A2 (nx8302)) ;
    or03 ix7306 (.Y (nx7305), .A0 (RST), .A1 (nx7135), .A2 (nx8302)) ;
    or03 ix7312 (.Y (nx7311), .A0 (RST), .A1 (nx7141), .A2 (nx8302)) ;
    or03 ix7318 (.Y (nx7317), .A0 (RST), .A1 (nx7147), .A2 (nx8302)) ;
    or03 ix7324 (.Y (nx7323), .A0 (RST), .A1 (nx7153), .A2 (nx8302)) ;
    or03 ix7330 (.Y (nx7329), .A0 (RST), .A1 (nx7159), .A2 (nx8302)) ;
    or03 ix7336 (.Y (nx7335), .A0 (RST), .A1 (nx7165), .A2 (nx8302)) ;
    or03 ix7342 (.Y (nx7341), .A0 (RST), .A1 (nx7171), .A2 (nx8304)) ;
    or03 ix7348 (.Y (nx7347), .A0 (RST), .A1 (nx7177), .A2 (nx8304)) ;
    or03 ix7354 (.Y (nx7353), .A0 (RST), .A1 (nx7183), .A2 (nx8304)) ;
    or03 ix7360 (.Y (nx7359), .A0 (RST), .A1 (nx7189), .A2 (nx8304)) ;
    or03 ix7366 (.Y (nx7365), .A0 (RST), .A1 (nx7195), .A2 (nx8304)) ;
    or03 ix7372 (.Y (nx7371), .A0 (RST), .A1 (nx7201), .A2 (nx8304)) ;
    or03 ix7378 (.Y (nx7377), .A0 (RST), .A1 (nx7207), .A2 (nx8304)) ;
    or03 ix7384 (.Y (nx7383), .A0 (RST), .A1 (nx7213), .A2 (nx8306)) ;
    or03 ix7462 (.Y (nx7461), .A0 (RST), .A1 (nx7291), .A2 (nx8306)) ;
    or03 ix7468 (.Y (nx7467), .A0 (RST), .A1 (nx7297), .A2 (nx8306)) ;
    or03 ix7474 (.Y (nx7473), .A0 (RST), .A1 (nx7303), .A2 (nx8306)) ;
    or03 ix7480 (.Y (nx7479), .A0 (RST), .A1 (nx7309), .A2 (nx8306)) ;
    or03 ix7486 (.Y (nx7485), .A0 (RST), .A1 (nx7315), .A2 (nx8306)) ;
    or03 ix7492 (.Y (nx7491), .A0 (RST), .A1 (nx7321), .A2 (nx8306)) ;
    or03 ix7498 (.Y (nx7497), .A0 (RST), .A1 (nx7327), .A2 (nx8222)) ;
    or03 ix7504 (.Y (nx7503), .A0 (RST), .A1 (nx7333), .A2 (nx8222)) ;
    or03 ix7510 (.Y (nx7509), .A0 (RST), .A1 (nx7339), .A2 (nx8222)) ;
    or03 ix7516 (.Y (nx7515), .A0 (RST), .A1 (nx7345), .A2 (nx8222)) ;
    or03 ix7522 (.Y (nx7521), .A0 (RST), .A1 (nx7351), .A2 (nx8224)) ;
    or03 ix7528 (.Y (nx7527), .A0 (RST), .A1 (nx7357), .A2 (nx8224)) ;
    or03 ix7534 (.Y (nx7533), .A0 (RST), .A1 (nx7363), .A2 (nx8224)) ;
    or03 ix7540 (.Y (nx7539), .A0 (RST), .A1 (nx7369), .A2 (nx8224)) ;
    or03 ix7546 (.Y (nx7545), .A0 (RST), .A1 (nx7375), .A2 (nx8224)) ;
    or03 ix7552 (.Y (nx7551), .A0 (RST), .A1 (nx7381), .A2 (nx8224)) ;
    or03 ix7702 (.Y (nx7701), .A0 (RST), .A1 (nx7459), .A2 (nx8312)) ;
    or03 ix7708 (.Y (nx7707), .A0 (RST), .A1 (nx7465), .A2 (nx8312)) ;
    or03 ix7714 (.Y (nx7713), .A0 (RST), .A1 (nx7471), .A2 (nx8312)) ;
    or03 ix7720 (.Y (nx7719), .A0 (RST), .A1 (nx7477), .A2 (nx8312)) ;
    or03 ix7726 (.Y (nx7725), .A0 (RST), .A1 (nx7483), .A2 (nx8312)) ;
    or03 ix7732 (.Y (nx7731), .A0 (RST), .A1 (nx7489), .A2 (nx8312)) ;
    or03 ix7738 (.Y (nx7737), .A0 (RST), .A1 (nx7495), .A2 (nx8312)) ;
    or03 ix7744 (.Y (nx7743), .A0 (RST), .A1 (nx7501), .A2 (nx8314)) ;
    or03 ix7750 (.Y (nx7749), .A0 (RST), .A1 (nx7507), .A2 (nx8314)) ;
    or03 ix7756 (.Y (nx7755), .A0 (RST), .A1 (nx7513), .A2 (nx8314)) ;
    or03 ix7762 (.Y (nx7761), .A0 (RST), .A1 (nx7519), .A2 (nx8314)) ;
    or03 ix7768 (.Y (nx7767), .A0 (RST), .A1 (nx7525), .A2 (nx8314)) ;
    or03 ix7774 (.Y (nx7773), .A0 (RST), .A1 (nx7531), .A2 (nx8314)) ;
    or03 ix7780 (.Y (nx7779), .A0 (RST), .A1 (nx7537), .A2 (nx8314)) ;
    or03 ix7786 (.Y (nx7785), .A0 (RST), .A1 (nx7543), .A2 (nx8226)) ;
    or03 ix7792 (.Y (nx7791), .A0 (RST), .A1 (nx7549), .A2 (nx8226)) ;
    or03 ix7798 (.Y (nx7797), .A0 (RST), .A1 (nx7555), .A2 (nx8226)) ;
    or03 ix7804 (.Y (nx7803), .A0 (RST), .A1 (nx7561), .A2 (nx8226)) ;
    or03 ix7810 (.Y (nx7809), .A0 (RST), .A1 (nx7567), .A2 (nx8226)) ;
    or03 ix7816 (.Y (nx7815), .A0 (RST), .A1 (nx7573), .A2 (nx8316)) ;
    or03 ix7822 (.Y (nx7821), .A0 (RST), .A1 (nx7579), .A2 (nx8318)) ;
    or03 ix7828 (.Y (nx7827), .A0 (RST), .A1 (nx7585), .A2 (nx8318)) ;
    or03 ix7834 (.Y (nx7833), .A0 (RST), .A1 (nx7591), .A2 (nx8318)) ;
    or03 ix7840 (.Y (nx7839), .A0 (RST), .A1 (nx7597), .A2 (nx8318)) ;
    or03 ix7846 (.Y (nx7845), .A0 (RST), .A1 (nx7603), .A2 (nx8318)) ;
    or03 ix7852 (.Y (nx7851), .A0 (RST), .A1 (nx7609), .A2 (nx8318)) ;
    or03 ix7858 (.Y (nx7857), .A0 (RST), .A1 (nx7615), .A2 (nx8318)) ;
    or03 ix7864 (.Y (nx7863), .A0 (RST), .A1 (nx7621), .A2 (nx8320)) ;
    or03 ix7870 (.Y (nx7869), .A0 (RST), .A1 (nx7627), .A2 (nx8320)) ;
    or03 ix7876 (.Y (nx7875), .A0 (RST), .A1 (nx7633), .A2 (nx8320)) ;
    or03 ix7882 (.Y (nx7881), .A0 (RST), .A1 (nx7639), .A2 (nx8320)) ;
    or03 ix7888 (.Y (nx7887), .A0 (RST), .A1 (nx7645), .A2 (nx8320)) ;
    or03 ix7894 (.Y (nx7893), .A0 (RST), .A1 (nx7651), .A2 (nx8320)) ;
    or03 ix7900 (.Y (nx7899), .A0 (RST), .A1 (nx7657), .A2 (nx8320)) ;
    or03 ix7906 (.Y (nx7905), .A0 (RST), .A1 (nx7663), .A2 (nx8228)) ;
    or03 ix7912 (.Y (nx7911), .A0 (RST), .A1 (nx7669), .A2 (nx8228)) ;
    or03 ix7918 (.Y (nx7917), .A0 (RST), .A1 (nx7675), .A2 (nx8228)) ;
    or03 ix7924 (.Y (nx7923), .A0 (RST), .A1 (nx7681), .A2 (nx8228)) ;
    or03 ix7930 (.Y (nx7929), .A0 (RST), .A1 (nx7687), .A2 (nx8228)) ;
    or03 ix7936 (.Y (nx7935), .A0 (RST), .A1 (nx7693), .A2 (nx8228)) ;
    inv02 ix8269 (.Y (nx8270), .A (nx8334)) ;
    inv02 ix8271 (.Y (nx8272), .A (nx8334)) ;
    inv02 ix8273 (.Y (nx8274), .A (nx8336)) ;
    inv02 ix8275 (.Y (nx8276), .A (nx8336)) ;
    inv02 ix8277 (.Y (nx8278), .A (nx8324)) ;
    inv02 ix8279 (.Y (nx8280), .A (nx8324)) ;
    inv02 ix8281 (.Y (nx8282), .A (nx8324)) ;
    inv02 ix8283 (.Y (nx8284), .A (nx8324)) ;
    inv02 ix8285 (.Y (nx8286), .A (nx8324)) ;
    inv02 ix8287 (.Y (nx8288), .A (nx8324)) ;
    inv02 ix8289 (.Y (nx8290), .A (nx8324)) ;
    inv02 ix8291 (.Y (nx8292), .A (nx8270)) ;
    inv02 ix8293 (.Y (nx8294), .A (nx8270)) ;
    inv02 ix8295 (.Y (nx8296), .A (nx8270)) ;
    inv02 ix8297 (.Y (nx8298), .A (nx8270)) ;
    inv02 ix8299 (.Y (nx8300), .A (nx8328)) ;
    inv02 ix8301 (.Y (nx8302), .A (nx8328)) ;
    inv02 ix8303 (.Y (nx8304), .A (nx8328)) ;
    inv02 ix8305 (.Y (nx8306), .A (nx8328)) ;
    inv02 ix8307 (.Y (nx8308), .A (nx8328)) ;
    inv02 ix8309 (.Y (nx8310), .A (nx8328)) ;
    inv02 ix8311 (.Y (nx8312), .A (nx8328)) ;
    inv02 ix8313 (.Y (nx8314), .A (nx8274)) ;
    inv02 ix8315 (.Y (nx8316), .A (nx8274)) ;
    inv02 ix8317 (.Y (nx8318), .A (nx8274)) ;
    inv02 ix8319 (.Y (nx8320), .A (nx8274)) ;
    inv02 ix8321 (.Y (nx8322), .A (nx8334)) ;
    inv02 ix8323 (.Y (nx8324), .A (nx8334)) ;
    inv02 ix8325 (.Y (nx8326), .A (nx8336)) ;
    inv02 ix8327 (.Y (nx8328), .A (nx8336)) ;
    inv01 ix8333 (.Y (nx8334), .A (nx84)) ;
    inv01 ix8335 (.Y (nx8336), .A (nx168)) ;
endmodule

