//
// Verilog description for cell calculator, 
// Sat May 12 15:09:22 2018
//
// LeonardoSpectrum Level 3, 2017a.2 
//


module calculator ( CLK, RST, Start, FilterSize, Instr, FilterDin_0__0__7, 
                    FilterDin_0__0__6, FilterDin_0__0__5, FilterDin_0__0__4, 
                    FilterDin_0__0__3, FilterDin_0__0__2, FilterDin_0__0__1, 
                    FilterDin_0__0__0, FilterDin_0__1__7, FilterDin_0__1__6, 
                    FilterDin_0__1__5, FilterDin_0__1__4, FilterDin_0__1__3, 
                    FilterDin_0__1__2, FilterDin_0__1__1, FilterDin_0__1__0, 
                    FilterDin_0__2__7, FilterDin_0__2__6, FilterDin_0__2__5, 
                    FilterDin_0__2__4, FilterDin_0__2__3, FilterDin_0__2__2, 
                    FilterDin_0__2__1, FilterDin_0__2__0, FilterDin_0__3__7, 
                    FilterDin_0__3__6, FilterDin_0__3__5, FilterDin_0__3__4, 
                    FilterDin_0__3__3, FilterDin_0__3__2, FilterDin_0__3__1, 
                    FilterDin_0__3__0, FilterDin_0__4__7, FilterDin_0__4__6, 
                    FilterDin_0__4__5, FilterDin_0__4__4, FilterDin_0__4__3, 
                    FilterDin_0__4__2, FilterDin_0__4__1, FilterDin_0__4__0, 
                    FilterDin_1__0__7, FilterDin_1__0__6, FilterDin_1__0__5, 
                    FilterDin_1__0__4, FilterDin_1__0__3, FilterDin_1__0__2, 
                    FilterDin_1__0__1, FilterDin_1__0__0, FilterDin_1__1__7, 
                    FilterDin_1__1__6, FilterDin_1__1__5, FilterDin_1__1__4, 
                    FilterDin_1__1__3, FilterDin_1__1__2, FilterDin_1__1__1, 
                    FilterDin_1__1__0, FilterDin_1__2__7, FilterDin_1__2__6, 
                    FilterDin_1__2__5, FilterDin_1__2__4, FilterDin_1__2__3, 
                    FilterDin_1__2__2, FilterDin_1__2__1, FilterDin_1__2__0, 
                    FilterDin_1__3__7, FilterDin_1__3__6, FilterDin_1__3__5, 
                    FilterDin_1__3__4, FilterDin_1__3__3, FilterDin_1__3__2, 
                    FilterDin_1__3__1, FilterDin_1__3__0, FilterDin_1__4__7, 
                    FilterDin_1__4__6, FilterDin_1__4__5, FilterDin_1__4__4, 
                    FilterDin_1__4__3, FilterDin_1__4__2, FilterDin_1__4__1, 
                    FilterDin_1__4__0, FilterDin_2__0__7, FilterDin_2__0__6, 
                    FilterDin_2__0__5, FilterDin_2__0__4, FilterDin_2__0__3, 
                    FilterDin_2__0__2, FilterDin_2__0__1, FilterDin_2__0__0, 
                    FilterDin_2__1__7, FilterDin_2__1__6, FilterDin_2__1__5, 
                    FilterDin_2__1__4, FilterDin_2__1__3, FilterDin_2__1__2, 
                    FilterDin_2__1__1, FilterDin_2__1__0, FilterDin_2__2__7, 
                    FilterDin_2__2__6, FilterDin_2__2__5, FilterDin_2__2__4, 
                    FilterDin_2__2__3, FilterDin_2__2__2, FilterDin_2__2__1, 
                    FilterDin_2__2__0, FilterDin_2__3__7, FilterDin_2__3__6, 
                    FilterDin_2__3__5, FilterDin_2__3__4, FilterDin_2__3__3, 
                    FilterDin_2__3__2, FilterDin_2__3__1, FilterDin_2__3__0, 
                    FilterDin_2__4__7, FilterDin_2__4__6, FilterDin_2__4__5, 
                    FilterDin_2__4__4, FilterDin_2__4__3, FilterDin_2__4__2, 
                    FilterDin_2__4__1, FilterDin_2__4__0, FilterDin_3__0__7, 
                    FilterDin_3__0__6, FilterDin_3__0__5, FilterDin_3__0__4, 
                    FilterDin_3__0__3, FilterDin_3__0__2, FilterDin_3__0__1, 
                    FilterDin_3__0__0, FilterDin_3__1__7, FilterDin_3__1__6, 
                    FilterDin_3__1__5, FilterDin_3__1__4, FilterDin_3__1__3, 
                    FilterDin_3__1__2, FilterDin_3__1__1, FilterDin_3__1__0, 
                    FilterDin_3__2__7, FilterDin_3__2__6, FilterDin_3__2__5, 
                    FilterDin_3__2__4, FilterDin_3__2__3, FilterDin_3__2__2, 
                    FilterDin_3__2__1, FilterDin_3__2__0, FilterDin_3__3__7, 
                    FilterDin_3__3__6, FilterDin_3__3__5, FilterDin_3__3__4, 
                    FilterDin_3__3__3, FilterDin_3__3__2, FilterDin_3__3__1, 
                    FilterDin_3__3__0, FilterDin_3__4__7, FilterDin_3__4__6, 
                    FilterDin_3__4__5, FilterDin_3__4__4, FilterDin_3__4__3, 
                    FilterDin_3__4__2, FilterDin_3__4__1, FilterDin_3__4__0, 
                    FilterDin_4__0__7, FilterDin_4__0__6, FilterDin_4__0__5, 
                    FilterDin_4__0__4, FilterDin_4__0__3, FilterDin_4__0__2, 
                    FilterDin_4__0__1, FilterDin_4__0__0, FilterDin_4__1__7, 
                    FilterDin_4__1__6, FilterDin_4__1__5, FilterDin_4__1__4, 
                    FilterDin_4__1__3, FilterDin_4__1__2, FilterDin_4__1__1, 
                    FilterDin_4__1__0, FilterDin_4__2__7, FilterDin_4__2__6, 
                    FilterDin_4__2__5, FilterDin_4__2__4, FilterDin_4__2__3, 
                    FilterDin_4__2__2, FilterDin_4__2__1, FilterDin_4__2__0, 
                    FilterDin_4__3__7, FilterDin_4__3__6, FilterDin_4__3__5, 
                    FilterDin_4__3__4, FilterDin_4__3__3, FilterDin_4__3__2, 
                    FilterDin_4__3__1, FilterDin_4__3__0, FilterDin_4__4__7, 
                    FilterDin_4__4__6, FilterDin_4__4__5, FilterDin_4__4__4, 
                    FilterDin_4__4__3, FilterDin_4__4__2, FilterDin_4__4__1, 
                    FilterDin_4__4__0, WindowDin_0__0__7, WindowDin_0__0__6, 
                    WindowDin_0__0__5, WindowDin_0__0__4, WindowDin_0__0__3, 
                    WindowDin_0__0__2, WindowDin_0__0__1, WindowDin_0__0__0, 
                    WindowDin_0__1__7, WindowDin_0__1__6, WindowDin_0__1__5, 
                    WindowDin_0__1__4, WindowDin_0__1__3, WindowDin_0__1__2, 
                    WindowDin_0__1__1, WindowDin_0__1__0, WindowDin_0__2__7, 
                    WindowDin_0__2__6, WindowDin_0__2__5, WindowDin_0__2__4, 
                    WindowDin_0__2__3, WindowDin_0__2__2, WindowDin_0__2__1, 
                    WindowDin_0__2__0, WindowDin_0__3__7, WindowDin_0__3__6, 
                    WindowDin_0__3__5, WindowDin_0__3__4, WindowDin_0__3__3, 
                    WindowDin_0__3__2, WindowDin_0__3__1, WindowDin_0__3__0, 
                    WindowDin_0__4__7, WindowDin_0__4__6, WindowDin_0__4__5, 
                    WindowDin_0__4__4, WindowDin_0__4__3, WindowDin_0__4__2, 
                    WindowDin_0__4__1, WindowDin_0__4__0, WindowDin_1__0__7, 
                    WindowDin_1__0__6, WindowDin_1__0__5, WindowDin_1__0__4, 
                    WindowDin_1__0__3, WindowDin_1__0__2, WindowDin_1__0__1, 
                    WindowDin_1__0__0, WindowDin_1__1__7, WindowDin_1__1__6, 
                    WindowDin_1__1__5, WindowDin_1__1__4, WindowDin_1__1__3, 
                    WindowDin_1__1__2, WindowDin_1__1__1, WindowDin_1__1__0, 
                    WindowDin_1__2__7, WindowDin_1__2__6, WindowDin_1__2__5, 
                    WindowDin_1__2__4, WindowDin_1__2__3, WindowDin_1__2__2, 
                    WindowDin_1__2__1, WindowDin_1__2__0, WindowDin_1__3__7, 
                    WindowDin_1__3__6, WindowDin_1__3__5, WindowDin_1__3__4, 
                    WindowDin_1__3__3, WindowDin_1__3__2, WindowDin_1__3__1, 
                    WindowDin_1__3__0, WindowDin_1__4__7, WindowDin_1__4__6, 
                    WindowDin_1__4__5, WindowDin_1__4__4, WindowDin_1__4__3, 
                    WindowDin_1__4__2, WindowDin_1__4__1, WindowDin_1__4__0, 
                    WindowDin_2__0__7, WindowDin_2__0__6, WindowDin_2__0__5, 
                    WindowDin_2__0__4, WindowDin_2__0__3, WindowDin_2__0__2, 
                    WindowDin_2__0__1, WindowDin_2__0__0, WindowDin_2__1__7, 
                    WindowDin_2__1__6, WindowDin_2__1__5, WindowDin_2__1__4, 
                    WindowDin_2__1__3, WindowDin_2__1__2, WindowDin_2__1__1, 
                    WindowDin_2__1__0, WindowDin_2__2__7, WindowDin_2__2__6, 
                    WindowDin_2__2__5, WindowDin_2__2__4, WindowDin_2__2__3, 
                    WindowDin_2__2__2, WindowDin_2__2__1, WindowDin_2__2__0, 
                    WindowDin_2__3__7, WindowDin_2__3__6, WindowDin_2__3__5, 
                    WindowDin_2__3__4, WindowDin_2__3__3, WindowDin_2__3__2, 
                    WindowDin_2__3__1, WindowDin_2__3__0, WindowDin_2__4__7, 
                    WindowDin_2__4__6, WindowDin_2__4__5, WindowDin_2__4__4, 
                    WindowDin_2__4__3, WindowDin_2__4__2, WindowDin_2__4__1, 
                    WindowDin_2__4__0, WindowDin_3__0__7, WindowDin_3__0__6, 
                    WindowDin_3__0__5, WindowDin_3__0__4, WindowDin_3__0__3, 
                    WindowDin_3__0__2, WindowDin_3__0__1, WindowDin_3__0__0, 
                    WindowDin_3__1__7, WindowDin_3__1__6, WindowDin_3__1__5, 
                    WindowDin_3__1__4, WindowDin_3__1__3, WindowDin_3__1__2, 
                    WindowDin_3__1__1, WindowDin_3__1__0, WindowDin_3__2__7, 
                    WindowDin_3__2__6, WindowDin_3__2__5, WindowDin_3__2__4, 
                    WindowDin_3__2__3, WindowDin_3__2__2, WindowDin_3__2__1, 
                    WindowDin_3__2__0, WindowDin_3__3__7, WindowDin_3__3__6, 
                    WindowDin_3__3__5, WindowDin_3__3__4, WindowDin_3__3__3, 
                    WindowDin_3__3__2, WindowDin_3__3__1, WindowDin_3__3__0, 
                    WindowDin_3__4__7, WindowDin_3__4__6, WindowDin_3__4__5, 
                    WindowDin_3__4__4, WindowDin_3__4__3, WindowDin_3__4__2, 
                    WindowDin_3__4__1, WindowDin_3__4__0, WindowDin_4__0__7, 
                    WindowDin_4__0__6, WindowDin_4__0__5, WindowDin_4__0__4, 
                    WindowDin_4__0__3, WindowDin_4__0__2, WindowDin_4__0__1, 
                    WindowDin_4__0__0, WindowDin_4__1__7, WindowDin_4__1__6, 
                    WindowDin_4__1__5, WindowDin_4__1__4, WindowDin_4__1__3, 
                    WindowDin_4__1__2, WindowDin_4__1__1, WindowDin_4__1__0, 
                    WindowDin_4__2__7, WindowDin_4__2__6, WindowDin_4__2__5, 
                    WindowDin_4__2__4, WindowDin_4__2__3, WindowDin_4__2__2, 
                    WindowDin_4__2__1, WindowDin_4__2__0, WindowDin_4__3__7, 
                    WindowDin_4__3__6, WindowDin_4__3__5, WindowDin_4__3__4, 
                    WindowDin_4__3__3, WindowDin_4__3__2, WindowDin_4__3__1, 
                    WindowDin_4__3__0, WindowDin_4__4__7, WindowDin_4__4__6, 
                    WindowDin_4__4__5, WindowDin_4__4__4, WindowDin_4__4__3, 
                    WindowDin_4__4__2, WindowDin_4__4__1, WindowDin_4__4__0, 
                    Done, Result ) ;

    input CLK ;
    input RST ;
    input Start ;
    input FilterSize ;
    input Instr ;
    input FilterDin_0__0__7 ;
    input FilterDin_0__0__6 ;
    input FilterDin_0__0__5 ;
    input FilterDin_0__0__4 ;
    input FilterDin_0__0__3 ;
    input FilterDin_0__0__2 ;
    input FilterDin_0__0__1 ;
    input FilterDin_0__0__0 ;
    input FilterDin_0__1__7 ;
    input FilterDin_0__1__6 ;
    input FilterDin_0__1__5 ;
    input FilterDin_0__1__4 ;
    input FilterDin_0__1__3 ;
    input FilterDin_0__1__2 ;
    input FilterDin_0__1__1 ;
    input FilterDin_0__1__0 ;
    input FilterDin_0__2__7 ;
    input FilterDin_0__2__6 ;
    input FilterDin_0__2__5 ;
    input FilterDin_0__2__4 ;
    input FilterDin_0__2__3 ;
    input FilterDin_0__2__2 ;
    input FilterDin_0__2__1 ;
    input FilterDin_0__2__0 ;
    input FilterDin_0__3__7 ;
    input FilterDin_0__3__6 ;
    input FilterDin_0__3__5 ;
    input FilterDin_0__3__4 ;
    input FilterDin_0__3__3 ;
    input FilterDin_0__3__2 ;
    input FilterDin_0__3__1 ;
    input FilterDin_0__3__0 ;
    input FilterDin_0__4__7 ;
    input FilterDin_0__4__6 ;
    input FilterDin_0__4__5 ;
    input FilterDin_0__4__4 ;
    input FilterDin_0__4__3 ;
    input FilterDin_0__4__2 ;
    input FilterDin_0__4__1 ;
    input FilterDin_0__4__0 ;
    input FilterDin_1__0__7 ;
    input FilterDin_1__0__6 ;
    input FilterDin_1__0__5 ;
    input FilterDin_1__0__4 ;
    input FilterDin_1__0__3 ;
    input FilterDin_1__0__2 ;
    input FilterDin_1__0__1 ;
    input FilterDin_1__0__0 ;
    input FilterDin_1__1__7 ;
    input FilterDin_1__1__6 ;
    input FilterDin_1__1__5 ;
    input FilterDin_1__1__4 ;
    input FilterDin_1__1__3 ;
    input FilterDin_1__1__2 ;
    input FilterDin_1__1__1 ;
    input FilterDin_1__1__0 ;
    input FilterDin_1__2__7 ;
    input FilterDin_1__2__6 ;
    input FilterDin_1__2__5 ;
    input FilterDin_1__2__4 ;
    input FilterDin_1__2__3 ;
    input FilterDin_1__2__2 ;
    input FilterDin_1__2__1 ;
    input FilterDin_1__2__0 ;
    input FilterDin_1__3__7 ;
    input FilterDin_1__3__6 ;
    input FilterDin_1__3__5 ;
    input FilterDin_1__3__4 ;
    input FilterDin_1__3__3 ;
    input FilterDin_1__3__2 ;
    input FilterDin_1__3__1 ;
    input FilterDin_1__3__0 ;
    input FilterDin_1__4__7 ;
    input FilterDin_1__4__6 ;
    input FilterDin_1__4__5 ;
    input FilterDin_1__4__4 ;
    input FilterDin_1__4__3 ;
    input FilterDin_1__4__2 ;
    input FilterDin_1__4__1 ;
    input FilterDin_1__4__0 ;
    input FilterDin_2__0__7 ;
    input FilterDin_2__0__6 ;
    input FilterDin_2__0__5 ;
    input FilterDin_2__0__4 ;
    input FilterDin_2__0__3 ;
    input FilterDin_2__0__2 ;
    input FilterDin_2__0__1 ;
    input FilterDin_2__0__0 ;
    input FilterDin_2__1__7 ;
    input FilterDin_2__1__6 ;
    input FilterDin_2__1__5 ;
    input FilterDin_2__1__4 ;
    input FilterDin_2__1__3 ;
    input FilterDin_2__1__2 ;
    input FilterDin_2__1__1 ;
    input FilterDin_2__1__0 ;
    input FilterDin_2__2__7 ;
    input FilterDin_2__2__6 ;
    input FilterDin_2__2__5 ;
    input FilterDin_2__2__4 ;
    input FilterDin_2__2__3 ;
    input FilterDin_2__2__2 ;
    input FilterDin_2__2__1 ;
    input FilterDin_2__2__0 ;
    input FilterDin_2__3__7 ;
    input FilterDin_2__3__6 ;
    input FilterDin_2__3__5 ;
    input FilterDin_2__3__4 ;
    input FilterDin_2__3__3 ;
    input FilterDin_2__3__2 ;
    input FilterDin_2__3__1 ;
    input FilterDin_2__3__0 ;
    input FilterDin_2__4__7 ;
    input FilterDin_2__4__6 ;
    input FilterDin_2__4__5 ;
    input FilterDin_2__4__4 ;
    input FilterDin_2__4__3 ;
    input FilterDin_2__4__2 ;
    input FilterDin_2__4__1 ;
    input FilterDin_2__4__0 ;
    input FilterDin_3__0__7 ;
    input FilterDin_3__0__6 ;
    input FilterDin_3__0__5 ;
    input FilterDin_3__0__4 ;
    input FilterDin_3__0__3 ;
    input FilterDin_3__0__2 ;
    input FilterDin_3__0__1 ;
    input FilterDin_3__0__0 ;
    input FilterDin_3__1__7 ;
    input FilterDin_3__1__6 ;
    input FilterDin_3__1__5 ;
    input FilterDin_3__1__4 ;
    input FilterDin_3__1__3 ;
    input FilterDin_3__1__2 ;
    input FilterDin_3__1__1 ;
    input FilterDin_3__1__0 ;
    input FilterDin_3__2__7 ;
    input FilterDin_3__2__6 ;
    input FilterDin_3__2__5 ;
    input FilterDin_3__2__4 ;
    input FilterDin_3__2__3 ;
    input FilterDin_3__2__2 ;
    input FilterDin_3__2__1 ;
    input FilterDin_3__2__0 ;
    input FilterDin_3__3__7 ;
    input FilterDin_3__3__6 ;
    input FilterDin_3__3__5 ;
    input FilterDin_3__3__4 ;
    input FilterDin_3__3__3 ;
    input FilterDin_3__3__2 ;
    input FilterDin_3__3__1 ;
    input FilterDin_3__3__0 ;
    input FilterDin_3__4__7 ;
    input FilterDin_3__4__6 ;
    input FilterDin_3__4__5 ;
    input FilterDin_3__4__4 ;
    input FilterDin_3__4__3 ;
    input FilterDin_3__4__2 ;
    input FilterDin_3__4__1 ;
    input FilterDin_3__4__0 ;
    input FilterDin_4__0__7 ;
    input FilterDin_4__0__6 ;
    input FilterDin_4__0__5 ;
    input FilterDin_4__0__4 ;
    input FilterDin_4__0__3 ;
    input FilterDin_4__0__2 ;
    input FilterDin_4__0__1 ;
    input FilterDin_4__0__0 ;
    input FilterDin_4__1__7 ;
    input FilterDin_4__1__6 ;
    input FilterDin_4__1__5 ;
    input FilterDin_4__1__4 ;
    input FilterDin_4__1__3 ;
    input FilterDin_4__1__2 ;
    input FilterDin_4__1__1 ;
    input FilterDin_4__1__0 ;
    input FilterDin_4__2__7 ;
    input FilterDin_4__2__6 ;
    input FilterDin_4__2__5 ;
    input FilterDin_4__2__4 ;
    input FilterDin_4__2__3 ;
    input FilterDin_4__2__2 ;
    input FilterDin_4__2__1 ;
    input FilterDin_4__2__0 ;
    input FilterDin_4__3__7 ;
    input FilterDin_4__3__6 ;
    input FilterDin_4__3__5 ;
    input FilterDin_4__3__4 ;
    input FilterDin_4__3__3 ;
    input FilterDin_4__3__2 ;
    input FilterDin_4__3__1 ;
    input FilterDin_4__3__0 ;
    input FilterDin_4__4__7 ;
    input FilterDin_4__4__6 ;
    input FilterDin_4__4__5 ;
    input FilterDin_4__4__4 ;
    input FilterDin_4__4__3 ;
    input FilterDin_4__4__2 ;
    input FilterDin_4__4__1 ;
    input FilterDin_4__4__0 ;
    input WindowDin_0__0__7 ;
    input WindowDin_0__0__6 ;
    input WindowDin_0__0__5 ;
    input WindowDin_0__0__4 ;
    input WindowDin_0__0__3 ;
    input WindowDin_0__0__2 ;
    input WindowDin_0__0__1 ;
    input WindowDin_0__0__0 ;
    input WindowDin_0__1__7 ;
    input WindowDin_0__1__6 ;
    input WindowDin_0__1__5 ;
    input WindowDin_0__1__4 ;
    input WindowDin_0__1__3 ;
    input WindowDin_0__1__2 ;
    input WindowDin_0__1__1 ;
    input WindowDin_0__1__0 ;
    input WindowDin_0__2__7 ;
    input WindowDin_0__2__6 ;
    input WindowDin_0__2__5 ;
    input WindowDin_0__2__4 ;
    input WindowDin_0__2__3 ;
    input WindowDin_0__2__2 ;
    input WindowDin_0__2__1 ;
    input WindowDin_0__2__0 ;
    input WindowDin_0__3__7 ;
    input WindowDin_0__3__6 ;
    input WindowDin_0__3__5 ;
    input WindowDin_0__3__4 ;
    input WindowDin_0__3__3 ;
    input WindowDin_0__3__2 ;
    input WindowDin_0__3__1 ;
    input WindowDin_0__3__0 ;
    input WindowDin_0__4__7 ;
    input WindowDin_0__4__6 ;
    input WindowDin_0__4__5 ;
    input WindowDin_0__4__4 ;
    input WindowDin_0__4__3 ;
    input WindowDin_0__4__2 ;
    input WindowDin_0__4__1 ;
    input WindowDin_0__4__0 ;
    input WindowDin_1__0__7 ;
    input WindowDin_1__0__6 ;
    input WindowDin_1__0__5 ;
    input WindowDin_1__0__4 ;
    input WindowDin_1__0__3 ;
    input WindowDin_1__0__2 ;
    input WindowDin_1__0__1 ;
    input WindowDin_1__0__0 ;
    input WindowDin_1__1__7 ;
    input WindowDin_1__1__6 ;
    input WindowDin_1__1__5 ;
    input WindowDin_1__1__4 ;
    input WindowDin_1__1__3 ;
    input WindowDin_1__1__2 ;
    input WindowDin_1__1__1 ;
    input WindowDin_1__1__0 ;
    input WindowDin_1__2__7 ;
    input WindowDin_1__2__6 ;
    input WindowDin_1__2__5 ;
    input WindowDin_1__2__4 ;
    input WindowDin_1__2__3 ;
    input WindowDin_1__2__2 ;
    input WindowDin_1__2__1 ;
    input WindowDin_1__2__0 ;
    input WindowDin_1__3__7 ;
    input WindowDin_1__3__6 ;
    input WindowDin_1__3__5 ;
    input WindowDin_1__3__4 ;
    input WindowDin_1__3__3 ;
    input WindowDin_1__3__2 ;
    input WindowDin_1__3__1 ;
    input WindowDin_1__3__0 ;
    input WindowDin_1__4__7 ;
    input WindowDin_1__4__6 ;
    input WindowDin_1__4__5 ;
    input WindowDin_1__4__4 ;
    input WindowDin_1__4__3 ;
    input WindowDin_1__4__2 ;
    input WindowDin_1__4__1 ;
    input WindowDin_1__4__0 ;
    input WindowDin_2__0__7 ;
    input WindowDin_2__0__6 ;
    input WindowDin_2__0__5 ;
    input WindowDin_2__0__4 ;
    input WindowDin_2__0__3 ;
    input WindowDin_2__0__2 ;
    input WindowDin_2__0__1 ;
    input WindowDin_2__0__0 ;
    input WindowDin_2__1__7 ;
    input WindowDin_2__1__6 ;
    input WindowDin_2__1__5 ;
    input WindowDin_2__1__4 ;
    input WindowDin_2__1__3 ;
    input WindowDin_2__1__2 ;
    input WindowDin_2__1__1 ;
    input WindowDin_2__1__0 ;
    input WindowDin_2__2__7 ;
    input WindowDin_2__2__6 ;
    input WindowDin_2__2__5 ;
    input WindowDin_2__2__4 ;
    input WindowDin_2__2__3 ;
    input WindowDin_2__2__2 ;
    input WindowDin_2__2__1 ;
    input WindowDin_2__2__0 ;
    input WindowDin_2__3__7 ;
    input WindowDin_2__3__6 ;
    input WindowDin_2__3__5 ;
    input WindowDin_2__3__4 ;
    input WindowDin_2__3__3 ;
    input WindowDin_2__3__2 ;
    input WindowDin_2__3__1 ;
    input WindowDin_2__3__0 ;
    input WindowDin_2__4__7 ;
    input WindowDin_2__4__6 ;
    input WindowDin_2__4__5 ;
    input WindowDin_2__4__4 ;
    input WindowDin_2__4__3 ;
    input WindowDin_2__4__2 ;
    input WindowDin_2__4__1 ;
    input WindowDin_2__4__0 ;
    input WindowDin_3__0__7 ;
    input WindowDin_3__0__6 ;
    input WindowDin_3__0__5 ;
    input WindowDin_3__0__4 ;
    input WindowDin_3__0__3 ;
    input WindowDin_3__0__2 ;
    input WindowDin_3__0__1 ;
    input WindowDin_3__0__0 ;
    input WindowDin_3__1__7 ;
    input WindowDin_3__1__6 ;
    input WindowDin_3__1__5 ;
    input WindowDin_3__1__4 ;
    input WindowDin_3__1__3 ;
    input WindowDin_3__1__2 ;
    input WindowDin_3__1__1 ;
    input WindowDin_3__1__0 ;
    input WindowDin_3__2__7 ;
    input WindowDin_3__2__6 ;
    input WindowDin_3__2__5 ;
    input WindowDin_3__2__4 ;
    input WindowDin_3__2__3 ;
    input WindowDin_3__2__2 ;
    input WindowDin_3__2__1 ;
    input WindowDin_3__2__0 ;
    input WindowDin_3__3__7 ;
    input WindowDin_3__3__6 ;
    input WindowDin_3__3__5 ;
    input WindowDin_3__3__4 ;
    input WindowDin_3__3__3 ;
    input WindowDin_3__3__2 ;
    input WindowDin_3__3__1 ;
    input WindowDin_3__3__0 ;
    input WindowDin_3__4__7 ;
    input WindowDin_3__4__6 ;
    input WindowDin_3__4__5 ;
    input WindowDin_3__4__4 ;
    input WindowDin_3__4__3 ;
    input WindowDin_3__4__2 ;
    input WindowDin_3__4__1 ;
    input WindowDin_3__4__0 ;
    input WindowDin_4__0__7 ;
    input WindowDin_4__0__6 ;
    input WindowDin_4__0__5 ;
    input WindowDin_4__0__4 ;
    input WindowDin_4__0__3 ;
    input WindowDin_4__0__2 ;
    input WindowDin_4__0__1 ;
    input WindowDin_4__0__0 ;
    input WindowDin_4__1__7 ;
    input WindowDin_4__1__6 ;
    input WindowDin_4__1__5 ;
    input WindowDin_4__1__4 ;
    input WindowDin_4__1__3 ;
    input WindowDin_4__1__2 ;
    input WindowDin_4__1__1 ;
    input WindowDin_4__1__0 ;
    input WindowDin_4__2__7 ;
    input WindowDin_4__2__6 ;
    input WindowDin_4__2__5 ;
    input WindowDin_4__2__4 ;
    input WindowDin_4__2__3 ;
    input WindowDin_4__2__2 ;
    input WindowDin_4__2__1 ;
    input WindowDin_4__2__0 ;
    input WindowDin_4__3__7 ;
    input WindowDin_4__3__6 ;
    input WindowDin_4__3__5 ;
    input WindowDin_4__3__4 ;
    input WindowDin_4__3__3 ;
    input WindowDin_4__3__2 ;
    input WindowDin_4__3__1 ;
    input WindowDin_4__3__0 ;
    input WindowDin_4__4__7 ;
    input WindowDin_4__4__6 ;
    input WindowDin_4__4__5 ;
    input WindowDin_4__4__4 ;
    input WindowDin_4__4__3 ;
    input WindowDin_4__4__2 ;
    input WindowDin_4__4__1 ;
    input WindowDin_4__4__0 ;
    output Done ;
    output [7:0]Result ;

    wire CounterEN, CounterRST, CalculatingBooth, CounterOut_3, CounterOut_2, 
         CounterOut_1, CounterOut_0, L1FirstOperands_0__7, L1FirstOperands_0__6, 
         L1FirstOperands_0__5, L1FirstOperands_0__4, L1FirstOperands_0__3, 
         L1FirstOperands_0__2, L1FirstOperands_0__1, L1FirstOperands_0__0, 
         L1FirstOperands_1__7, L1FirstOperands_1__6, L1FirstOperands_1__5, 
         L1FirstOperands_1__4, L1FirstOperands_1__3, L1FirstOperands_1__2, 
         L1FirstOperands_1__1, L1FirstOperands_1__0, L1FirstOperands_2__7, 
         L1FirstOperands_2__6, L1FirstOperands_2__5, L1FirstOperands_2__4, 
         L1FirstOperands_2__3, L1FirstOperands_2__2, L1FirstOperands_2__1, 
         L1FirstOperands_2__0, L1FirstOperands_3__7, L1FirstOperands_3__6, 
         L1FirstOperands_3__5, L1FirstOperands_3__4, L1FirstOperands_3__3, 
         L1FirstOperands_3__2, L1FirstOperands_3__1, L1FirstOperands_3__0, 
         L1FirstOperands_4__7, L1FirstOperands_4__6, L1FirstOperands_4__5, 
         L1FirstOperands_4__4, L1FirstOperands_4__3, L1FirstOperands_4__2, 
         L1FirstOperands_4__1, L1FirstOperands_4__0, L1FirstOperands_5__7, 
         L1FirstOperands_5__6, L1FirstOperands_5__5, L1FirstOperands_5__4, 
         L1FirstOperands_5__3, L1FirstOperands_5__2, L1FirstOperands_5__1, 
         L1FirstOperands_5__0, L1FirstOperands_6__7, L1FirstOperands_6__6, 
         L1FirstOperands_6__5, L1FirstOperands_6__4, L1FirstOperands_6__3, 
         L1FirstOperands_6__2, L1FirstOperands_6__1, L1FirstOperands_6__0, 
         L1FirstOperands_7__7, L1FirstOperands_7__6, L1FirstOperands_7__5, 
         L1FirstOperands_7__4, L1FirstOperands_7__3, L1FirstOperands_7__2, 
         L1FirstOperands_7__1, L1FirstOperands_7__0, L1FirstOperands_8__7, 
         L1FirstOperands_8__6, L1FirstOperands_8__5, L1FirstOperands_8__4, 
         L1FirstOperands_8__3, L1FirstOperands_8__2, L1FirstOperands_8__1, 
         L1FirstOperands_8__0, L1FirstOperands_9__7, L1FirstOperands_9__6, 
         L1FirstOperands_9__5, L1FirstOperands_9__4, L1FirstOperands_9__3, 
         L1FirstOperands_9__2, L1FirstOperands_9__1, L1FirstOperands_9__0, 
         L1FirstOperands_10__7, L1FirstOperands_10__6, L1FirstOperands_10__5, 
         L1FirstOperands_10__4, L1FirstOperands_10__3, L1FirstOperands_10__2, 
         L1FirstOperands_10__1, L1FirstOperands_10__0, L1FirstOperands_11__7, 
         L1FirstOperands_11__6, L1FirstOperands_11__5, L1FirstOperands_11__4, 
         L1FirstOperands_11__3, L1FirstOperands_11__2, L1FirstOperands_11__1, 
         L1FirstOperands_11__0, L1SecondOperands_0__7, L1SecondOperands_0__6, 
         L1SecondOperands_0__5, L1SecondOperands_0__4, L1SecondOperands_0__3, 
         L1SecondOperands_0__2, L1SecondOperands_0__1, L1SecondOperands_0__0, 
         L1SecondOperands_1__7, L1SecondOperands_1__6, L1SecondOperands_1__5, 
         L1SecondOperands_1__4, L1SecondOperands_1__3, L1SecondOperands_1__2, 
         L1SecondOperands_1__1, L1SecondOperands_1__0, L1SecondOperands_2__7, 
         L1SecondOperands_2__6, L1SecondOperands_2__5, L1SecondOperands_2__4, 
         L1SecondOperands_2__3, L1SecondOperands_2__2, L1SecondOperands_2__1, 
         L1SecondOperands_2__0, L1SecondOperands_3__7, L1SecondOperands_3__6, 
         L1SecondOperands_3__5, L1SecondOperands_3__4, L1SecondOperands_3__3, 
         L1SecondOperands_3__2, L1SecondOperands_3__1, L1SecondOperands_3__0, 
         L1SecondOperands_4__7, L1SecondOperands_4__6, L1SecondOperands_4__5, 
         L1SecondOperands_4__4, L1SecondOperands_4__3, L1SecondOperands_4__2, 
         L1SecondOperands_4__1, L1SecondOperands_4__0, L1SecondOperands_5__7, 
         L1SecondOperands_5__6, L1SecondOperands_5__5, L1SecondOperands_5__4, 
         L1SecondOperands_5__3, L1SecondOperands_5__2, L1SecondOperands_5__1, 
         L1SecondOperands_5__0, L1SecondOperands_6__7, L1SecondOperands_6__6, 
         L1SecondOperands_6__5, L1SecondOperands_6__4, L1SecondOperands_6__3, 
         L1SecondOperands_6__2, L1SecondOperands_6__1, L1SecondOperands_6__0, 
         L1SecondOperands_7__7, L1SecondOperands_7__6, L1SecondOperands_7__5, 
         L1SecondOperands_7__4, L1SecondOperands_7__3, L1SecondOperands_7__2, 
         L1SecondOperands_7__1, L1SecondOperands_7__0, L1SecondOperands_8__7, 
         L1SecondOperands_8__6, L1SecondOperands_8__5, L1SecondOperands_8__4, 
         L1SecondOperands_8__3, L1SecondOperands_8__2, L1SecondOperands_8__1, 
         L1SecondOperands_8__0, L1SecondOperands_9__7, L1SecondOperands_9__6, 
         L1SecondOperands_9__5, L1SecondOperands_9__4, L1SecondOperands_9__3, 
         L1SecondOperands_9__2, L1SecondOperands_9__1, L1SecondOperands_9__0, 
         L1SecondOperands_10__7, L1SecondOperands_10__6, L1SecondOperands_10__5, 
         L1SecondOperands_10__4, L1SecondOperands_10__3, L1SecondOperands_10__2, 
         L1SecondOperands_10__1, L1SecondOperands_10__0, L1SecondOperands_11__7, 
         L1SecondOperands_11__6, L1SecondOperands_11__5, L1SecondOperands_11__4, 
         L1SecondOperands_11__3, L1SecondOperands_11__2, L1SecondOperands_11__1, 
         L1SecondOperands_11__0, L1Results_0__7, L1Results_0__6, L1Results_0__5, 
         L1Results_0__4, L1Results_0__3, L1Results_0__2, L1Results_0__1, 
         L1Results_0__0, L1Results_1__7, L1Results_1__6, L1Results_1__5, 
         L1Results_1__4, L1Results_1__3, L1Results_1__2, L1Results_1__1, 
         L1Results_1__0, L1Results_2__7, L1Results_2__6, L1Results_2__5, 
         L1Results_2__4, L1Results_2__3, L1Results_2__2, L1Results_2__1, 
         L1Results_2__0, L1Results_3__7, L1Results_3__6, L1Results_3__5, 
         L1Results_3__4, L1Results_3__3, L1Results_3__2, L1Results_3__1, 
         L1Results_3__0, L1Results_4__7, L1Results_4__6, L1Results_4__5, 
         L1Results_4__4, L1Results_4__3, L1Results_4__2, L1Results_4__1, 
         L1Results_4__0, L1Results_5__7, L1Results_5__6, L1Results_5__5, 
         L1Results_5__4, L1Results_5__3, L1Results_5__2, L1Results_5__1, 
         L1Results_5__0, L1Results_6__7, L1Results_6__6, L1Results_6__5, 
         L1Results_6__4, L1Results_6__3, L1Results_6__2, L1Results_6__1, 
         L1Results_6__0, L1Results_7__7, L1Results_7__6, L1Results_7__5, 
         L1Results_7__4, L1Results_7__3, L1Results_7__2, L1Results_7__1, 
         L1Results_7__0, L1Results_8__7, L1Results_8__6, L1Results_8__5, 
         L1Results_8__4, L1Results_8__3, L1Results_8__2, L1Results_8__1, 
         L1Results_8__0, L1Results_9__7, L1Results_9__6, L1Results_9__5, 
         L1Results_9__4, L1Results_9__3, L1Results_9__2, L1Results_9__1, 
         L1Results_9__0, L1Results_10__7, L1Results_10__6, L1Results_10__5, 
         L1Results_10__4, L1Results_10__3, L1Results_10__2, L1Results_10__1, 
         L1Results_10__0, L1Results_11__7, L1Results_11__6, L1Results_11__5, 
         L1Results_11__4, L1Results_11__3, L1Results_11__2, L1Results_11__1, 
         L1Results_11__0, L2Results_0__7, L2Results_0__6, L2Results_0__5, 
         L2Results_0__4, L2Results_0__3, L2Results_0__2, L2Results_0__1, 
         L2Results_0__0, L2Results_1__7, L2Results_1__6, L2Results_1__5, 
         L2Results_1__4, L2Results_1__3, L2Results_1__2, L2Results_1__1, 
         L2Results_1__0, L2Results_2__7, L2Results_2__6, L2Results_2__5, 
         L2Results_2__4, L2Results_2__3, L2Results_2__2, L2Results_2__1, 
         L2Results_2__0, L2Results_3__7, L2Results_3__6, L2Results_3__5, 
         L2Results_3__4, L2Results_3__3, L2Results_3__2, L2Results_3__1, 
         L2Results_3__0, L2Results_4__7, L2Results_4__6, L2Results_4__5, 
         L2Results_4__4, L2Results_4__3, L2Results_4__2, L2Results_4__1, 
         L2Results_4__0, L2Results_5__7, L2Results_5__6, L2Results_5__5, 
         L2Results_5__4, L2Results_5__3, L2Results_5__2, L2Results_5__1, 
         L2Results_5__0, L3Results_0__7, L3Results_0__6, L3Results_0__5, 
         L3Results_0__4, L3Results_0__3, L3Results_0__2, L3Results_0__1, 
         L3Results_0__0, L3Results_1__7, L3Results_1__6, L3Results_1__5, 
         L3Results_1__4, L3Results_1__3, L3Results_1__2, L3Results_1__1, 
         L3Results_1__0, L3Results_2__7, L3Results_2__6, L3Results_2__5, 
         L3Results_2__4, L3Results_2__3, L3Results_2__2, L3Results_2__1, 
         L3Results_2__0, L4Results_0__7, L4Results_0__6, L4Results_0__5, 
         L4Results_0__4, L4Results_0__3, L4Results_0__2, L4Results_0__1, 
         L4Results_0__0, L5FirstOperands_1__7, L5FirstOperands_1__6, 
         L5FirstOperands_1__5, L5FirstOperands_1__4, L5FirstOperands_1__3, 
         L5FirstOperands_1__2, L5FirstOperands_1__1, L5FirstOperands_1__0, 
         L5SecondOperands_1__7, L5SecondOperands_1__6, L5SecondOperands_1__5, 
         L5SecondOperands_1__4, L5SecondOperands_1__3, L5SecondOperands_1__2, 
         L5SecondOperands_1__1, L5SecondOperands_1__0, L5Results_1__7, 
         L5Results_1__6, L5Results_1__5, L5Results_1__4, L5Results_1__3, 
         L5Results_1__2, L5Results_1__1, L5Results_1__0, nx22, nx78, nx990, 
         nx993, nx995, nx1001, nx1003, nx1007, nx1009, nx1012, nx1014, nx1043, 
         CalculatingBooth_dup_1084, CalculatingBooth_dup_1119, 
         CalculatingBooth_dup_1162, CalculatingBooth_dup_1253, 
         ACCELERATOR_COUNTER_nx6, ACCELERATOR_COUNTER_nx12, 
         ACCELERATOR_COUNTER_nx18, ACCELERATOR_COUNTER_nx81, 
         ACCELERATOR_COUNTER_nx91, ACCELERATOR_COUNTER_nx101, 
         ACCELERATOR_COUNTER_nx111, ACCELERATOR_COUNTER_nx133, 
         ACCELERATOR_COUNTER_nx139, L1_0_L2_0_G1_MINI_ALU_AddPToBoothOperand, 
         L1_0_L2_0_G1_MINI_ALU_BoothOperand_16, 
         L1_0_L2_0_G1_MINI_ALU_BoothOperand_15, 
         L1_0_L2_0_G1_MINI_ALU_BoothOperand_14, 
         L1_0_L2_0_G1_MINI_ALU_BoothOperand_13, 
         L1_0_L2_0_G1_MINI_ALU_BoothOperand_12, 
         L1_0_L2_0_G1_MINI_ALU_BoothOperand_11, 
         L1_0_L2_0_G1_MINI_ALU_BoothOperand_10, 
         L1_0_L2_0_G1_MINI_ALU_BoothOperand_9, 
         L1_0_L2_0_G1_MINI_ALU_BoothOperand_8, 
         L1_0_L2_0_G1_MINI_ALU_BoothOperand_7, 
         L1_0_L2_0_G1_MINI_ALU_BoothOperand_6, 
         L1_0_L2_0_G1_MINI_ALU_BoothOperand_5, 
         L1_0_L2_0_G1_MINI_ALU_BoothOperand_4, 
         L1_0_L2_0_G1_MINI_ALU_BoothOperand_3, 
         L1_0_L2_0_G1_MINI_ALU_BoothOperand_2, 
         L1_0_L2_0_G1_MINI_ALU_BoothOperand_1, 
         L1_0_L2_0_G1_MINI_ALU_BoothOperand_0, 
         L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_16, 
         L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_15, 
         L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_14, 
         L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_13, 
         L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_12, 
         L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_11, 
         L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_10, 
         L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_9, 
         L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_8, 
         L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_7, 
         L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_6, 
         L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_5, 
         L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_4, 
         L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_3, 
         L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_2, 
         L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_1, 
         L1_0_L2_0_G1_MINI_ALU_BoothP_16, L1_0_L2_0_G1_MINI_ALU_BoothP_15, 
         L1_0_L2_0_G1_MINI_ALU_BoothP_14, L1_0_L2_0_G1_MINI_ALU_BoothP_13, 
         L1_0_L2_0_G1_MINI_ALU_BoothP_12, L1_0_L2_0_G1_MINI_ALU_BoothP_11, 
         L1_0_L2_0_G1_MINI_ALU_BoothP_10, L1_0_L2_0_G1_MINI_ALU_BoothP_9, 
         L1_0_L2_0_G1_MINI_ALU_BoothP_8, L1_0_L2_0_G1_MINI_ALU_BoothP_7, 
         L1_0_L2_0_G1_MINI_ALU_BoothP_6, L1_0_L2_0_G1_MINI_ALU_BoothP_5, 
         L1_0_L2_0_G1_MINI_ALU_BoothP_4, L1_0_L2_0_G1_MINI_ALU_BoothP_3, 
         L1_0_L2_0_G1_MINI_ALU_BoothP_2, L1_0_L2_0_G1_MINI_ALU_BoothP_1, 
         L1_0_L2_0_G1_MINI_ALU_BoothP_0, L1_0_L2_0_G1_MINI_ALU_nx0, 
         L1_0_L2_0_G1_MINI_ALU_nx6, L1_0_L2_0_G1_MINI_ALU_nx12, 
         L1_0_L2_0_G1_MINI_ALU_nx18, L1_0_L2_0_G1_MINI_ALU_nx24, 
         L1_0_L2_0_G1_MINI_ALU_nx30, L1_0_L2_0_G1_MINI_ALU_nx40, 
         L1_0_L2_0_G1_MINI_ALU_nx44, L1_0_L2_0_G1_MINI_ALU_nx48, 
         L1_0_L2_0_G1_MINI_ALU_nx52, L1_0_L2_0_G1_MINI_ALU_nx56, 
         L1_0_L2_0_G1_MINI_ALU_nx62, L1_0_L2_0_G1_MINI_ALU_nx154, 
         L1_0_L2_0_G1_MINI_ALU_nx316, L1_0_L2_0_G1_MINI_ALU_nx336, 
         L1_0_L2_0_G1_MINI_ALU_nx356, L1_0_L2_0_G1_MINI_ALU_nx376, 
         L1_0_L2_0_G1_MINI_ALU_nx396, L1_0_L2_0_G1_MINI_ALU_nx416, 
         L1_0_L2_0_G1_MINI_ALU_nx436, L1_0_L2_0_G1_MINI_ALU_nx454, 
         L1_0_L2_0_G1_MINI_ALU_nx456, L1_0_L2_0_G1_MINI_ALU_nx379, 
         L1_0_L2_0_G1_MINI_ALU_nx381, L1_0_L2_0_G1_MINI_ALU_nx383, 
         L1_0_L2_0_G1_MINI_ALU_nx387, L1_0_L2_0_G1_MINI_ALU_nx389, 
         L1_0_L2_0_G1_MINI_ALU_nx391, L1_0_L2_0_G1_MINI_ALU_nx395, 
         L1_0_L2_0_G1_MINI_ALU_nx399, L1_0_L2_0_G1_MINI_ALU_nx401, 
         L1_0_L2_0_G1_MINI_ALU_nx403, L1_0_L2_0_G1_MINI_ALU_nx405, 
         L1_0_L2_0_G1_MINI_ALU_nx409, L1_0_L2_0_G1_MINI_ALU_nx411, 
         L1_0_L2_0_G1_MINI_ALU_nx413, L1_0_L2_0_G1_MINI_ALU_nx415, 
         L1_0_L2_0_G1_MINI_ALU_nx419, L1_0_L2_0_G1_MINI_ALU_nx421, 
         L1_0_L2_0_G1_MINI_ALU_nx423, L1_0_L2_0_G1_MINI_ALU_nx425, 
         L1_0_L2_0_G1_MINI_ALU_nx429, L1_0_L2_0_G1_MINI_ALU_nx431, 
         L1_0_L2_0_G1_MINI_ALU_nx433, L1_0_L2_0_G1_MINI_ALU_nx435, 
         L1_0_L2_0_G1_MINI_ALU_nx439, L1_0_L2_0_G1_MINI_ALU_nx441, 
         L1_0_L2_0_G1_MINI_ALU_nx443, L1_0_L2_0_G1_MINI_ALU_nx445, 
         L1_0_L2_0_G1_MINI_ALU_nx449, L1_0_L2_0_G1_MINI_ALU_nx451, 
         L1_0_L2_0_G1_MINI_ALU_nx453, L1_0_L2_0_G1_MINI_ALU_nx455, 
         L1_0_L2_0_G1_MINI_ALU_nx461, L1_0_L2_0_G1_MINI_ALU_nx463, 
         L1_0_L2_0_G1_MINI_ALU_nx467, L1_0_L2_0_G1_MINI_ALU_nx469, 
         L1_0_L2_0_G1_MINI_ALU_nx471, L1_0_L2_0_G1_MINI_ALU_nx475, 
         L1_0_L2_0_G1_MINI_ALU_nx477, L1_0_L2_0_G1_MINI_ALU_nx479, 
         L1_0_L2_0_G1_MINI_ALU_nx483, L1_0_L2_0_G1_MINI_ALU_nx485, 
         L1_0_L2_0_G1_MINI_ALU_nx487, L1_0_L2_0_G1_MINI_ALU_nx491, 
         L1_0_L2_0_G1_MINI_ALU_nx493, L1_0_L2_0_G1_MINI_ALU_nx495, 
         L1_0_L2_0_G1_MINI_ALU_nx499, L1_0_L2_0_G1_MINI_ALU_nx501, 
         L1_0_L2_0_G1_MINI_ALU_nx503, L1_0_L2_0_G1_MINI_ALU_nx507, 
         L1_0_L2_0_G1_MINI_ALU_nx509, L1_0_L2_0_G1_MINI_ALU_nx511, 
         L1_0_L2_0_G1_MINI_ALU_nx515, L1_0_L2_0_G1_MINI_ALU_nx517, 
         L1_0_L2_0_G1_MINI_ALU_nx529, L1_0_L2_0_G1_MINI_ALU_nx531, 
         L1_0_L2_0_G1_MINI_ALU_nx534, L1_0_L2_0_G1_MINI_ALU_nx537, 
         L1_0_L2_0_G1_MINI_ALU_nx540, L1_0_L2_0_G1_MINI_ALU_nx544, 
         L1_0_L2_0_G1_MINI_ALU_nx547, L1_0_L2_0_G1_MINI_ALU_nx551, 
         L1_0_L2_0_G1_MINI_ALU_nx554, L1_0_L2_0_G1_MINI_ALU_nx558, 
         L1_0_L2_0_G1_MINI_ALU_nx561, L1_0_L2_0_G1_MINI_ALU_nx565, 
         L1_0_L2_0_G1_MINI_ALU_nx568, 
         L1_0_L2_0_G1_MINI_ALU_WindowCellShiftedLeft_16, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_16, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_15, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_14, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_13, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_12, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_11, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_10, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_16, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_15, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_14, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_13, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_12, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_11, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_10, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_9, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_8, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_7, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_6, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_5, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_4, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_3, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_2, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_1, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_0, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_16, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_15, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_14, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_13, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_12, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_11, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_10, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_9, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_8, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_7, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_6, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_5, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_4, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_3, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_2, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_1, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_0, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_16, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_15, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_14, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_13, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_12, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_11, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_10, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_9, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_8, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_7, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_6, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_5, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_4, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_3, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_2, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_1, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_0, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx4, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx8, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx12, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx16, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx20, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx24, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx80, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx328, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx384, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx564, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642, 
         L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644, 
         L1_0_L2_1_G1_MINI_ALU_AddPToBoothOperand, 
         L1_0_L2_1_G1_MINI_ALU_BoothOperand_16, 
         L1_0_L2_1_G1_MINI_ALU_BoothOperand_15, 
         L1_0_L2_1_G1_MINI_ALU_BoothOperand_14, 
         L1_0_L2_1_G1_MINI_ALU_BoothOperand_13, 
         L1_0_L2_1_G1_MINI_ALU_BoothOperand_12, 
         L1_0_L2_1_G1_MINI_ALU_BoothOperand_11, 
         L1_0_L2_1_G1_MINI_ALU_BoothOperand_10, 
         L1_0_L2_1_G1_MINI_ALU_BoothOperand_9, 
         L1_0_L2_1_G1_MINI_ALU_BoothOperand_8, 
         L1_0_L2_1_G1_MINI_ALU_BoothOperand_7, 
         L1_0_L2_1_G1_MINI_ALU_BoothOperand_6, 
         L1_0_L2_1_G1_MINI_ALU_BoothOperand_5, 
         L1_0_L2_1_G1_MINI_ALU_BoothOperand_4, 
         L1_0_L2_1_G1_MINI_ALU_BoothOperand_3, 
         L1_0_L2_1_G1_MINI_ALU_BoothOperand_2, 
         L1_0_L2_1_G1_MINI_ALU_BoothOperand_1, 
         L1_0_L2_1_G1_MINI_ALU_BoothOperand_0, 
         L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_16, 
         L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_15, 
         L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_14, 
         L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_13, 
         L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_12, 
         L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_11, 
         L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_10, 
         L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_9, 
         L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_8, 
         L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_7, 
         L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_6, 
         L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_5, 
         L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_4, 
         L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_3, 
         L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_2, 
         L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_1, 
         L1_0_L2_1_G1_MINI_ALU_BoothP_16, L1_0_L2_1_G1_MINI_ALU_BoothP_15, 
         L1_0_L2_1_G1_MINI_ALU_BoothP_14, L1_0_L2_1_G1_MINI_ALU_BoothP_13, 
         L1_0_L2_1_G1_MINI_ALU_BoothP_12, L1_0_L2_1_G1_MINI_ALU_BoothP_11, 
         L1_0_L2_1_G1_MINI_ALU_BoothP_10, L1_0_L2_1_G1_MINI_ALU_BoothP_9, 
         L1_0_L2_1_G1_MINI_ALU_BoothP_8, L1_0_L2_1_G1_MINI_ALU_BoothP_7, 
         L1_0_L2_1_G1_MINI_ALU_BoothP_6, L1_0_L2_1_G1_MINI_ALU_BoothP_5, 
         L1_0_L2_1_G1_MINI_ALU_BoothP_4, L1_0_L2_1_G1_MINI_ALU_BoothP_3, 
         L1_0_L2_1_G1_MINI_ALU_BoothP_2, L1_0_L2_1_G1_MINI_ALU_BoothP_1, 
         L1_0_L2_1_G1_MINI_ALU_BoothP_0, L1_0_L2_1_G1_MINI_ALU_nx0, 
         L1_0_L2_1_G1_MINI_ALU_nx6, L1_0_L2_1_G1_MINI_ALU_nx12, 
         L1_0_L2_1_G1_MINI_ALU_nx18, L1_0_L2_1_G1_MINI_ALU_nx24, 
         L1_0_L2_1_G1_MINI_ALU_nx30, L1_0_L2_1_G1_MINI_ALU_nx40, 
         L1_0_L2_1_G1_MINI_ALU_nx44, L1_0_L2_1_G1_MINI_ALU_nx48, 
         L1_0_L2_1_G1_MINI_ALU_nx52, L1_0_L2_1_G1_MINI_ALU_nx56, 
         L1_0_L2_1_G1_MINI_ALU_nx62, L1_0_L2_1_G1_MINI_ALU_nx154, 
         L1_0_L2_1_G1_MINI_ALU_nx316, L1_0_L2_1_G1_MINI_ALU_nx336, 
         L1_0_L2_1_G1_MINI_ALU_nx356, L1_0_L2_1_G1_MINI_ALU_nx376, 
         L1_0_L2_1_G1_MINI_ALU_nx396, L1_0_L2_1_G1_MINI_ALU_nx416, 
         L1_0_L2_1_G1_MINI_ALU_nx436, L1_0_L2_1_G1_MINI_ALU_nx454, 
         L1_0_L2_1_G1_MINI_ALU_nx456, L1_0_L2_1_G1_MINI_ALU_nx379, 
         L1_0_L2_1_G1_MINI_ALU_nx381, L1_0_L2_1_G1_MINI_ALU_nx383, 
         L1_0_L2_1_G1_MINI_ALU_nx387, L1_0_L2_1_G1_MINI_ALU_nx389, 
         L1_0_L2_1_G1_MINI_ALU_nx391, L1_0_L2_1_G1_MINI_ALU_nx395, 
         L1_0_L2_1_G1_MINI_ALU_nx399, L1_0_L2_1_G1_MINI_ALU_nx401, 
         L1_0_L2_1_G1_MINI_ALU_nx403, L1_0_L2_1_G1_MINI_ALU_nx405, 
         L1_0_L2_1_G1_MINI_ALU_nx409, L1_0_L2_1_G1_MINI_ALU_nx411, 
         L1_0_L2_1_G1_MINI_ALU_nx413, L1_0_L2_1_G1_MINI_ALU_nx415, 
         L1_0_L2_1_G1_MINI_ALU_nx419, L1_0_L2_1_G1_MINI_ALU_nx421, 
         L1_0_L2_1_G1_MINI_ALU_nx423, L1_0_L2_1_G1_MINI_ALU_nx425, 
         L1_0_L2_1_G1_MINI_ALU_nx429, L1_0_L2_1_G1_MINI_ALU_nx431, 
         L1_0_L2_1_G1_MINI_ALU_nx433, L1_0_L2_1_G1_MINI_ALU_nx435, 
         L1_0_L2_1_G1_MINI_ALU_nx439, L1_0_L2_1_G1_MINI_ALU_nx441, 
         L1_0_L2_1_G1_MINI_ALU_nx443, L1_0_L2_1_G1_MINI_ALU_nx445, 
         L1_0_L2_1_G1_MINI_ALU_nx449, L1_0_L2_1_G1_MINI_ALU_nx451, 
         L1_0_L2_1_G1_MINI_ALU_nx453, L1_0_L2_1_G1_MINI_ALU_nx455, 
         L1_0_L2_1_G1_MINI_ALU_nx461, L1_0_L2_1_G1_MINI_ALU_nx463, 
         L1_0_L2_1_G1_MINI_ALU_nx467, L1_0_L2_1_G1_MINI_ALU_nx469, 
         L1_0_L2_1_G1_MINI_ALU_nx471, L1_0_L2_1_G1_MINI_ALU_nx475, 
         L1_0_L2_1_G1_MINI_ALU_nx477, L1_0_L2_1_G1_MINI_ALU_nx479, 
         L1_0_L2_1_G1_MINI_ALU_nx483, L1_0_L2_1_G1_MINI_ALU_nx485, 
         L1_0_L2_1_G1_MINI_ALU_nx487, L1_0_L2_1_G1_MINI_ALU_nx491, 
         L1_0_L2_1_G1_MINI_ALU_nx493, L1_0_L2_1_G1_MINI_ALU_nx495, 
         L1_0_L2_1_G1_MINI_ALU_nx499, L1_0_L2_1_G1_MINI_ALU_nx501, 
         L1_0_L2_1_G1_MINI_ALU_nx503, L1_0_L2_1_G1_MINI_ALU_nx507, 
         L1_0_L2_1_G1_MINI_ALU_nx509, L1_0_L2_1_G1_MINI_ALU_nx511, 
         L1_0_L2_1_G1_MINI_ALU_nx515, L1_0_L2_1_G1_MINI_ALU_nx517, 
         L1_0_L2_1_G1_MINI_ALU_nx529, L1_0_L2_1_G1_MINI_ALU_nx531, 
         L1_0_L2_1_G1_MINI_ALU_nx534, L1_0_L2_1_G1_MINI_ALU_nx537, 
         L1_0_L2_1_G1_MINI_ALU_nx540, L1_0_L2_1_G1_MINI_ALU_nx544, 
         L1_0_L2_1_G1_MINI_ALU_nx547, L1_0_L2_1_G1_MINI_ALU_nx551, 
         L1_0_L2_1_G1_MINI_ALU_nx554, L1_0_L2_1_G1_MINI_ALU_nx558, 
         L1_0_L2_1_G1_MINI_ALU_nx561, L1_0_L2_1_G1_MINI_ALU_nx565, 
         L1_0_L2_1_G1_MINI_ALU_nx568, 
         L1_0_L2_1_G1_MINI_ALU_WindowCellShiftedLeft_16, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_16, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_15, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_14, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_13, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_12, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_11, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_10, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_16, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_15, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_14, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_13, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_12, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_11, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_10, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_9, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_8, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_7, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_6, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_5, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_4, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_3, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_2, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_1, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_0, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_16, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_15, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_14, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_13, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_12, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_11, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_10, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_9, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_8, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_7, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_6, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_5, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_4, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_3, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_2, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_1, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_0, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_16, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_15, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_14, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_13, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_12, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_11, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_10, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_9, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_8, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_7, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_6, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_5, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_4, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_3, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_2, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_1, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_0, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx4, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx8, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx12, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx16, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx20, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx24, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx80, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx328, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx384, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642, 
         L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644, 
         L1_0_L2_2_G1_MINI_ALU_AddPToBoothOperand, 
         L1_0_L2_2_G1_MINI_ALU_BoothOperand_16, 
         L1_0_L2_2_G1_MINI_ALU_BoothOperand_15, 
         L1_0_L2_2_G1_MINI_ALU_BoothOperand_14, 
         L1_0_L2_2_G1_MINI_ALU_BoothOperand_13, 
         L1_0_L2_2_G1_MINI_ALU_BoothOperand_12, 
         L1_0_L2_2_G1_MINI_ALU_BoothOperand_11, 
         L1_0_L2_2_G1_MINI_ALU_BoothOperand_10, 
         L1_0_L2_2_G1_MINI_ALU_BoothOperand_9, 
         L1_0_L2_2_G1_MINI_ALU_BoothOperand_8, 
         L1_0_L2_2_G1_MINI_ALU_BoothOperand_7, 
         L1_0_L2_2_G1_MINI_ALU_BoothOperand_6, 
         L1_0_L2_2_G1_MINI_ALU_BoothOperand_5, 
         L1_0_L2_2_G1_MINI_ALU_BoothOperand_4, 
         L1_0_L2_2_G1_MINI_ALU_BoothOperand_3, 
         L1_0_L2_2_G1_MINI_ALU_BoothOperand_2, 
         L1_0_L2_2_G1_MINI_ALU_BoothOperand_1, 
         L1_0_L2_2_G1_MINI_ALU_BoothOperand_0, 
         L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_16, 
         L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_15, 
         L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_14, 
         L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_13, 
         L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_12, 
         L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_11, 
         L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_10, 
         L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_9, 
         L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_8, 
         L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_7, 
         L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_6, 
         L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_5, 
         L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_4, 
         L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_3, 
         L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_2, 
         L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_1, 
         L1_0_L2_2_G1_MINI_ALU_BoothP_16, L1_0_L2_2_G1_MINI_ALU_BoothP_15, 
         L1_0_L2_2_G1_MINI_ALU_BoothP_14, L1_0_L2_2_G1_MINI_ALU_BoothP_13, 
         L1_0_L2_2_G1_MINI_ALU_BoothP_12, L1_0_L2_2_G1_MINI_ALU_BoothP_11, 
         L1_0_L2_2_G1_MINI_ALU_BoothP_10, L1_0_L2_2_G1_MINI_ALU_BoothP_9, 
         L1_0_L2_2_G1_MINI_ALU_BoothP_8, L1_0_L2_2_G1_MINI_ALU_BoothP_7, 
         L1_0_L2_2_G1_MINI_ALU_BoothP_6, L1_0_L2_2_G1_MINI_ALU_BoothP_5, 
         L1_0_L2_2_G1_MINI_ALU_BoothP_4, L1_0_L2_2_G1_MINI_ALU_BoothP_3, 
         L1_0_L2_2_G1_MINI_ALU_BoothP_2, L1_0_L2_2_G1_MINI_ALU_BoothP_1, 
         L1_0_L2_2_G1_MINI_ALU_BoothP_0, L1_0_L2_2_G1_MINI_ALU_nx0, 
         L1_0_L2_2_G1_MINI_ALU_nx6, L1_0_L2_2_G1_MINI_ALU_nx12, 
         L1_0_L2_2_G1_MINI_ALU_nx18, L1_0_L2_2_G1_MINI_ALU_nx24, 
         L1_0_L2_2_G1_MINI_ALU_nx30, L1_0_L2_2_G1_MINI_ALU_nx40, 
         L1_0_L2_2_G1_MINI_ALU_nx44, L1_0_L2_2_G1_MINI_ALU_nx48, 
         L1_0_L2_2_G1_MINI_ALU_nx52, L1_0_L2_2_G1_MINI_ALU_nx56, 
         L1_0_L2_2_G1_MINI_ALU_nx62, L1_0_L2_2_G1_MINI_ALU_nx154, 
         L1_0_L2_2_G1_MINI_ALU_nx316, L1_0_L2_2_G1_MINI_ALU_nx336, 
         L1_0_L2_2_G1_MINI_ALU_nx356, L1_0_L2_2_G1_MINI_ALU_nx376, 
         L1_0_L2_2_G1_MINI_ALU_nx396, L1_0_L2_2_G1_MINI_ALU_nx416, 
         L1_0_L2_2_G1_MINI_ALU_nx436, L1_0_L2_2_G1_MINI_ALU_nx454, 
         L1_0_L2_2_G1_MINI_ALU_nx456, L1_0_L2_2_G1_MINI_ALU_nx379, 
         L1_0_L2_2_G1_MINI_ALU_nx381, L1_0_L2_2_G1_MINI_ALU_nx383, 
         L1_0_L2_2_G1_MINI_ALU_nx387, L1_0_L2_2_G1_MINI_ALU_nx389, 
         L1_0_L2_2_G1_MINI_ALU_nx391, L1_0_L2_2_G1_MINI_ALU_nx395, 
         L1_0_L2_2_G1_MINI_ALU_nx399, L1_0_L2_2_G1_MINI_ALU_nx401, 
         L1_0_L2_2_G1_MINI_ALU_nx403, L1_0_L2_2_G1_MINI_ALU_nx405, 
         L1_0_L2_2_G1_MINI_ALU_nx409, L1_0_L2_2_G1_MINI_ALU_nx411, 
         L1_0_L2_2_G1_MINI_ALU_nx413, L1_0_L2_2_G1_MINI_ALU_nx415, 
         L1_0_L2_2_G1_MINI_ALU_nx419, L1_0_L2_2_G1_MINI_ALU_nx421, 
         L1_0_L2_2_G1_MINI_ALU_nx423, L1_0_L2_2_G1_MINI_ALU_nx425, 
         L1_0_L2_2_G1_MINI_ALU_nx429, L1_0_L2_2_G1_MINI_ALU_nx431, 
         L1_0_L2_2_G1_MINI_ALU_nx433, L1_0_L2_2_G1_MINI_ALU_nx435, 
         L1_0_L2_2_G1_MINI_ALU_nx439, L1_0_L2_2_G1_MINI_ALU_nx441, 
         L1_0_L2_2_G1_MINI_ALU_nx443, L1_0_L2_2_G1_MINI_ALU_nx445, 
         L1_0_L2_2_G1_MINI_ALU_nx449, L1_0_L2_2_G1_MINI_ALU_nx451, 
         L1_0_L2_2_G1_MINI_ALU_nx453, L1_0_L2_2_G1_MINI_ALU_nx455, 
         L1_0_L2_2_G1_MINI_ALU_nx461, L1_0_L2_2_G1_MINI_ALU_nx463, 
         L1_0_L2_2_G1_MINI_ALU_nx467, L1_0_L2_2_G1_MINI_ALU_nx469, 
         L1_0_L2_2_G1_MINI_ALU_nx471, L1_0_L2_2_G1_MINI_ALU_nx475, 
         L1_0_L2_2_G1_MINI_ALU_nx477, L1_0_L2_2_G1_MINI_ALU_nx479, 
         L1_0_L2_2_G1_MINI_ALU_nx483, L1_0_L2_2_G1_MINI_ALU_nx485, 
         L1_0_L2_2_G1_MINI_ALU_nx487, L1_0_L2_2_G1_MINI_ALU_nx491, 
         L1_0_L2_2_G1_MINI_ALU_nx493, L1_0_L2_2_G1_MINI_ALU_nx495, 
         L1_0_L2_2_G1_MINI_ALU_nx499, L1_0_L2_2_G1_MINI_ALU_nx501, 
         L1_0_L2_2_G1_MINI_ALU_nx503, L1_0_L2_2_G1_MINI_ALU_nx507, 
         L1_0_L2_2_G1_MINI_ALU_nx509, L1_0_L2_2_G1_MINI_ALU_nx511, 
         L1_0_L2_2_G1_MINI_ALU_nx515, L1_0_L2_2_G1_MINI_ALU_nx517, 
         L1_0_L2_2_G1_MINI_ALU_nx529, L1_0_L2_2_G1_MINI_ALU_nx531, 
         L1_0_L2_2_G1_MINI_ALU_nx534, L1_0_L2_2_G1_MINI_ALU_nx537, 
         L1_0_L2_2_G1_MINI_ALU_nx540, L1_0_L2_2_G1_MINI_ALU_nx544, 
         L1_0_L2_2_G1_MINI_ALU_nx547, L1_0_L2_2_G1_MINI_ALU_nx551, 
         L1_0_L2_2_G1_MINI_ALU_nx554, L1_0_L2_2_G1_MINI_ALU_nx558, 
         L1_0_L2_2_G1_MINI_ALU_nx561, L1_0_L2_2_G1_MINI_ALU_nx565, 
         L1_0_L2_2_G1_MINI_ALU_nx568, 
         L1_0_L2_2_G1_MINI_ALU_WindowCellShiftedLeft_16, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_16, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_15, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_14, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_13, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_12, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_11, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_10, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_16, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_15, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_14, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_13, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_12, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_11, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_10, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_9, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_8, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_7, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_6, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_5, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_4, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_3, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_2, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_1, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_0, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_16, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_15, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_14, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_13, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_12, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_11, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_10, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_9, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_8, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_7, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_6, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_5, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_4, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_3, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_2, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_1, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_0, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_16, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_15, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_14, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_13, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_12, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_11, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_10, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_9, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_8, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_7, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_6, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_5, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_4, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_3, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_2, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_1, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_0, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx4, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx8, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx12, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx16, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx20, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx24, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx80, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx328, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx384, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642, 
         L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644, 
         L1_0_L2_3_G1_MINI_ALU_AddPToBoothOperand, 
         L1_0_L2_3_G1_MINI_ALU_BoothOperand_16, 
         L1_0_L2_3_G1_MINI_ALU_BoothOperand_15, 
         L1_0_L2_3_G1_MINI_ALU_BoothOperand_14, 
         L1_0_L2_3_G1_MINI_ALU_BoothOperand_13, 
         L1_0_L2_3_G1_MINI_ALU_BoothOperand_12, 
         L1_0_L2_3_G1_MINI_ALU_BoothOperand_11, 
         L1_0_L2_3_G1_MINI_ALU_BoothOperand_10, 
         L1_0_L2_3_G1_MINI_ALU_BoothOperand_9, 
         L1_0_L2_3_G1_MINI_ALU_BoothOperand_8, 
         L1_0_L2_3_G1_MINI_ALU_BoothOperand_7, 
         L1_0_L2_3_G1_MINI_ALU_BoothOperand_6, 
         L1_0_L2_3_G1_MINI_ALU_BoothOperand_5, 
         L1_0_L2_3_G1_MINI_ALU_BoothOperand_4, 
         L1_0_L2_3_G1_MINI_ALU_BoothOperand_3, 
         L1_0_L2_3_G1_MINI_ALU_BoothOperand_2, 
         L1_0_L2_3_G1_MINI_ALU_BoothOperand_1, 
         L1_0_L2_3_G1_MINI_ALU_BoothOperand_0, 
         L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_16, 
         L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_15, 
         L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_14, 
         L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_13, 
         L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_12, 
         L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_11, 
         L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_10, 
         L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_9, 
         L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_8, 
         L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_7, 
         L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_6, 
         L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_5, 
         L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_4, 
         L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_3, 
         L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_2, 
         L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_1, 
         L1_0_L2_3_G1_MINI_ALU_BoothP_16, L1_0_L2_3_G1_MINI_ALU_BoothP_15, 
         L1_0_L2_3_G1_MINI_ALU_BoothP_14, L1_0_L2_3_G1_MINI_ALU_BoothP_13, 
         L1_0_L2_3_G1_MINI_ALU_BoothP_12, L1_0_L2_3_G1_MINI_ALU_BoothP_11, 
         L1_0_L2_3_G1_MINI_ALU_BoothP_10, L1_0_L2_3_G1_MINI_ALU_BoothP_9, 
         L1_0_L2_3_G1_MINI_ALU_BoothP_8, L1_0_L2_3_G1_MINI_ALU_BoothP_7, 
         L1_0_L2_3_G1_MINI_ALU_BoothP_6, L1_0_L2_3_G1_MINI_ALU_BoothP_5, 
         L1_0_L2_3_G1_MINI_ALU_BoothP_4, L1_0_L2_3_G1_MINI_ALU_BoothP_3, 
         L1_0_L2_3_G1_MINI_ALU_BoothP_2, L1_0_L2_3_G1_MINI_ALU_BoothP_1, 
         L1_0_L2_3_G1_MINI_ALU_BoothP_0, L1_0_L2_3_G1_MINI_ALU_nx0, 
         L1_0_L2_3_G1_MINI_ALU_nx6, L1_0_L2_3_G1_MINI_ALU_nx12, 
         L1_0_L2_3_G1_MINI_ALU_nx18, L1_0_L2_3_G1_MINI_ALU_nx24, 
         L1_0_L2_3_G1_MINI_ALU_nx30, L1_0_L2_3_G1_MINI_ALU_nx40, 
         L1_0_L2_3_G1_MINI_ALU_nx44, L1_0_L2_3_G1_MINI_ALU_nx48, 
         L1_0_L2_3_G1_MINI_ALU_nx52, L1_0_L2_3_G1_MINI_ALU_nx56, 
         L1_0_L2_3_G1_MINI_ALU_nx62, L1_0_L2_3_G1_MINI_ALU_nx154, 
         L1_0_L2_3_G1_MINI_ALU_nx316, L1_0_L2_3_G1_MINI_ALU_nx336, 
         L1_0_L2_3_G1_MINI_ALU_nx356, L1_0_L2_3_G1_MINI_ALU_nx376, 
         L1_0_L2_3_G1_MINI_ALU_nx396, L1_0_L2_3_G1_MINI_ALU_nx416, 
         L1_0_L2_3_G1_MINI_ALU_nx436, L1_0_L2_3_G1_MINI_ALU_nx454, 
         L1_0_L2_3_G1_MINI_ALU_nx456, L1_0_L2_3_G1_MINI_ALU_nx379, 
         L1_0_L2_3_G1_MINI_ALU_nx381, L1_0_L2_3_G1_MINI_ALU_nx383, 
         L1_0_L2_3_G1_MINI_ALU_nx387, L1_0_L2_3_G1_MINI_ALU_nx389, 
         L1_0_L2_3_G1_MINI_ALU_nx391, L1_0_L2_3_G1_MINI_ALU_nx395, 
         L1_0_L2_3_G1_MINI_ALU_nx399, L1_0_L2_3_G1_MINI_ALU_nx401, 
         L1_0_L2_3_G1_MINI_ALU_nx403, L1_0_L2_3_G1_MINI_ALU_nx405, 
         L1_0_L2_3_G1_MINI_ALU_nx409, L1_0_L2_3_G1_MINI_ALU_nx411, 
         L1_0_L2_3_G1_MINI_ALU_nx413, L1_0_L2_3_G1_MINI_ALU_nx415, 
         L1_0_L2_3_G1_MINI_ALU_nx419, L1_0_L2_3_G1_MINI_ALU_nx421, 
         L1_0_L2_3_G1_MINI_ALU_nx423, L1_0_L2_3_G1_MINI_ALU_nx425, 
         L1_0_L2_3_G1_MINI_ALU_nx429, L1_0_L2_3_G1_MINI_ALU_nx431, 
         L1_0_L2_3_G1_MINI_ALU_nx433, L1_0_L2_3_G1_MINI_ALU_nx435, 
         L1_0_L2_3_G1_MINI_ALU_nx439, L1_0_L2_3_G1_MINI_ALU_nx441, 
         L1_0_L2_3_G1_MINI_ALU_nx443, L1_0_L2_3_G1_MINI_ALU_nx445, 
         L1_0_L2_3_G1_MINI_ALU_nx449, L1_0_L2_3_G1_MINI_ALU_nx451, 
         L1_0_L2_3_G1_MINI_ALU_nx453, L1_0_L2_3_G1_MINI_ALU_nx455, 
         L1_0_L2_3_G1_MINI_ALU_nx461, L1_0_L2_3_G1_MINI_ALU_nx463, 
         L1_0_L2_3_G1_MINI_ALU_nx467, L1_0_L2_3_G1_MINI_ALU_nx469, 
         L1_0_L2_3_G1_MINI_ALU_nx471, L1_0_L2_3_G1_MINI_ALU_nx475, 
         L1_0_L2_3_G1_MINI_ALU_nx477, L1_0_L2_3_G1_MINI_ALU_nx479, 
         L1_0_L2_3_G1_MINI_ALU_nx483, L1_0_L2_3_G1_MINI_ALU_nx485, 
         L1_0_L2_3_G1_MINI_ALU_nx487, L1_0_L2_3_G1_MINI_ALU_nx491, 
         L1_0_L2_3_G1_MINI_ALU_nx493, L1_0_L2_3_G1_MINI_ALU_nx495, 
         L1_0_L2_3_G1_MINI_ALU_nx499, L1_0_L2_3_G1_MINI_ALU_nx501, 
         L1_0_L2_3_G1_MINI_ALU_nx503, L1_0_L2_3_G1_MINI_ALU_nx507, 
         L1_0_L2_3_G1_MINI_ALU_nx509, L1_0_L2_3_G1_MINI_ALU_nx511, 
         L1_0_L2_3_G1_MINI_ALU_nx515, L1_0_L2_3_G1_MINI_ALU_nx517, 
         L1_0_L2_3_G1_MINI_ALU_nx529, L1_0_L2_3_G1_MINI_ALU_nx531, 
         L1_0_L2_3_G1_MINI_ALU_nx534, L1_0_L2_3_G1_MINI_ALU_nx537, 
         L1_0_L2_3_G1_MINI_ALU_nx540, L1_0_L2_3_G1_MINI_ALU_nx544, 
         L1_0_L2_3_G1_MINI_ALU_nx547, L1_0_L2_3_G1_MINI_ALU_nx551, 
         L1_0_L2_3_G1_MINI_ALU_nx554, L1_0_L2_3_G1_MINI_ALU_nx558, 
         L1_0_L2_3_G1_MINI_ALU_nx561, L1_0_L2_3_G1_MINI_ALU_nx565, 
         L1_0_L2_3_G1_MINI_ALU_nx568, 
         L1_0_L2_3_G1_MINI_ALU_WindowCellShiftedLeft_16, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_16, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_15, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_14, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_13, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_12, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_11, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_10, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_16, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_15, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_14, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_13, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_12, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_11, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_10, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_9, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_8, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_7, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_6, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_5, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_4, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_3, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_2, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_1, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_0, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_16, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_15, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_14, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_13, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_12, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_11, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_10, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_9, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_8, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_7, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_6, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_5, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_4, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_3, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_2, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_1, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_0, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_16, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_15, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_14, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_13, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_12, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_11, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_10, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_9, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_8, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_7, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_6, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_5, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_4, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_3, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_2, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_1, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_0, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx4, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx8, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx12, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx16, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx20, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx24, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx80, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx328, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx384, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642, 
         L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644, 
         L1_0_L2_4_G1_MINI_ALU_AddPToBoothOperand, 
         L1_0_L2_4_G1_MINI_ALU_BoothOperand_16, 
         L1_0_L2_4_G1_MINI_ALU_BoothOperand_15, 
         L1_0_L2_4_G1_MINI_ALU_BoothOperand_14, 
         L1_0_L2_4_G1_MINI_ALU_BoothOperand_13, 
         L1_0_L2_4_G1_MINI_ALU_BoothOperand_12, 
         L1_0_L2_4_G1_MINI_ALU_BoothOperand_11, 
         L1_0_L2_4_G1_MINI_ALU_BoothOperand_10, 
         L1_0_L2_4_G1_MINI_ALU_BoothOperand_9, 
         L1_0_L2_4_G1_MINI_ALU_BoothOperand_8, 
         L1_0_L2_4_G1_MINI_ALU_BoothOperand_7, 
         L1_0_L2_4_G1_MINI_ALU_BoothOperand_6, 
         L1_0_L2_4_G1_MINI_ALU_BoothOperand_5, 
         L1_0_L2_4_G1_MINI_ALU_BoothOperand_4, 
         L1_0_L2_4_G1_MINI_ALU_BoothOperand_3, 
         L1_0_L2_4_G1_MINI_ALU_BoothOperand_2, 
         L1_0_L2_4_G1_MINI_ALU_BoothOperand_1, 
         L1_0_L2_4_G1_MINI_ALU_BoothOperand_0, 
         L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_16, 
         L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_15, 
         L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_14, 
         L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_13, 
         L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_12, 
         L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_11, 
         L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_10, 
         L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_9, 
         L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_8, 
         L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_7, 
         L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_6, 
         L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_5, 
         L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_4, 
         L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_3, 
         L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_2, 
         L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_1, 
         L1_0_L2_4_G1_MINI_ALU_BoothP_16, L1_0_L2_4_G1_MINI_ALU_BoothP_15, 
         L1_0_L2_4_G1_MINI_ALU_BoothP_14, L1_0_L2_4_G1_MINI_ALU_BoothP_13, 
         L1_0_L2_4_G1_MINI_ALU_BoothP_12, L1_0_L2_4_G1_MINI_ALU_BoothP_11, 
         L1_0_L2_4_G1_MINI_ALU_BoothP_10, L1_0_L2_4_G1_MINI_ALU_BoothP_9, 
         L1_0_L2_4_G1_MINI_ALU_BoothP_8, L1_0_L2_4_G1_MINI_ALU_BoothP_7, 
         L1_0_L2_4_G1_MINI_ALU_BoothP_6, L1_0_L2_4_G1_MINI_ALU_BoothP_5, 
         L1_0_L2_4_G1_MINI_ALU_BoothP_4, L1_0_L2_4_G1_MINI_ALU_BoothP_3, 
         L1_0_L2_4_G1_MINI_ALU_BoothP_2, L1_0_L2_4_G1_MINI_ALU_BoothP_1, 
         L1_0_L2_4_G1_MINI_ALU_BoothP_0, L1_0_L2_4_G1_MINI_ALU_nx0, 
         L1_0_L2_4_G1_MINI_ALU_nx6, L1_0_L2_4_G1_MINI_ALU_nx12, 
         L1_0_L2_4_G1_MINI_ALU_nx18, L1_0_L2_4_G1_MINI_ALU_nx24, 
         L1_0_L2_4_G1_MINI_ALU_nx30, L1_0_L2_4_G1_MINI_ALU_nx40, 
         L1_0_L2_4_G1_MINI_ALU_nx44, L1_0_L2_4_G1_MINI_ALU_nx48, 
         L1_0_L2_4_G1_MINI_ALU_nx52, L1_0_L2_4_G1_MINI_ALU_nx56, 
         L1_0_L2_4_G1_MINI_ALU_nx62, L1_0_L2_4_G1_MINI_ALU_nx154, 
         L1_0_L2_4_G1_MINI_ALU_nx316, L1_0_L2_4_G1_MINI_ALU_nx336, 
         L1_0_L2_4_G1_MINI_ALU_nx356, L1_0_L2_4_G1_MINI_ALU_nx376, 
         L1_0_L2_4_G1_MINI_ALU_nx396, L1_0_L2_4_G1_MINI_ALU_nx416, 
         L1_0_L2_4_G1_MINI_ALU_nx436, L1_0_L2_4_G1_MINI_ALU_nx454, 
         L1_0_L2_4_G1_MINI_ALU_nx456, L1_0_L2_4_G1_MINI_ALU_nx379, 
         L1_0_L2_4_G1_MINI_ALU_nx381, L1_0_L2_4_G1_MINI_ALU_nx383, 
         L1_0_L2_4_G1_MINI_ALU_nx387, L1_0_L2_4_G1_MINI_ALU_nx389, 
         L1_0_L2_4_G1_MINI_ALU_nx391, L1_0_L2_4_G1_MINI_ALU_nx395, 
         L1_0_L2_4_G1_MINI_ALU_nx399, L1_0_L2_4_G1_MINI_ALU_nx401, 
         L1_0_L2_4_G1_MINI_ALU_nx403, L1_0_L2_4_G1_MINI_ALU_nx405, 
         L1_0_L2_4_G1_MINI_ALU_nx409, L1_0_L2_4_G1_MINI_ALU_nx411, 
         L1_0_L2_4_G1_MINI_ALU_nx413, L1_0_L2_4_G1_MINI_ALU_nx415, 
         L1_0_L2_4_G1_MINI_ALU_nx419, L1_0_L2_4_G1_MINI_ALU_nx421, 
         L1_0_L2_4_G1_MINI_ALU_nx423, L1_0_L2_4_G1_MINI_ALU_nx425, 
         L1_0_L2_4_G1_MINI_ALU_nx429, L1_0_L2_4_G1_MINI_ALU_nx431, 
         L1_0_L2_4_G1_MINI_ALU_nx433, L1_0_L2_4_G1_MINI_ALU_nx435, 
         L1_0_L2_4_G1_MINI_ALU_nx439, L1_0_L2_4_G1_MINI_ALU_nx441, 
         L1_0_L2_4_G1_MINI_ALU_nx443, L1_0_L2_4_G1_MINI_ALU_nx445, 
         L1_0_L2_4_G1_MINI_ALU_nx449, L1_0_L2_4_G1_MINI_ALU_nx451, 
         L1_0_L2_4_G1_MINI_ALU_nx453, L1_0_L2_4_G1_MINI_ALU_nx455, 
         L1_0_L2_4_G1_MINI_ALU_nx461, L1_0_L2_4_G1_MINI_ALU_nx463, 
         L1_0_L2_4_G1_MINI_ALU_nx467, L1_0_L2_4_G1_MINI_ALU_nx469, 
         L1_0_L2_4_G1_MINI_ALU_nx471, L1_0_L2_4_G1_MINI_ALU_nx475, 
         L1_0_L2_4_G1_MINI_ALU_nx477, L1_0_L2_4_G1_MINI_ALU_nx479, 
         L1_0_L2_4_G1_MINI_ALU_nx483, L1_0_L2_4_G1_MINI_ALU_nx485, 
         L1_0_L2_4_G1_MINI_ALU_nx487, L1_0_L2_4_G1_MINI_ALU_nx491, 
         L1_0_L2_4_G1_MINI_ALU_nx493, L1_0_L2_4_G1_MINI_ALU_nx495, 
         L1_0_L2_4_G1_MINI_ALU_nx499, L1_0_L2_4_G1_MINI_ALU_nx501, 
         L1_0_L2_4_G1_MINI_ALU_nx503, L1_0_L2_4_G1_MINI_ALU_nx507, 
         L1_0_L2_4_G1_MINI_ALU_nx509, L1_0_L2_4_G1_MINI_ALU_nx511, 
         L1_0_L2_4_G1_MINI_ALU_nx515, L1_0_L2_4_G1_MINI_ALU_nx517, 
         L1_0_L2_4_G1_MINI_ALU_nx529, L1_0_L2_4_G1_MINI_ALU_nx531, 
         L1_0_L2_4_G1_MINI_ALU_nx534, L1_0_L2_4_G1_MINI_ALU_nx537, 
         L1_0_L2_4_G1_MINI_ALU_nx540, L1_0_L2_4_G1_MINI_ALU_nx544, 
         L1_0_L2_4_G1_MINI_ALU_nx547, L1_0_L2_4_G1_MINI_ALU_nx551, 
         L1_0_L2_4_G1_MINI_ALU_nx554, L1_0_L2_4_G1_MINI_ALU_nx558, 
         L1_0_L2_4_G1_MINI_ALU_nx561, L1_0_L2_4_G1_MINI_ALU_nx565, 
         L1_0_L2_4_G1_MINI_ALU_nx568, 
         L1_0_L2_4_G1_MINI_ALU_WindowCellShiftedLeft_16, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_16, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_15, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_14, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_13, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_12, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_11, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_10, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_16, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_15, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_14, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_13, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_12, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_11, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_10, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_9, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_8, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_7, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_6, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_5, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_4, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_3, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_2, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_1, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_0, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_16, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_15, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_14, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_13, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_12, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_11, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_10, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_9, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_8, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_7, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_6, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_5, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_4, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_3, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_2, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_1, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_0, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_16, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_15, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_14, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_13, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_12, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_11, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_10, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_9, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_8, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_7, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_6, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_5, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_4, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_3, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_2, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_1, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_0, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx4, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx8, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx12, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx16, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx20, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx24, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx80, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx328, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx384, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642, 
         L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644, 
         L1_1_L2_0_G1_MINI_ALU_AddPToBoothOperand, 
         L1_1_L2_0_G1_MINI_ALU_BoothOperand_16, 
         L1_1_L2_0_G1_MINI_ALU_BoothOperand_15, 
         L1_1_L2_0_G1_MINI_ALU_BoothOperand_14, 
         L1_1_L2_0_G1_MINI_ALU_BoothOperand_13, 
         L1_1_L2_0_G1_MINI_ALU_BoothOperand_12, 
         L1_1_L2_0_G1_MINI_ALU_BoothOperand_11, 
         L1_1_L2_0_G1_MINI_ALU_BoothOperand_10, 
         L1_1_L2_0_G1_MINI_ALU_BoothOperand_9, 
         L1_1_L2_0_G1_MINI_ALU_BoothOperand_8, 
         L1_1_L2_0_G1_MINI_ALU_BoothOperand_7, 
         L1_1_L2_0_G1_MINI_ALU_BoothOperand_6, 
         L1_1_L2_0_G1_MINI_ALU_BoothOperand_5, 
         L1_1_L2_0_G1_MINI_ALU_BoothOperand_4, 
         L1_1_L2_0_G1_MINI_ALU_BoothOperand_3, 
         L1_1_L2_0_G1_MINI_ALU_BoothOperand_2, 
         L1_1_L2_0_G1_MINI_ALU_BoothOperand_1, 
         L1_1_L2_0_G1_MINI_ALU_BoothOperand_0, 
         L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_16, 
         L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_15, 
         L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_14, 
         L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_13, 
         L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_12, 
         L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_11, 
         L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_10, 
         L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_9, 
         L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_8, 
         L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_7, 
         L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_6, 
         L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_5, 
         L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_4, 
         L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_3, 
         L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_2, 
         L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_1, 
         L1_1_L2_0_G1_MINI_ALU_BoothP_16, L1_1_L2_0_G1_MINI_ALU_BoothP_15, 
         L1_1_L2_0_G1_MINI_ALU_BoothP_14, L1_1_L2_0_G1_MINI_ALU_BoothP_13, 
         L1_1_L2_0_G1_MINI_ALU_BoothP_12, L1_1_L2_0_G1_MINI_ALU_BoothP_11, 
         L1_1_L2_0_G1_MINI_ALU_BoothP_10, L1_1_L2_0_G1_MINI_ALU_BoothP_9, 
         L1_1_L2_0_G1_MINI_ALU_BoothP_8, L1_1_L2_0_G1_MINI_ALU_BoothP_7, 
         L1_1_L2_0_G1_MINI_ALU_BoothP_6, L1_1_L2_0_G1_MINI_ALU_BoothP_5, 
         L1_1_L2_0_G1_MINI_ALU_BoothP_4, L1_1_L2_0_G1_MINI_ALU_BoothP_3, 
         L1_1_L2_0_G1_MINI_ALU_BoothP_2, L1_1_L2_0_G1_MINI_ALU_BoothP_1, 
         L1_1_L2_0_G1_MINI_ALU_BoothP_0, L1_1_L2_0_G1_MINI_ALU_nx0, 
         L1_1_L2_0_G1_MINI_ALU_nx6, L1_1_L2_0_G1_MINI_ALU_nx12, 
         L1_1_L2_0_G1_MINI_ALU_nx18, L1_1_L2_0_G1_MINI_ALU_nx24, 
         L1_1_L2_0_G1_MINI_ALU_nx30, L1_1_L2_0_G1_MINI_ALU_nx40, 
         L1_1_L2_0_G1_MINI_ALU_nx44, L1_1_L2_0_G1_MINI_ALU_nx48, 
         L1_1_L2_0_G1_MINI_ALU_nx52, L1_1_L2_0_G1_MINI_ALU_nx56, 
         L1_1_L2_0_G1_MINI_ALU_nx62, L1_1_L2_0_G1_MINI_ALU_nx154, 
         L1_1_L2_0_G1_MINI_ALU_nx316, L1_1_L2_0_G1_MINI_ALU_nx336, 
         L1_1_L2_0_G1_MINI_ALU_nx356, L1_1_L2_0_G1_MINI_ALU_nx376, 
         L1_1_L2_0_G1_MINI_ALU_nx396, L1_1_L2_0_G1_MINI_ALU_nx416, 
         L1_1_L2_0_G1_MINI_ALU_nx436, L1_1_L2_0_G1_MINI_ALU_nx454, 
         L1_1_L2_0_G1_MINI_ALU_nx456, L1_1_L2_0_G1_MINI_ALU_nx379, 
         L1_1_L2_0_G1_MINI_ALU_nx381, L1_1_L2_0_G1_MINI_ALU_nx383, 
         L1_1_L2_0_G1_MINI_ALU_nx387, L1_1_L2_0_G1_MINI_ALU_nx389, 
         L1_1_L2_0_G1_MINI_ALU_nx391, L1_1_L2_0_G1_MINI_ALU_nx395, 
         L1_1_L2_0_G1_MINI_ALU_nx399, L1_1_L2_0_G1_MINI_ALU_nx401, 
         L1_1_L2_0_G1_MINI_ALU_nx403, L1_1_L2_0_G1_MINI_ALU_nx405, 
         L1_1_L2_0_G1_MINI_ALU_nx409, L1_1_L2_0_G1_MINI_ALU_nx411, 
         L1_1_L2_0_G1_MINI_ALU_nx413, L1_1_L2_0_G1_MINI_ALU_nx415, 
         L1_1_L2_0_G1_MINI_ALU_nx419, L1_1_L2_0_G1_MINI_ALU_nx421, 
         L1_1_L2_0_G1_MINI_ALU_nx423, L1_1_L2_0_G1_MINI_ALU_nx425, 
         L1_1_L2_0_G1_MINI_ALU_nx429, L1_1_L2_0_G1_MINI_ALU_nx431, 
         L1_1_L2_0_G1_MINI_ALU_nx433, L1_1_L2_0_G1_MINI_ALU_nx435, 
         L1_1_L2_0_G1_MINI_ALU_nx439, L1_1_L2_0_G1_MINI_ALU_nx441, 
         L1_1_L2_0_G1_MINI_ALU_nx443, L1_1_L2_0_G1_MINI_ALU_nx445, 
         L1_1_L2_0_G1_MINI_ALU_nx449, L1_1_L2_0_G1_MINI_ALU_nx451, 
         L1_1_L2_0_G1_MINI_ALU_nx453, L1_1_L2_0_G1_MINI_ALU_nx455, 
         L1_1_L2_0_G1_MINI_ALU_nx461, L1_1_L2_0_G1_MINI_ALU_nx463, 
         L1_1_L2_0_G1_MINI_ALU_nx467, L1_1_L2_0_G1_MINI_ALU_nx469, 
         L1_1_L2_0_G1_MINI_ALU_nx471, L1_1_L2_0_G1_MINI_ALU_nx475, 
         L1_1_L2_0_G1_MINI_ALU_nx477, L1_1_L2_0_G1_MINI_ALU_nx479, 
         L1_1_L2_0_G1_MINI_ALU_nx483, L1_1_L2_0_G1_MINI_ALU_nx485, 
         L1_1_L2_0_G1_MINI_ALU_nx487, L1_1_L2_0_G1_MINI_ALU_nx491, 
         L1_1_L2_0_G1_MINI_ALU_nx493, L1_1_L2_0_G1_MINI_ALU_nx495, 
         L1_1_L2_0_G1_MINI_ALU_nx499, L1_1_L2_0_G1_MINI_ALU_nx501, 
         L1_1_L2_0_G1_MINI_ALU_nx503, L1_1_L2_0_G1_MINI_ALU_nx507, 
         L1_1_L2_0_G1_MINI_ALU_nx509, L1_1_L2_0_G1_MINI_ALU_nx511, 
         L1_1_L2_0_G1_MINI_ALU_nx515, L1_1_L2_0_G1_MINI_ALU_nx517, 
         L1_1_L2_0_G1_MINI_ALU_nx529, L1_1_L2_0_G1_MINI_ALU_nx531, 
         L1_1_L2_0_G1_MINI_ALU_nx534, L1_1_L2_0_G1_MINI_ALU_nx537, 
         L1_1_L2_0_G1_MINI_ALU_nx540, L1_1_L2_0_G1_MINI_ALU_nx544, 
         L1_1_L2_0_G1_MINI_ALU_nx547, L1_1_L2_0_G1_MINI_ALU_nx551, 
         L1_1_L2_0_G1_MINI_ALU_nx554, L1_1_L2_0_G1_MINI_ALU_nx558, 
         L1_1_L2_0_G1_MINI_ALU_nx561, L1_1_L2_0_G1_MINI_ALU_nx565, 
         L1_1_L2_0_G1_MINI_ALU_nx568, 
         L1_1_L2_0_G1_MINI_ALU_WindowCellShiftedLeft_16, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_16, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_15, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_14, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_13, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_12, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_11, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_10, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_16, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_15, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_14, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_13, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_12, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_11, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_10, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_9, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_8, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_7, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_6, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_5, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_4, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_3, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_2, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_1, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_0, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_16, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_15, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_14, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_13, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_12, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_11, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_10, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_9, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_8, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_7, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_6, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_5, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_4, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_3, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_2, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_1, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_0, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_16, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_15, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_14, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_13, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_12, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_11, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_10, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_9, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_8, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_7, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_6, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_5, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_4, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_3, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_2, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_1, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_0, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx4, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx8, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx12, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx16, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx20, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx24, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx80, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx328, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx384, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642, 
         L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644, 
         L1_1_L2_1_G1_MINI_ALU_AddPToBoothOperand, 
         L1_1_L2_1_G1_MINI_ALU_BoothOperand_16, 
         L1_1_L2_1_G1_MINI_ALU_BoothOperand_15, 
         L1_1_L2_1_G1_MINI_ALU_BoothOperand_14, 
         L1_1_L2_1_G1_MINI_ALU_BoothOperand_13, 
         L1_1_L2_1_G1_MINI_ALU_BoothOperand_12, 
         L1_1_L2_1_G1_MINI_ALU_BoothOperand_11, 
         L1_1_L2_1_G1_MINI_ALU_BoothOperand_10, 
         L1_1_L2_1_G1_MINI_ALU_BoothOperand_9, 
         L1_1_L2_1_G1_MINI_ALU_BoothOperand_8, 
         L1_1_L2_1_G1_MINI_ALU_BoothOperand_7, 
         L1_1_L2_1_G1_MINI_ALU_BoothOperand_6, 
         L1_1_L2_1_G1_MINI_ALU_BoothOperand_5, 
         L1_1_L2_1_G1_MINI_ALU_BoothOperand_4, 
         L1_1_L2_1_G1_MINI_ALU_BoothOperand_3, 
         L1_1_L2_1_G1_MINI_ALU_BoothOperand_2, 
         L1_1_L2_1_G1_MINI_ALU_BoothOperand_1, 
         L1_1_L2_1_G1_MINI_ALU_BoothOperand_0, 
         L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_16, 
         L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_15, 
         L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_14, 
         L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_13, 
         L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_12, 
         L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_11, 
         L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_10, 
         L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_9, 
         L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_8, 
         L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_7, 
         L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_6, 
         L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_5, 
         L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_4, 
         L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_3, 
         L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_2, 
         L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_1, 
         L1_1_L2_1_G1_MINI_ALU_BoothP_16, L1_1_L2_1_G1_MINI_ALU_BoothP_15, 
         L1_1_L2_1_G1_MINI_ALU_BoothP_14, L1_1_L2_1_G1_MINI_ALU_BoothP_13, 
         L1_1_L2_1_G1_MINI_ALU_BoothP_12, L1_1_L2_1_G1_MINI_ALU_BoothP_11, 
         L1_1_L2_1_G1_MINI_ALU_BoothP_10, L1_1_L2_1_G1_MINI_ALU_BoothP_9, 
         L1_1_L2_1_G1_MINI_ALU_BoothP_8, L1_1_L2_1_G1_MINI_ALU_BoothP_7, 
         L1_1_L2_1_G1_MINI_ALU_BoothP_6, L1_1_L2_1_G1_MINI_ALU_BoothP_5, 
         L1_1_L2_1_G1_MINI_ALU_BoothP_4, L1_1_L2_1_G1_MINI_ALU_BoothP_3, 
         L1_1_L2_1_G1_MINI_ALU_BoothP_2, L1_1_L2_1_G1_MINI_ALU_BoothP_1, 
         L1_1_L2_1_G1_MINI_ALU_BoothP_0, L1_1_L2_1_G1_MINI_ALU_nx0, 
         L1_1_L2_1_G1_MINI_ALU_nx6, L1_1_L2_1_G1_MINI_ALU_nx12, 
         L1_1_L2_1_G1_MINI_ALU_nx18, L1_1_L2_1_G1_MINI_ALU_nx24, 
         L1_1_L2_1_G1_MINI_ALU_nx30, L1_1_L2_1_G1_MINI_ALU_nx40, 
         L1_1_L2_1_G1_MINI_ALU_nx44, L1_1_L2_1_G1_MINI_ALU_nx48, 
         L1_1_L2_1_G1_MINI_ALU_nx52, L1_1_L2_1_G1_MINI_ALU_nx56, 
         L1_1_L2_1_G1_MINI_ALU_nx62, L1_1_L2_1_G1_MINI_ALU_nx154, 
         L1_1_L2_1_G1_MINI_ALU_nx316, L1_1_L2_1_G1_MINI_ALU_nx336, 
         L1_1_L2_1_G1_MINI_ALU_nx356, L1_1_L2_1_G1_MINI_ALU_nx376, 
         L1_1_L2_1_G1_MINI_ALU_nx396, L1_1_L2_1_G1_MINI_ALU_nx416, 
         L1_1_L2_1_G1_MINI_ALU_nx436, L1_1_L2_1_G1_MINI_ALU_nx454, 
         L1_1_L2_1_G1_MINI_ALU_nx456, L1_1_L2_1_G1_MINI_ALU_nx379, 
         L1_1_L2_1_G1_MINI_ALU_nx381, L1_1_L2_1_G1_MINI_ALU_nx383, 
         L1_1_L2_1_G1_MINI_ALU_nx387, L1_1_L2_1_G1_MINI_ALU_nx389, 
         L1_1_L2_1_G1_MINI_ALU_nx391, L1_1_L2_1_G1_MINI_ALU_nx395, 
         L1_1_L2_1_G1_MINI_ALU_nx399, L1_1_L2_1_G1_MINI_ALU_nx401, 
         L1_1_L2_1_G1_MINI_ALU_nx403, L1_1_L2_1_G1_MINI_ALU_nx405, 
         L1_1_L2_1_G1_MINI_ALU_nx409, L1_1_L2_1_G1_MINI_ALU_nx411, 
         L1_1_L2_1_G1_MINI_ALU_nx413, L1_1_L2_1_G1_MINI_ALU_nx415, 
         L1_1_L2_1_G1_MINI_ALU_nx419, L1_1_L2_1_G1_MINI_ALU_nx421, 
         L1_1_L2_1_G1_MINI_ALU_nx423, L1_1_L2_1_G1_MINI_ALU_nx425, 
         L1_1_L2_1_G1_MINI_ALU_nx429, L1_1_L2_1_G1_MINI_ALU_nx431, 
         L1_1_L2_1_G1_MINI_ALU_nx433, L1_1_L2_1_G1_MINI_ALU_nx435, 
         L1_1_L2_1_G1_MINI_ALU_nx439, L1_1_L2_1_G1_MINI_ALU_nx441, 
         L1_1_L2_1_G1_MINI_ALU_nx443, L1_1_L2_1_G1_MINI_ALU_nx445, 
         L1_1_L2_1_G1_MINI_ALU_nx449, L1_1_L2_1_G1_MINI_ALU_nx451, 
         L1_1_L2_1_G1_MINI_ALU_nx453, L1_1_L2_1_G1_MINI_ALU_nx455, 
         L1_1_L2_1_G1_MINI_ALU_nx461, L1_1_L2_1_G1_MINI_ALU_nx463, 
         L1_1_L2_1_G1_MINI_ALU_nx467, L1_1_L2_1_G1_MINI_ALU_nx469, 
         L1_1_L2_1_G1_MINI_ALU_nx471, L1_1_L2_1_G1_MINI_ALU_nx475, 
         L1_1_L2_1_G1_MINI_ALU_nx477, L1_1_L2_1_G1_MINI_ALU_nx479, 
         L1_1_L2_1_G1_MINI_ALU_nx483, L1_1_L2_1_G1_MINI_ALU_nx485, 
         L1_1_L2_1_G1_MINI_ALU_nx487, L1_1_L2_1_G1_MINI_ALU_nx491, 
         L1_1_L2_1_G1_MINI_ALU_nx493, L1_1_L2_1_G1_MINI_ALU_nx495, 
         L1_1_L2_1_G1_MINI_ALU_nx499, L1_1_L2_1_G1_MINI_ALU_nx501, 
         L1_1_L2_1_G1_MINI_ALU_nx503, L1_1_L2_1_G1_MINI_ALU_nx507, 
         L1_1_L2_1_G1_MINI_ALU_nx509, L1_1_L2_1_G1_MINI_ALU_nx511, 
         L1_1_L2_1_G1_MINI_ALU_nx515, L1_1_L2_1_G1_MINI_ALU_nx517, 
         L1_1_L2_1_G1_MINI_ALU_nx529, L1_1_L2_1_G1_MINI_ALU_nx531, 
         L1_1_L2_1_G1_MINI_ALU_nx534, L1_1_L2_1_G1_MINI_ALU_nx537, 
         L1_1_L2_1_G1_MINI_ALU_nx540, L1_1_L2_1_G1_MINI_ALU_nx544, 
         L1_1_L2_1_G1_MINI_ALU_nx547, L1_1_L2_1_G1_MINI_ALU_nx551, 
         L1_1_L2_1_G1_MINI_ALU_nx554, L1_1_L2_1_G1_MINI_ALU_nx558, 
         L1_1_L2_1_G1_MINI_ALU_nx561, L1_1_L2_1_G1_MINI_ALU_nx565, 
         L1_1_L2_1_G1_MINI_ALU_nx568, 
         L1_1_L2_1_G1_MINI_ALU_WindowCellShiftedLeft_16, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_16, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_15, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_14, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_13, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_12, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_11, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_10, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_16, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_15, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_14, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_13, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_12, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_11, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_10, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_9, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_8, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_7, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_6, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_5, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_4, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_3, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_2, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_1, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_0, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_16, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_15, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_14, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_13, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_12, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_11, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_10, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_9, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_8, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_7, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_6, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_5, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_4, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_3, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_2, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_1, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_0, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_16, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_15, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_14, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_13, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_12, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_11, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_10, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_9, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_8, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_7, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_6, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_5, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_4, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_3, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_2, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_1, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_0, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx4, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx8, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx12, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx16, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx20, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx24, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx80, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx328, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx384, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642, 
         L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644, 
         L1_1_L2_2_G1_MINI_ALU_AddPToBoothOperand, 
         L1_1_L2_2_G1_MINI_ALU_BoothOperand_16, 
         L1_1_L2_2_G1_MINI_ALU_BoothOperand_15, 
         L1_1_L2_2_G1_MINI_ALU_BoothOperand_14, 
         L1_1_L2_2_G1_MINI_ALU_BoothOperand_13, 
         L1_1_L2_2_G1_MINI_ALU_BoothOperand_12, 
         L1_1_L2_2_G1_MINI_ALU_BoothOperand_11, 
         L1_1_L2_2_G1_MINI_ALU_BoothOperand_10, 
         L1_1_L2_2_G1_MINI_ALU_BoothOperand_9, 
         L1_1_L2_2_G1_MINI_ALU_BoothOperand_8, 
         L1_1_L2_2_G1_MINI_ALU_BoothOperand_7, 
         L1_1_L2_2_G1_MINI_ALU_BoothOperand_6, 
         L1_1_L2_2_G1_MINI_ALU_BoothOperand_5, 
         L1_1_L2_2_G1_MINI_ALU_BoothOperand_4, 
         L1_1_L2_2_G1_MINI_ALU_BoothOperand_3, 
         L1_1_L2_2_G1_MINI_ALU_BoothOperand_2, 
         L1_1_L2_2_G1_MINI_ALU_BoothOperand_1, 
         L1_1_L2_2_G1_MINI_ALU_BoothOperand_0, 
         L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_16, 
         L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_15, 
         L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_14, 
         L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_13, 
         L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_12, 
         L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_11, 
         L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_10, 
         L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_9, 
         L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_8, 
         L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_7, 
         L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_6, 
         L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_5, 
         L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_4, 
         L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_3, 
         L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_2, 
         L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_1, 
         L1_1_L2_2_G1_MINI_ALU_BoothP_16, L1_1_L2_2_G1_MINI_ALU_BoothP_15, 
         L1_1_L2_2_G1_MINI_ALU_BoothP_14, L1_1_L2_2_G1_MINI_ALU_BoothP_13, 
         L1_1_L2_2_G1_MINI_ALU_BoothP_12, L1_1_L2_2_G1_MINI_ALU_BoothP_11, 
         L1_1_L2_2_G1_MINI_ALU_BoothP_10, L1_1_L2_2_G1_MINI_ALU_BoothP_9, 
         L1_1_L2_2_G1_MINI_ALU_BoothP_8, L1_1_L2_2_G1_MINI_ALU_BoothP_7, 
         L1_1_L2_2_G1_MINI_ALU_BoothP_6, L1_1_L2_2_G1_MINI_ALU_BoothP_5, 
         L1_1_L2_2_G1_MINI_ALU_BoothP_4, L1_1_L2_2_G1_MINI_ALU_BoothP_3, 
         L1_1_L2_2_G1_MINI_ALU_BoothP_2, L1_1_L2_2_G1_MINI_ALU_BoothP_1, 
         L1_1_L2_2_G1_MINI_ALU_BoothP_0, L1_1_L2_2_G1_MINI_ALU_nx0, 
         L1_1_L2_2_G1_MINI_ALU_nx6, L1_1_L2_2_G1_MINI_ALU_nx12, 
         L1_1_L2_2_G1_MINI_ALU_nx18, L1_1_L2_2_G1_MINI_ALU_nx24, 
         L1_1_L2_2_G1_MINI_ALU_nx30, L1_1_L2_2_G1_MINI_ALU_nx40, 
         L1_1_L2_2_G1_MINI_ALU_nx44, L1_1_L2_2_G1_MINI_ALU_nx48, 
         L1_1_L2_2_G1_MINI_ALU_nx52, L1_1_L2_2_G1_MINI_ALU_nx56, 
         L1_1_L2_2_G1_MINI_ALU_nx62, L1_1_L2_2_G1_MINI_ALU_nx154, 
         L1_1_L2_2_G1_MINI_ALU_nx316, L1_1_L2_2_G1_MINI_ALU_nx336, 
         L1_1_L2_2_G1_MINI_ALU_nx356, L1_1_L2_2_G1_MINI_ALU_nx376, 
         L1_1_L2_2_G1_MINI_ALU_nx396, L1_1_L2_2_G1_MINI_ALU_nx416, 
         L1_1_L2_2_G1_MINI_ALU_nx436, L1_1_L2_2_G1_MINI_ALU_nx454, 
         L1_1_L2_2_G1_MINI_ALU_nx456, L1_1_L2_2_G1_MINI_ALU_nx379, 
         L1_1_L2_2_G1_MINI_ALU_nx381, L1_1_L2_2_G1_MINI_ALU_nx383, 
         L1_1_L2_2_G1_MINI_ALU_nx387, L1_1_L2_2_G1_MINI_ALU_nx389, 
         L1_1_L2_2_G1_MINI_ALU_nx391, L1_1_L2_2_G1_MINI_ALU_nx395, 
         L1_1_L2_2_G1_MINI_ALU_nx399, L1_1_L2_2_G1_MINI_ALU_nx401, 
         L1_1_L2_2_G1_MINI_ALU_nx403, L1_1_L2_2_G1_MINI_ALU_nx405, 
         L1_1_L2_2_G1_MINI_ALU_nx409, L1_1_L2_2_G1_MINI_ALU_nx411, 
         L1_1_L2_2_G1_MINI_ALU_nx413, L1_1_L2_2_G1_MINI_ALU_nx415, 
         L1_1_L2_2_G1_MINI_ALU_nx419, L1_1_L2_2_G1_MINI_ALU_nx421, 
         L1_1_L2_2_G1_MINI_ALU_nx423, L1_1_L2_2_G1_MINI_ALU_nx425, 
         L1_1_L2_2_G1_MINI_ALU_nx429, L1_1_L2_2_G1_MINI_ALU_nx431, 
         L1_1_L2_2_G1_MINI_ALU_nx433, L1_1_L2_2_G1_MINI_ALU_nx435, 
         L1_1_L2_2_G1_MINI_ALU_nx439, L1_1_L2_2_G1_MINI_ALU_nx441, 
         L1_1_L2_2_G1_MINI_ALU_nx443, L1_1_L2_2_G1_MINI_ALU_nx445, 
         L1_1_L2_2_G1_MINI_ALU_nx449, L1_1_L2_2_G1_MINI_ALU_nx451, 
         L1_1_L2_2_G1_MINI_ALU_nx453, L1_1_L2_2_G1_MINI_ALU_nx455, 
         L1_1_L2_2_G1_MINI_ALU_nx461, L1_1_L2_2_G1_MINI_ALU_nx463, 
         L1_1_L2_2_G1_MINI_ALU_nx467, L1_1_L2_2_G1_MINI_ALU_nx469, 
         L1_1_L2_2_G1_MINI_ALU_nx471, L1_1_L2_2_G1_MINI_ALU_nx475, 
         L1_1_L2_2_G1_MINI_ALU_nx477, L1_1_L2_2_G1_MINI_ALU_nx479, 
         L1_1_L2_2_G1_MINI_ALU_nx483, L1_1_L2_2_G1_MINI_ALU_nx485, 
         L1_1_L2_2_G1_MINI_ALU_nx487, L1_1_L2_2_G1_MINI_ALU_nx491, 
         L1_1_L2_2_G1_MINI_ALU_nx493, L1_1_L2_2_G1_MINI_ALU_nx495, 
         L1_1_L2_2_G1_MINI_ALU_nx499, L1_1_L2_2_G1_MINI_ALU_nx501, 
         L1_1_L2_2_G1_MINI_ALU_nx503, L1_1_L2_2_G1_MINI_ALU_nx507, 
         L1_1_L2_2_G1_MINI_ALU_nx509, L1_1_L2_2_G1_MINI_ALU_nx511, 
         L1_1_L2_2_G1_MINI_ALU_nx515, L1_1_L2_2_G1_MINI_ALU_nx517, 
         L1_1_L2_2_G1_MINI_ALU_nx529, L1_1_L2_2_G1_MINI_ALU_nx531, 
         L1_1_L2_2_G1_MINI_ALU_nx534, L1_1_L2_2_G1_MINI_ALU_nx537, 
         L1_1_L2_2_G1_MINI_ALU_nx540, L1_1_L2_2_G1_MINI_ALU_nx544, 
         L1_1_L2_2_G1_MINI_ALU_nx547, L1_1_L2_2_G1_MINI_ALU_nx551, 
         L1_1_L2_2_G1_MINI_ALU_nx554, L1_1_L2_2_G1_MINI_ALU_nx558, 
         L1_1_L2_2_G1_MINI_ALU_nx561, L1_1_L2_2_G1_MINI_ALU_nx565, 
         L1_1_L2_2_G1_MINI_ALU_nx568, 
         L1_1_L2_2_G1_MINI_ALU_WindowCellShiftedLeft_16, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_16, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_15, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_14, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_13, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_12, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_11, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_10, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_16, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_15, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_14, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_13, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_12, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_11, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_10, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_9, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_8, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_7, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_6, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_5, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_4, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_3, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_2, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_1, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_0, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_16, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_15, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_14, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_13, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_12, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_11, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_10, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_9, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_8, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_7, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_6, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_5, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_4, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_3, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_2, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_1, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_0, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_16, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_15, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_14, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_13, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_12, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_11, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_10, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_9, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_8, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_7, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_6, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_5, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_4, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_3, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_2, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_1, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_0, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx4, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx8, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx12, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx16, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx20, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx24, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx80, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx328, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx384, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642, 
         L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644, 
         L1_1_L2_3_G1_MINI_ALU_AddPToBoothOperand, 
         L1_1_L2_3_G1_MINI_ALU_BoothOperand_16, 
         L1_1_L2_3_G1_MINI_ALU_BoothOperand_15, 
         L1_1_L2_3_G1_MINI_ALU_BoothOperand_14, 
         L1_1_L2_3_G1_MINI_ALU_BoothOperand_13, 
         L1_1_L2_3_G1_MINI_ALU_BoothOperand_12, 
         L1_1_L2_3_G1_MINI_ALU_BoothOperand_11, 
         L1_1_L2_3_G1_MINI_ALU_BoothOperand_10, 
         L1_1_L2_3_G1_MINI_ALU_BoothOperand_9, 
         L1_1_L2_3_G1_MINI_ALU_BoothOperand_8, 
         L1_1_L2_3_G1_MINI_ALU_BoothOperand_7, 
         L1_1_L2_3_G1_MINI_ALU_BoothOperand_6, 
         L1_1_L2_3_G1_MINI_ALU_BoothOperand_5, 
         L1_1_L2_3_G1_MINI_ALU_BoothOperand_4, 
         L1_1_L2_3_G1_MINI_ALU_BoothOperand_3, 
         L1_1_L2_3_G1_MINI_ALU_BoothOperand_2, 
         L1_1_L2_3_G1_MINI_ALU_BoothOperand_1, 
         L1_1_L2_3_G1_MINI_ALU_BoothOperand_0, 
         L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_16, 
         L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_15, 
         L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_14, 
         L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_13, 
         L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_12, 
         L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_11, 
         L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_10, 
         L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_9, 
         L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_8, 
         L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_7, 
         L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_6, 
         L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_5, 
         L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_4, 
         L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_3, 
         L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_2, 
         L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_1, 
         L1_1_L2_3_G1_MINI_ALU_BoothP_16, L1_1_L2_3_G1_MINI_ALU_BoothP_15, 
         L1_1_L2_3_G1_MINI_ALU_BoothP_14, L1_1_L2_3_G1_MINI_ALU_BoothP_13, 
         L1_1_L2_3_G1_MINI_ALU_BoothP_12, L1_1_L2_3_G1_MINI_ALU_BoothP_11, 
         L1_1_L2_3_G1_MINI_ALU_BoothP_10, L1_1_L2_3_G1_MINI_ALU_BoothP_9, 
         L1_1_L2_3_G1_MINI_ALU_BoothP_8, L1_1_L2_3_G1_MINI_ALU_BoothP_7, 
         L1_1_L2_3_G1_MINI_ALU_BoothP_6, L1_1_L2_3_G1_MINI_ALU_BoothP_5, 
         L1_1_L2_3_G1_MINI_ALU_BoothP_4, L1_1_L2_3_G1_MINI_ALU_BoothP_3, 
         L1_1_L2_3_G1_MINI_ALU_BoothP_2, L1_1_L2_3_G1_MINI_ALU_BoothP_1, 
         L1_1_L2_3_G1_MINI_ALU_BoothP_0, L1_1_L2_3_G1_MINI_ALU_nx0, 
         L1_1_L2_3_G1_MINI_ALU_nx6, L1_1_L2_3_G1_MINI_ALU_nx12, 
         L1_1_L2_3_G1_MINI_ALU_nx18, L1_1_L2_3_G1_MINI_ALU_nx24, 
         L1_1_L2_3_G1_MINI_ALU_nx30, L1_1_L2_3_G1_MINI_ALU_nx40, 
         L1_1_L2_3_G1_MINI_ALU_nx44, L1_1_L2_3_G1_MINI_ALU_nx48, 
         L1_1_L2_3_G1_MINI_ALU_nx52, L1_1_L2_3_G1_MINI_ALU_nx56, 
         L1_1_L2_3_G1_MINI_ALU_nx62, L1_1_L2_3_G1_MINI_ALU_nx154, 
         L1_1_L2_3_G1_MINI_ALU_nx316, L1_1_L2_3_G1_MINI_ALU_nx336, 
         L1_1_L2_3_G1_MINI_ALU_nx356, L1_1_L2_3_G1_MINI_ALU_nx376, 
         L1_1_L2_3_G1_MINI_ALU_nx396, L1_1_L2_3_G1_MINI_ALU_nx416, 
         L1_1_L2_3_G1_MINI_ALU_nx436, L1_1_L2_3_G1_MINI_ALU_nx454, 
         L1_1_L2_3_G1_MINI_ALU_nx456, L1_1_L2_3_G1_MINI_ALU_nx379, 
         L1_1_L2_3_G1_MINI_ALU_nx381, L1_1_L2_3_G1_MINI_ALU_nx383, 
         L1_1_L2_3_G1_MINI_ALU_nx387, L1_1_L2_3_G1_MINI_ALU_nx389, 
         L1_1_L2_3_G1_MINI_ALU_nx391, L1_1_L2_3_G1_MINI_ALU_nx395, 
         L1_1_L2_3_G1_MINI_ALU_nx399, L1_1_L2_3_G1_MINI_ALU_nx401, 
         L1_1_L2_3_G1_MINI_ALU_nx403, L1_1_L2_3_G1_MINI_ALU_nx405, 
         L1_1_L2_3_G1_MINI_ALU_nx409, L1_1_L2_3_G1_MINI_ALU_nx411, 
         L1_1_L2_3_G1_MINI_ALU_nx413, L1_1_L2_3_G1_MINI_ALU_nx415, 
         L1_1_L2_3_G1_MINI_ALU_nx419, L1_1_L2_3_G1_MINI_ALU_nx421, 
         L1_1_L2_3_G1_MINI_ALU_nx423, L1_1_L2_3_G1_MINI_ALU_nx425, 
         L1_1_L2_3_G1_MINI_ALU_nx429, L1_1_L2_3_G1_MINI_ALU_nx431, 
         L1_1_L2_3_G1_MINI_ALU_nx433, L1_1_L2_3_G1_MINI_ALU_nx435, 
         L1_1_L2_3_G1_MINI_ALU_nx439, L1_1_L2_3_G1_MINI_ALU_nx441, 
         L1_1_L2_3_G1_MINI_ALU_nx443, L1_1_L2_3_G1_MINI_ALU_nx445, 
         L1_1_L2_3_G1_MINI_ALU_nx449, L1_1_L2_3_G1_MINI_ALU_nx451, 
         L1_1_L2_3_G1_MINI_ALU_nx453, L1_1_L2_3_G1_MINI_ALU_nx455, 
         L1_1_L2_3_G1_MINI_ALU_nx461, L1_1_L2_3_G1_MINI_ALU_nx463, 
         L1_1_L2_3_G1_MINI_ALU_nx467, L1_1_L2_3_G1_MINI_ALU_nx469, 
         L1_1_L2_3_G1_MINI_ALU_nx471, L1_1_L2_3_G1_MINI_ALU_nx475, 
         L1_1_L2_3_G1_MINI_ALU_nx477, L1_1_L2_3_G1_MINI_ALU_nx479, 
         L1_1_L2_3_G1_MINI_ALU_nx483, L1_1_L2_3_G1_MINI_ALU_nx485, 
         L1_1_L2_3_G1_MINI_ALU_nx487, L1_1_L2_3_G1_MINI_ALU_nx491, 
         L1_1_L2_3_G1_MINI_ALU_nx493, L1_1_L2_3_G1_MINI_ALU_nx495, 
         L1_1_L2_3_G1_MINI_ALU_nx499, L1_1_L2_3_G1_MINI_ALU_nx501, 
         L1_1_L2_3_G1_MINI_ALU_nx503, L1_1_L2_3_G1_MINI_ALU_nx507, 
         L1_1_L2_3_G1_MINI_ALU_nx509, L1_1_L2_3_G1_MINI_ALU_nx511, 
         L1_1_L2_3_G1_MINI_ALU_nx515, L1_1_L2_3_G1_MINI_ALU_nx517, 
         L1_1_L2_3_G1_MINI_ALU_nx529, L1_1_L2_3_G1_MINI_ALU_nx531, 
         L1_1_L2_3_G1_MINI_ALU_nx534, L1_1_L2_3_G1_MINI_ALU_nx537, 
         L1_1_L2_3_G1_MINI_ALU_nx540, L1_1_L2_3_G1_MINI_ALU_nx544, 
         L1_1_L2_3_G1_MINI_ALU_nx547, L1_1_L2_3_G1_MINI_ALU_nx551, 
         L1_1_L2_3_G1_MINI_ALU_nx554, L1_1_L2_3_G1_MINI_ALU_nx558, 
         L1_1_L2_3_G1_MINI_ALU_nx561, L1_1_L2_3_G1_MINI_ALU_nx565, 
         L1_1_L2_3_G1_MINI_ALU_nx568, 
         L1_1_L2_3_G1_MINI_ALU_WindowCellShiftedLeft_16, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_16, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_15, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_14, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_13, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_12, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_11, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_10, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_16, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_15, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_14, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_13, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_12, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_11, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_10, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_9, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_8, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_7, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_6, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_5, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_4, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_3, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_2, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_1, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_0, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_16, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_15, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_14, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_13, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_12, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_11, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_10, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_9, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_8, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_7, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_6, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_5, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_4, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_3, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_2, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_1, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_0, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_16, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_15, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_14, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_13, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_12, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_11, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_10, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_9, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_8, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_7, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_6, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_5, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_4, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_3, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_2, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_1, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_0, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx4, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx8, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx12, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx16, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx20, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx24, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx80, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx328, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx384, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642, 
         L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644, 
         L1_1_L2_4_G1_MINI_ALU_AddPToBoothOperand, 
         L1_1_L2_4_G1_MINI_ALU_BoothOperand_16, 
         L1_1_L2_4_G1_MINI_ALU_BoothOperand_15, 
         L1_1_L2_4_G1_MINI_ALU_BoothOperand_14, 
         L1_1_L2_4_G1_MINI_ALU_BoothOperand_13, 
         L1_1_L2_4_G1_MINI_ALU_BoothOperand_12, 
         L1_1_L2_4_G1_MINI_ALU_BoothOperand_11, 
         L1_1_L2_4_G1_MINI_ALU_BoothOperand_10, 
         L1_1_L2_4_G1_MINI_ALU_BoothOperand_9, 
         L1_1_L2_4_G1_MINI_ALU_BoothOperand_8, 
         L1_1_L2_4_G1_MINI_ALU_BoothOperand_7, 
         L1_1_L2_4_G1_MINI_ALU_BoothOperand_6, 
         L1_1_L2_4_G1_MINI_ALU_BoothOperand_5, 
         L1_1_L2_4_G1_MINI_ALU_BoothOperand_4, 
         L1_1_L2_4_G1_MINI_ALU_BoothOperand_3, 
         L1_1_L2_4_G1_MINI_ALU_BoothOperand_2, 
         L1_1_L2_4_G1_MINI_ALU_BoothOperand_1, 
         L1_1_L2_4_G1_MINI_ALU_BoothOperand_0, 
         L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_16, 
         L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_15, 
         L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_14, 
         L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_13, 
         L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_12, 
         L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_11, 
         L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_10, 
         L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_9, 
         L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_8, 
         L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_7, 
         L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_6, 
         L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_5, 
         L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_4, 
         L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_3, 
         L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_2, 
         L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_1, 
         L1_1_L2_4_G1_MINI_ALU_BoothP_16, L1_1_L2_4_G1_MINI_ALU_BoothP_15, 
         L1_1_L2_4_G1_MINI_ALU_BoothP_14, L1_1_L2_4_G1_MINI_ALU_BoothP_13, 
         L1_1_L2_4_G1_MINI_ALU_BoothP_12, L1_1_L2_4_G1_MINI_ALU_BoothP_11, 
         L1_1_L2_4_G1_MINI_ALU_BoothP_10, L1_1_L2_4_G1_MINI_ALU_BoothP_9, 
         L1_1_L2_4_G1_MINI_ALU_BoothP_8, L1_1_L2_4_G1_MINI_ALU_BoothP_7, 
         L1_1_L2_4_G1_MINI_ALU_BoothP_6, L1_1_L2_4_G1_MINI_ALU_BoothP_5, 
         L1_1_L2_4_G1_MINI_ALU_BoothP_4, L1_1_L2_4_G1_MINI_ALU_BoothP_3, 
         L1_1_L2_4_G1_MINI_ALU_BoothP_2, L1_1_L2_4_G1_MINI_ALU_BoothP_1, 
         L1_1_L2_4_G1_MINI_ALU_BoothP_0, L1_1_L2_4_G1_MINI_ALU_nx0, 
         L1_1_L2_4_G1_MINI_ALU_nx6, L1_1_L2_4_G1_MINI_ALU_nx12, 
         L1_1_L2_4_G1_MINI_ALU_nx18, L1_1_L2_4_G1_MINI_ALU_nx24, 
         L1_1_L2_4_G1_MINI_ALU_nx30, L1_1_L2_4_G1_MINI_ALU_nx40, 
         L1_1_L2_4_G1_MINI_ALU_nx44, L1_1_L2_4_G1_MINI_ALU_nx48, 
         L1_1_L2_4_G1_MINI_ALU_nx52, L1_1_L2_4_G1_MINI_ALU_nx56, 
         L1_1_L2_4_G1_MINI_ALU_nx62, L1_1_L2_4_G1_MINI_ALU_nx154, 
         L1_1_L2_4_G1_MINI_ALU_nx316, L1_1_L2_4_G1_MINI_ALU_nx336, 
         L1_1_L2_4_G1_MINI_ALU_nx356, L1_1_L2_4_G1_MINI_ALU_nx376, 
         L1_1_L2_4_G1_MINI_ALU_nx396, L1_1_L2_4_G1_MINI_ALU_nx416, 
         L1_1_L2_4_G1_MINI_ALU_nx436, L1_1_L2_4_G1_MINI_ALU_nx454, 
         L1_1_L2_4_G1_MINI_ALU_nx456, L1_1_L2_4_G1_MINI_ALU_nx379, 
         L1_1_L2_4_G1_MINI_ALU_nx381, L1_1_L2_4_G1_MINI_ALU_nx383, 
         L1_1_L2_4_G1_MINI_ALU_nx387, L1_1_L2_4_G1_MINI_ALU_nx389, 
         L1_1_L2_4_G1_MINI_ALU_nx391, L1_1_L2_4_G1_MINI_ALU_nx395, 
         L1_1_L2_4_G1_MINI_ALU_nx399, L1_1_L2_4_G1_MINI_ALU_nx401, 
         L1_1_L2_4_G1_MINI_ALU_nx403, L1_1_L2_4_G1_MINI_ALU_nx405, 
         L1_1_L2_4_G1_MINI_ALU_nx409, L1_1_L2_4_G1_MINI_ALU_nx411, 
         L1_1_L2_4_G1_MINI_ALU_nx413, L1_1_L2_4_G1_MINI_ALU_nx415, 
         L1_1_L2_4_G1_MINI_ALU_nx419, L1_1_L2_4_G1_MINI_ALU_nx421, 
         L1_1_L2_4_G1_MINI_ALU_nx423, L1_1_L2_4_G1_MINI_ALU_nx425, 
         L1_1_L2_4_G1_MINI_ALU_nx429, L1_1_L2_4_G1_MINI_ALU_nx431, 
         L1_1_L2_4_G1_MINI_ALU_nx433, L1_1_L2_4_G1_MINI_ALU_nx435, 
         L1_1_L2_4_G1_MINI_ALU_nx439, L1_1_L2_4_G1_MINI_ALU_nx441, 
         L1_1_L2_4_G1_MINI_ALU_nx443, L1_1_L2_4_G1_MINI_ALU_nx445, 
         L1_1_L2_4_G1_MINI_ALU_nx449, L1_1_L2_4_G1_MINI_ALU_nx451, 
         L1_1_L2_4_G1_MINI_ALU_nx453, L1_1_L2_4_G1_MINI_ALU_nx455, 
         L1_1_L2_4_G1_MINI_ALU_nx461, L1_1_L2_4_G1_MINI_ALU_nx463, 
         L1_1_L2_4_G1_MINI_ALU_nx467, L1_1_L2_4_G1_MINI_ALU_nx469, 
         L1_1_L2_4_G1_MINI_ALU_nx471, L1_1_L2_4_G1_MINI_ALU_nx475, 
         L1_1_L2_4_G1_MINI_ALU_nx477, L1_1_L2_4_G1_MINI_ALU_nx479, 
         L1_1_L2_4_G1_MINI_ALU_nx483, L1_1_L2_4_G1_MINI_ALU_nx485, 
         L1_1_L2_4_G1_MINI_ALU_nx487, L1_1_L2_4_G1_MINI_ALU_nx491, 
         L1_1_L2_4_G1_MINI_ALU_nx493, L1_1_L2_4_G1_MINI_ALU_nx495, 
         L1_1_L2_4_G1_MINI_ALU_nx499, L1_1_L2_4_G1_MINI_ALU_nx501, 
         L1_1_L2_4_G1_MINI_ALU_nx503, L1_1_L2_4_G1_MINI_ALU_nx507, 
         L1_1_L2_4_G1_MINI_ALU_nx509, L1_1_L2_4_G1_MINI_ALU_nx511, 
         L1_1_L2_4_G1_MINI_ALU_nx515, L1_1_L2_4_G1_MINI_ALU_nx517, 
         L1_1_L2_4_G1_MINI_ALU_nx529, L1_1_L2_4_G1_MINI_ALU_nx531, 
         L1_1_L2_4_G1_MINI_ALU_nx534, L1_1_L2_4_G1_MINI_ALU_nx537, 
         L1_1_L2_4_G1_MINI_ALU_nx540, L1_1_L2_4_G1_MINI_ALU_nx544, 
         L1_1_L2_4_G1_MINI_ALU_nx547, L1_1_L2_4_G1_MINI_ALU_nx551, 
         L1_1_L2_4_G1_MINI_ALU_nx554, L1_1_L2_4_G1_MINI_ALU_nx558, 
         L1_1_L2_4_G1_MINI_ALU_nx561, L1_1_L2_4_G1_MINI_ALU_nx565, 
         L1_1_L2_4_G1_MINI_ALU_nx568, 
         L1_1_L2_4_G1_MINI_ALU_WindowCellShiftedLeft_16, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_16, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_15, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_14, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_13, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_12, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_11, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_10, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_16, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_15, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_14, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_13, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_12, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_11, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_10, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_9, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_8, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_7, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_6, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_5, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_4, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_3, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_2, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_1, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_0, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_16, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_15, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_14, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_13, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_12, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_11, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_10, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_9, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_8, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_7, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_6, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_5, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_4, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_3, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_2, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_1, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_0, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_16, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_15, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_14, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_13, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_12, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_11, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_10, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_9, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_8, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_7, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_6, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_5, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_4, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_3, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_2, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_1, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_0, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx4, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx8, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx12, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx16, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx20, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx24, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx80, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx328, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx384, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642, 
         L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644, 
         L1_2_L2_0_G1_MINI_ALU_AddPToBoothOperand, 
         L1_2_L2_0_G1_MINI_ALU_BoothOperand_16, 
         L1_2_L2_0_G1_MINI_ALU_BoothOperand_15, 
         L1_2_L2_0_G1_MINI_ALU_BoothOperand_14, 
         L1_2_L2_0_G1_MINI_ALU_BoothOperand_13, 
         L1_2_L2_0_G1_MINI_ALU_BoothOperand_12, 
         L1_2_L2_0_G1_MINI_ALU_BoothOperand_11, 
         L1_2_L2_0_G1_MINI_ALU_BoothOperand_10, 
         L1_2_L2_0_G1_MINI_ALU_BoothOperand_9, 
         L1_2_L2_0_G1_MINI_ALU_BoothOperand_8, 
         L1_2_L2_0_G1_MINI_ALU_BoothOperand_7, 
         L1_2_L2_0_G1_MINI_ALU_BoothOperand_6, 
         L1_2_L2_0_G1_MINI_ALU_BoothOperand_5, 
         L1_2_L2_0_G1_MINI_ALU_BoothOperand_4, 
         L1_2_L2_0_G1_MINI_ALU_BoothOperand_3, 
         L1_2_L2_0_G1_MINI_ALU_BoothOperand_2, 
         L1_2_L2_0_G1_MINI_ALU_BoothOperand_1, 
         L1_2_L2_0_G1_MINI_ALU_BoothOperand_0, 
         L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_16, 
         L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_15, 
         L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_14, 
         L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_13, 
         L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_12, 
         L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_11, 
         L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_10, 
         L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_9, 
         L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_8, 
         L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_7, 
         L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_6, 
         L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_5, 
         L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_4, 
         L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_3, 
         L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_2, 
         L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_1, 
         L1_2_L2_0_G1_MINI_ALU_BoothP_16, L1_2_L2_0_G1_MINI_ALU_BoothP_15, 
         L1_2_L2_0_G1_MINI_ALU_BoothP_14, L1_2_L2_0_G1_MINI_ALU_BoothP_13, 
         L1_2_L2_0_G1_MINI_ALU_BoothP_12, L1_2_L2_0_G1_MINI_ALU_BoothP_11, 
         L1_2_L2_0_G1_MINI_ALU_BoothP_10, L1_2_L2_0_G1_MINI_ALU_BoothP_9, 
         L1_2_L2_0_G1_MINI_ALU_BoothP_8, L1_2_L2_0_G1_MINI_ALU_BoothP_7, 
         L1_2_L2_0_G1_MINI_ALU_BoothP_6, L1_2_L2_0_G1_MINI_ALU_BoothP_5, 
         L1_2_L2_0_G1_MINI_ALU_BoothP_4, L1_2_L2_0_G1_MINI_ALU_BoothP_3, 
         L1_2_L2_0_G1_MINI_ALU_BoothP_2, L1_2_L2_0_G1_MINI_ALU_BoothP_1, 
         L1_2_L2_0_G1_MINI_ALU_BoothP_0, L1_2_L2_0_G1_MINI_ALU_nx0, 
         L1_2_L2_0_G1_MINI_ALU_nx6, L1_2_L2_0_G1_MINI_ALU_nx12, 
         L1_2_L2_0_G1_MINI_ALU_nx18, L1_2_L2_0_G1_MINI_ALU_nx24, 
         L1_2_L2_0_G1_MINI_ALU_nx30, L1_2_L2_0_G1_MINI_ALU_nx40, 
         L1_2_L2_0_G1_MINI_ALU_nx44, L1_2_L2_0_G1_MINI_ALU_nx48, 
         L1_2_L2_0_G1_MINI_ALU_nx52, L1_2_L2_0_G1_MINI_ALU_nx56, 
         L1_2_L2_0_G1_MINI_ALU_nx62, L1_2_L2_0_G1_MINI_ALU_nx154, 
         L1_2_L2_0_G1_MINI_ALU_nx316, L1_2_L2_0_G1_MINI_ALU_nx336, 
         L1_2_L2_0_G1_MINI_ALU_nx356, L1_2_L2_0_G1_MINI_ALU_nx376, 
         L1_2_L2_0_G1_MINI_ALU_nx396, L1_2_L2_0_G1_MINI_ALU_nx416, 
         L1_2_L2_0_G1_MINI_ALU_nx436, L1_2_L2_0_G1_MINI_ALU_nx454, 
         L1_2_L2_0_G1_MINI_ALU_nx456, L1_2_L2_0_G1_MINI_ALU_nx379, 
         L1_2_L2_0_G1_MINI_ALU_nx381, L1_2_L2_0_G1_MINI_ALU_nx383, 
         L1_2_L2_0_G1_MINI_ALU_nx387, L1_2_L2_0_G1_MINI_ALU_nx389, 
         L1_2_L2_0_G1_MINI_ALU_nx391, L1_2_L2_0_G1_MINI_ALU_nx395, 
         L1_2_L2_0_G1_MINI_ALU_nx399, L1_2_L2_0_G1_MINI_ALU_nx401, 
         L1_2_L2_0_G1_MINI_ALU_nx403, L1_2_L2_0_G1_MINI_ALU_nx405, 
         L1_2_L2_0_G1_MINI_ALU_nx409, L1_2_L2_0_G1_MINI_ALU_nx411, 
         L1_2_L2_0_G1_MINI_ALU_nx413, L1_2_L2_0_G1_MINI_ALU_nx415, 
         L1_2_L2_0_G1_MINI_ALU_nx419, L1_2_L2_0_G1_MINI_ALU_nx421, 
         L1_2_L2_0_G1_MINI_ALU_nx423, L1_2_L2_0_G1_MINI_ALU_nx425, 
         L1_2_L2_0_G1_MINI_ALU_nx429, L1_2_L2_0_G1_MINI_ALU_nx431, 
         L1_2_L2_0_G1_MINI_ALU_nx433, L1_2_L2_0_G1_MINI_ALU_nx435, 
         L1_2_L2_0_G1_MINI_ALU_nx439, L1_2_L2_0_G1_MINI_ALU_nx441, 
         L1_2_L2_0_G1_MINI_ALU_nx443, L1_2_L2_0_G1_MINI_ALU_nx445, 
         L1_2_L2_0_G1_MINI_ALU_nx449, L1_2_L2_0_G1_MINI_ALU_nx451, 
         L1_2_L2_0_G1_MINI_ALU_nx453, L1_2_L2_0_G1_MINI_ALU_nx455, 
         L1_2_L2_0_G1_MINI_ALU_nx461, L1_2_L2_0_G1_MINI_ALU_nx463, 
         L1_2_L2_0_G1_MINI_ALU_nx467, L1_2_L2_0_G1_MINI_ALU_nx469, 
         L1_2_L2_0_G1_MINI_ALU_nx471, L1_2_L2_0_G1_MINI_ALU_nx475, 
         L1_2_L2_0_G1_MINI_ALU_nx477, L1_2_L2_0_G1_MINI_ALU_nx479, 
         L1_2_L2_0_G1_MINI_ALU_nx483, L1_2_L2_0_G1_MINI_ALU_nx485, 
         L1_2_L2_0_G1_MINI_ALU_nx487, L1_2_L2_0_G1_MINI_ALU_nx491, 
         L1_2_L2_0_G1_MINI_ALU_nx493, L1_2_L2_0_G1_MINI_ALU_nx495, 
         L1_2_L2_0_G1_MINI_ALU_nx499, L1_2_L2_0_G1_MINI_ALU_nx501, 
         L1_2_L2_0_G1_MINI_ALU_nx503, L1_2_L2_0_G1_MINI_ALU_nx507, 
         L1_2_L2_0_G1_MINI_ALU_nx509, L1_2_L2_0_G1_MINI_ALU_nx511, 
         L1_2_L2_0_G1_MINI_ALU_nx515, L1_2_L2_0_G1_MINI_ALU_nx517, 
         L1_2_L2_0_G1_MINI_ALU_nx529, L1_2_L2_0_G1_MINI_ALU_nx531, 
         L1_2_L2_0_G1_MINI_ALU_nx534, L1_2_L2_0_G1_MINI_ALU_nx537, 
         L1_2_L2_0_G1_MINI_ALU_nx540, L1_2_L2_0_G1_MINI_ALU_nx544, 
         L1_2_L2_0_G1_MINI_ALU_nx547, L1_2_L2_0_G1_MINI_ALU_nx551, 
         L1_2_L2_0_G1_MINI_ALU_nx554, L1_2_L2_0_G1_MINI_ALU_nx558, 
         L1_2_L2_0_G1_MINI_ALU_nx561, L1_2_L2_0_G1_MINI_ALU_nx565, 
         L1_2_L2_0_G1_MINI_ALU_nx568, 
         L1_2_L2_0_G1_MINI_ALU_WindowCellShiftedLeft_16, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_16, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_15, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_14, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_13, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_12, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_11, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_10, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_16, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_15, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_14, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_13, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_12, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_11, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_10, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_9, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_8, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_7, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_6, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_5, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_4, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_3, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_2, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_1, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_0, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_16, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_15, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_14, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_13, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_12, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_11, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_10, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_9, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_8, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_7, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_6, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_5, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_4, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_3, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_2, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_1, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_0, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_16, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_15, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_14, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_13, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_12, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_11, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_10, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_9, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_8, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_7, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_6, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_5, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_4, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_3, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_2, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_1, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_0, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx4, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx8, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx12, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx16, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx20, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx24, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx80, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx328, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx384, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642, 
         L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644, 
         L1_2_L2_1_G1_MINI_ALU_AddPToBoothOperand, 
         L1_2_L2_1_G1_MINI_ALU_BoothOperand_16, 
         L1_2_L2_1_G1_MINI_ALU_BoothOperand_15, 
         L1_2_L2_1_G1_MINI_ALU_BoothOperand_14, 
         L1_2_L2_1_G1_MINI_ALU_BoothOperand_13, 
         L1_2_L2_1_G1_MINI_ALU_BoothOperand_12, 
         L1_2_L2_1_G1_MINI_ALU_BoothOperand_11, 
         L1_2_L2_1_G1_MINI_ALU_BoothOperand_10, 
         L1_2_L2_1_G1_MINI_ALU_BoothOperand_9, 
         L1_2_L2_1_G1_MINI_ALU_BoothOperand_8, 
         L1_2_L2_1_G1_MINI_ALU_BoothOperand_7, 
         L1_2_L2_1_G1_MINI_ALU_BoothOperand_6, 
         L1_2_L2_1_G1_MINI_ALU_BoothOperand_5, 
         L1_2_L2_1_G1_MINI_ALU_BoothOperand_4, 
         L1_2_L2_1_G1_MINI_ALU_BoothOperand_3, 
         L1_2_L2_1_G1_MINI_ALU_BoothOperand_2, 
         L1_2_L2_1_G1_MINI_ALU_BoothOperand_1, 
         L1_2_L2_1_G1_MINI_ALU_BoothOperand_0, 
         L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_16, 
         L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_15, 
         L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_14, 
         L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_13, 
         L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_12, 
         L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_11, 
         L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_10, 
         L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_9, 
         L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_8, 
         L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_7, 
         L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_6, 
         L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_5, 
         L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_4, 
         L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_3, 
         L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_2, 
         L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_1, 
         L1_2_L2_1_G1_MINI_ALU_BoothP_16, L1_2_L2_1_G1_MINI_ALU_BoothP_15, 
         L1_2_L2_1_G1_MINI_ALU_BoothP_14, L1_2_L2_1_G1_MINI_ALU_BoothP_13, 
         L1_2_L2_1_G1_MINI_ALU_BoothP_12, L1_2_L2_1_G1_MINI_ALU_BoothP_11, 
         L1_2_L2_1_G1_MINI_ALU_BoothP_10, L1_2_L2_1_G1_MINI_ALU_BoothP_9, 
         L1_2_L2_1_G1_MINI_ALU_BoothP_8, L1_2_L2_1_G1_MINI_ALU_BoothP_7, 
         L1_2_L2_1_G1_MINI_ALU_BoothP_6, L1_2_L2_1_G1_MINI_ALU_BoothP_5, 
         L1_2_L2_1_G1_MINI_ALU_BoothP_4, L1_2_L2_1_G1_MINI_ALU_BoothP_3, 
         L1_2_L2_1_G1_MINI_ALU_BoothP_2, L1_2_L2_1_G1_MINI_ALU_BoothP_1, 
         L1_2_L2_1_G1_MINI_ALU_BoothP_0, L1_2_L2_1_G1_MINI_ALU_nx0, 
         L1_2_L2_1_G1_MINI_ALU_nx6, L1_2_L2_1_G1_MINI_ALU_nx12, 
         L1_2_L2_1_G1_MINI_ALU_nx18, L1_2_L2_1_G1_MINI_ALU_nx24, 
         L1_2_L2_1_G1_MINI_ALU_nx30, L1_2_L2_1_G1_MINI_ALU_nx40, 
         L1_2_L2_1_G1_MINI_ALU_nx44, L1_2_L2_1_G1_MINI_ALU_nx48, 
         L1_2_L2_1_G1_MINI_ALU_nx52, L1_2_L2_1_G1_MINI_ALU_nx56, 
         L1_2_L2_1_G1_MINI_ALU_nx62, L1_2_L2_1_G1_MINI_ALU_nx154, 
         L1_2_L2_1_G1_MINI_ALU_nx316, L1_2_L2_1_G1_MINI_ALU_nx336, 
         L1_2_L2_1_G1_MINI_ALU_nx356, L1_2_L2_1_G1_MINI_ALU_nx376, 
         L1_2_L2_1_G1_MINI_ALU_nx396, L1_2_L2_1_G1_MINI_ALU_nx416, 
         L1_2_L2_1_G1_MINI_ALU_nx436, L1_2_L2_1_G1_MINI_ALU_nx454, 
         L1_2_L2_1_G1_MINI_ALU_nx456, L1_2_L2_1_G1_MINI_ALU_nx379, 
         L1_2_L2_1_G1_MINI_ALU_nx381, L1_2_L2_1_G1_MINI_ALU_nx383, 
         L1_2_L2_1_G1_MINI_ALU_nx387, L1_2_L2_1_G1_MINI_ALU_nx389, 
         L1_2_L2_1_G1_MINI_ALU_nx391, L1_2_L2_1_G1_MINI_ALU_nx395, 
         L1_2_L2_1_G1_MINI_ALU_nx399, L1_2_L2_1_G1_MINI_ALU_nx401, 
         L1_2_L2_1_G1_MINI_ALU_nx403, L1_2_L2_1_G1_MINI_ALU_nx405, 
         L1_2_L2_1_G1_MINI_ALU_nx409, L1_2_L2_1_G1_MINI_ALU_nx411, 
         L1_2_L2_1_G1_MINI_ALU_nx413, L1_2_L2_1_G1_MINI_ALU_nx415, 
         L1_2_L2_1_G1_MINI_ALU_nx419, L1_2_L2_1_G1_MINI_ALU_nx421, 
         L1_2_L2_1_G1_MINI_ALU_nx423, L1_2_L2_1_G1_MINI_ALU_nx425, 
         L1_2_L2_1_G1_MINI_ALU_nx429, L1_2_L2_1_G1_MINI_ALU_nx431, 
         L1_2_L2_1_G1_MINI_ALU_nx433, L1_2_L2_1_G1_MINI_ALU_nx435, 
         L1_2_L2_1_G1_MINI_ALU_nx439, L1_2_L2_1_G1_MINI_ALU_nx441, 
         L1_2_L2_1_G1_MINI_ALU_nx443, L1_2_L2_1_G1_MINI_ALU_nx445, 
         L1_2_L2_1_G1_MINI_ALU_nx449, L1_2_L2_1_G1_MINI_ALU_nx451, 
         L1_2_L2_1_G1_MINI_ALU_nx453, L1_2_L2_1_G1_MINI_ALU_nx455, 
         L1_2_L2_1_G1_MINI_ALU_nx461, L1_2_L2_1_G1_MINI_ALU_nx463, 
         L1_2_L2_1_G1_MINI_ALU_nx467, L1_2_L2_1_G1_MINI_ALU_nx469, 
         L1_2_L2_1_G1_MINI_ALU_nx471, L1_2_L2_1_G1_MINI_ALU_nx475, 
         L1_2_L2_1_G1_MINI_ALU_nx477, L1_2_L2_1_G1_MINI_ALU_nx479, 
         L1_2_L2_1_G1_MINI_ALU_nx483, L1_2_L2_1_G1_MINI_ALU_nx485, 
         L1_2_L2_1_G1_MINI_ALU_nx487, L1_2_L2_1_G1_MINI_ALU_nx491, 
         L1_2_L2_1_G1_MINI_ALU_nx493, L1_2_L2_1_G1_MINI_ALU_nx495, 
         L1_2_L2_1_G1_MINI_ALU_nx499, L1_2_L2_1_G1_MINI_ALU_nx501, 
         L1_2_L2_1_G1_MINI_ALU_nx503, L1_2_L2_1_G1_MINI_ALU_nx507, 
         L1_2_L2_1_G1_MINI_ALU_nx509, L1_2_L2_1_G1_MINI_ALU_nx511, 
         L1_2_L2_1_G1_MINI_ALU_nx515, L1_2_L2_1_G1_MINI_ALU_nx517, 
         L1_2_L2_1_G1_MINI_ALU_nx529, L1_2_L2_1_G1_MINI_ALU_nx531, 
         L1_2_L2_1_G1_MINI_ALU_nx534, L1_2_L2_1_G1_MINI_ALU_nx537, 
         L1_2_L2_1_G1_MINI_ALU_nx540, L1_2_L2_1_G1_MINI_ALU_nx544, 
         L1_2_L2_1_G1_MINI_ALU_nx547, L1_2_L2_1_G1_MINI_ALU_nx551, 
         L1_2_L2_1_G1_MINI_ALU_nx554, L1_2_L2_1_G1_MINI_ALU_nx558, 
         L1_2_L2_1_G1_MINI_ALU_nx561, L1_2_L2_1_G1_MINI_ALU_nx565, 
         L1_2_L2_1_G1_MINI_ALU_nx568, 
         L1_2_L2_1_G1_MINI_ALU_WindowCellShiftedLeft_16, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_16, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_15, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_14, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_13, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_12, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_11, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_10, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_16, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_15, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_14, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_13, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_12, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_11, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_10, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_9, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_8, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_7, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_6, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_5, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_4, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_3, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_2, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_1, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_0, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_16, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_15, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_14, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_13, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_12, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_11, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_10, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_9, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_8, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_7, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_6, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_5, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_4, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_3, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_2, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_1, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_0, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_16, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_15, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_14, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_13, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_12, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_11, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_10, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_9, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_8, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_7, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_6, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_5, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_4, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_3, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_2, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_1, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_0, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx4, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx8, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx12, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx16, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx20, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx24, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx80, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx328, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx384, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642, 
         L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644, 
         L1_2_L2_2_G1_MINI_ALU_AddPToBoothOperand, 
         L1_2_L2_2_G1_MINI_ALU_BoothOperand_16, 
         L1_2_L2_2_G1_MINI_ALU_BoothOperand_15, 
         L1_2_L2_2_G1_MINI_ALU_BoothOperand_14, 
         L1_2_L2_2_G1_MINI_ALU_BoothOperand_13, 
         L1_2_L2_2_G1_MINI_ALU_BoothOperand_12, 
         L1_2_L2_2_G1_MINI_ALU_BoothOperand_11, 
         L1_2_L2_2_G1_MINI_ALU_BoothOperand_10, 
         L1_2_L2_2_G1_MINI_ALU_BoothOperand_9, 
         L1_2_L2_2_G1_MINI_ALU_BoothOperand_8, 
         L1_2_L2_2_G1_MINI_ALU_BoothOperand_7, 
         L1_2_L2_2_G1_MINI_ALU_BoothOperand_6, 
         L1_2_L2_2_G1_MINI_ALU_BoothOperand_5, 
         L1_2_L2_2_G1_MINI_ALU_BoothOperand_4, 
         L1_2_L2_2_G1_MINI_ALU_BoothOperand_3, 
         L1_2_L2_2_G1_MINI_ALU_BoothOperand_2, 
         L1_2_L2_2_G1_MINI_ALU_BoothOperand_1, 
         L1_2_L2_2_G1_MINI_ALU_BoothOperand_0, 
         L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_16, 
         L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_15, 
         L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_14, 
         L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_13, 
         L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_12, 
         L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_11, 
         L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_10, 
         L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_9, 
         L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_8, 
         L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_7, 
         L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_6, 
         L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_5, 
         L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_4, 
         L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_3, 
         L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_2, 
         L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_1, 
         L1_2_L2_2_G1_MINI_ALU_BoothP_16, L1_2_L2_2_G1_MINI_ALU_BoothP_15, 
         L1_2_L2_2_G1_MINI_ALU_BoothP_14, L1_2_L2_2_G1_MINI_ALU_BoothP_13, 
         L1_2_L2_2_G1_MINI_ALU_BoothP_12, L1_2_L2_2_G1_MINI_ALU_BoothP_11, 
         L1_2_L2_2_G1_MINI_ALU_BoothP_10, L1_2_L2_2_G1_MINI_ALU_BoothP_9, 
         L1_2_L2_2_G1_MINI_ALU_BoothP_8, L1_2_L2_2_G1_MINI_ALU_BoothP_7, 
         L1_2_L2_2_G1_MINI_ALU_BoothP_6, L1_2_L2_2_G1_MINI_ALU_BoothP_5, 
         L1_2_L2_2_G1_MINI_ALU_BoothP_4, L1_2_L2_2_G1_MINI_ALU_BoothP_3, 
         L1_2_L2_2_G1_MINI_ALU_BoothP_2, L1_2_L2_2_G1_MINI_ALU_BoothP_1, 
         L1_2_L2_2_G1_MINI_ALU_BoothP_0, L1_2_L2_2_G1_MINI_ALU_nx154, 
         L1_2_L2_2_G1_MINI_ALU_nx316, L1_2_L2_2_G1_MINI_ALU_nx336, 
         L1_2_L2_2_G1_MINI_ALU_nx356, L1_2_L2_2_G1_MINI_ALU_nx376, 
         L1_2_L2_2_G1_MINI_ALU_nx396, L1_2_L2_2_G1_MINI_ALU_nx416, 
         L1_2_L2_2_G1_MINI_ALU_nx436, L1_2_L2_2_G1_MINI_ALU_nx454, 
         L1_2_L2_2_G1_MINI_ALU_nx456, L1_2_L2_2_G1_MINI_ALU_nx379, 
         L1_2_L2_2_G1_MINI_ALU_nx381, L1_2_L2_2_G1_MINI_ALU_nx383, 
         L1_2_L2_2_G1_MINI_ALU_nx387, L1_2_L2_2_G1_MINI_ALU_nx389, 
         L1_2_L2_2_G1_MINI_ALU_nx391, L1_2_L2_2_G1_MINI_ALU_nx395, 
         L1_2_L2_2_G1_MINI_ALU_nx399, L1_2_L2_2_G1_MINI_ALU_nx401, 
         L1_2_L2_2_G1_MINI_ALU_nx403, L1_2_L2_2_G1_MINI_ALU_nx405, 
         L1_2_L2_2_G1_MINI_ALU_nx409, L1_2_L2_2_G1_MINI_ALU_nx411, 
         L1_2_L2_2_G1_MINI_ALU_nx413, L1_2_L2_2_G1_MINI_ALU_nx415, 
         L1_2_L2_2_G1_MINI_ALU_nx419, L1_2_L2_2_G1_MINI_ALU_nx421, 
         L1_2_L2_2_G1_MINI_ALU_nx423, L1_2_L2_2_G1_MINI_ALU_nx425, 
         L1_2_L2_2_G1_MINI_ALU_nx429, L1_2_L2_2_G1_MINI_ALU_nx431, 
         L1_2_L2_2_G1_MINI_ALU_nx433, L1_2_L2_2_G1_MINI_ALU_nx435, 
         L1_2_L2_2_G1_MINI_ALU_nx439, L1_2_L2_2_G1_MINI_ALU_nx441, 
         L1_2_L2_2_G1_MINI_ALU_nx443, L1_2_L2_2_G1_MINI_ALU_nx445, 
         L1_2_L2_2_G1_MINI_ALU_nx449, L1_2_L2_2_G1_MINI_ALU_nx451, 
         L1_2_L2_2_G1_MINI_ALU_nx453, L1_2_L2_2_G1_MINI_ALU_nx455, 
         L1_2_L2_2_G1_MINI_ALU_nx461, L1_2_L2_2_G1_MINI_ALU_nx463, 
         L1_2_L2_2_G1_MINI_ALU_nx467, L1_2_L2_2_G1_MINI_ALU_nx469, 
         L1_2_L2_2_G1_MINI_ALU_nx471, L1_2_L2_2_G1_MINI_ALU_nx475, 
         L1_2_L2_2_G1_MINI_ALU_nx477, L1_2_L2_2_G1_MINI_ALU_nx479, 
         L1_2_L2_2_G1_MINI_ALU_nx483, L1_2_L2_2_G1_MINI_ALU_nx485, 
         L1_2_L2_2_G1_MINI_ALU_nx487, L1_2_L2_2_G1_MINI_ALU_nx491, 
         L1_2_L2_2_G1_MINI_ALU_nx493, L1_2_L2_2_G1_MINI_ALU_nx495, 
         L1_2_L2_2_G1_MINI_ALU_nx499, L1_2_L2_2_G1_MINI_ALU_nx501, 
         L1_2_L2_2_G1_MINI_ALU_nx503, L1_2_L2_2_G1_MINI_ALU_nx507, 
         L1_2_L2_2_G1_MINI_ALU_nx509, L1_2_L2_2_G1_MINI_ALU_nx511, 
         L1_2_L2_2_G1_MINI_ALU_nx515, L1_2_L2_2_G1_MINI_ALU_nx517, 
         L1_2_L2_2_G1_MINI_ALU_WindowCellShiftedLeft_16, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_16, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_15, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_14, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_13, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_12, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_11, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_10, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_16, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_15, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_14, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_13, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_12, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_11, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_10, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_9, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_8, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_7, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_6, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_5, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_4, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_3, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_2, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_1, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_0, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_16, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_15, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_14, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_13, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_12, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_11, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_10, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_9, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_8, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_7, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_6, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_5, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_4, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_3, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_2, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_1, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_0, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_16, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_15, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_14, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_13, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_12, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_11, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_10, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_9, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_8, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_7, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_6, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_5, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_4, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_3, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_2, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_1, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_0, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx4, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx8, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx12, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx16, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx20, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx24, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx80, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx328, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx384, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642, 
         L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644, 
         L1_2_L2_3_G2_MINI_ALU_AddPToBoothOperand, 
         L1_2_L2_3_G2_MINI_ALU_BoothOperand_16, 
         L1_2_L2_3_G2_MINI_ALU_BoothOperand_15, 
         L1_2_L2_3_G2_MINI_ALU_BoothOperand_14, 
         L1_2_L2_3_G2_MINI_ALU_BoothOperand_13, 
         L1_2_L2_3_G2_MINI_ALU_BoothOperand_12, 
         L1_2_L2_3_G2_MINI_ALU_BoothOperand_11, 
         L1_2_L2_3_G2_MINI_ALU_BoothOperand_10, 
         L1_2_L2_3_G2_MINI_ALU_BoothOperand_9, 
         L1_2_L2_3_G2_MINI_ALU_BoothOperand_8, 
         L1_2_L2_3_G2_MINI_ALU_BoothOperand_7, 
         L1_2_L2_3_G2_MINI_ALU_BoothOperand_6, 
         L1_2_L2_3_G2_MINI_ALU_BoothOperand_5, 
         L1_2_L2_3_G2_MINI_ALU_BoothOperand_4, 
         L1_2_L2_3_G2_MINI_ALU_BoothOperand_3, 
         L1_2_L2_3_G2_MINI_ALU_BoothOperand_2, 
         L1_2_L2_3_G2_MINI_ALU_BoothOperand_1, 
         L1_2_L2_3_G2_MINI_ALU_BoothOperand_0, 
         L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_16, 
         L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_15, 
         L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_14, 
         L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_13, 
         L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_12, 
         L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_11, 
         L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_10, 
         L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_9, 
         L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_8, 
         L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_7, 
         L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_6, 
         L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_5, 
         L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_4, 
         L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_3, 
         L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_2, 
         L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_1, 
         L1_2_L2_3_G2_MINI_ALU_BoothP_16, L1_2_L2_3_G2_MINI_ALU_BoothP_15, 
         L1_2_L2_3_G2_MINI_ALU_BoothP_14, L1_2_L2_3_G2_MINI_ALU_BoothP_13, 
         L1_2_L2_3_G2_MINI_ALU_BoothP_12, L1_2_L2_3_G2_MINI_ALU_BoothP_11, 
         L1_2_L2_3_G2_MINI_ALU_BoothP_10, L1_2_L2_3_G2_MINI_ALU_BoothP_9, 
         L1_2_L2_3_G2_MINI_ALU_BoothP_8, L1_2_L2_3_G2_MINI_ALU_BoothP_7, 
         L1_2_L2_3_G2_MINI_ALU_BoothP_6, L1_2_L2_3_G2_MINI_ALU_BoothP_5, 
         L1_2_L2_3_G2_MINI_ALU_BoothP_4, L1_2_L2_3_G2_MINI_ALU_BoothP_3, 
         L1_2_L2_3_G2_MINI_ALU_BoothP_2, L1_2_L2_3_G2_MINI_ALU_BoothP_1, 
         L1_2_L2_3_G2_MINI_ALU_BoothP_0, L1_2_L2_3_G2_MINI_ALU_nx0, 
         L1_2_L2_3_G2_MINI_ALU_nx6, L1_2_L2_3_G2_MINI_ALU_nx12, 
         L1_2_L2_3_G2_MINI_ALU_nx18, L1_2_L2_3_G2_MINI_ALU_nx24, 
         L1_2_L2_3_G2_MINI_ALU_nx30, L1_2_L2_3_G2_MINI_ALU_nx40, 
         L1_2_L2_3_G2_MINI_ALU_nx44, L1_2_L2_3_G2_MINI_ALU_nx48, 
         L1_2_L2_3_G2_MINI_ALU_nx52, L1_2_L2_3_G2_MINI_ALU_nx56, 
         L1_2_L2_3_G2_MINI_ALU_nx62, L1_2_L2_3_G2_MINI_ALU_nx154, 
         L1_2_L2_3_G2_MINI_ALU_nx316, L1_2_L2_3_G2_MINI_ALU_nx336, 
         L1_2_L2_3_G2_MINI_ALU_nx356, L1_2_L2_3_G2_MINI_ALU_nx376, 
         L1_2_L2_3_G2_MINI_ALU_nx396, L1_2_L2_3_G2_MINI_ALU_nx416, 
         L1_2_L2_3_G2_MINI_ALU_nx436, L1_2_L2_3_G2_MINI_ALU_nx454, 
         L1_2_L2_3_G2_MINI_ALU_nx456, L1_2_L2_3_G2_MINI_ALU_nx379, 
         L1_2_L2_3_G2_MINI_ALU_nx381, L1_2_L2_3_G2_MINI_ALU_nx383, 
         L1_2_L2_3_G2_MINI_ALU_nx387, L1_2_L2_3_G2_MINI_ALU_nx389, 
         L1_2_L2_3_G2_MINI_ALU_nx391, L1_2_L2_3_G2_MINI_ALU_nx395, 
         L1_2_L2_3_G2_MINI_ALU_nx399, L1_2_L2_3_G2_MINI_ALU_nx401, 
         L1_2_L2_3_G2_MINI_ALU_nx403, L1_2_L2_3_G2_MINI_ALU_nx405, 
         L1_2_L2_3_G2_MINI_ALU_nx409, L1_2_L2_3_G2_MINI_ALU_nx411, 
         L1_2_L2_3_G2_MINI_ALU_nx413, L1_2_L2_3_G2_MINI_ALU_nx415, 
         L1_2_L2_3_G2_MINI_ALU_nx419, L1_2_L2_3_G2_MINI_ALU_nx421, 
         L1_2_L2_3_G2_MINI_ALU_nx423, L1_2_L2_3_G2_MINI_ALU_nx425, 
         L1_2_L2_3_G2_MINI_ALU_nx429, L1_2_L2_3_G2_MINI_ALU_nx431, 
         L1_2_L2_3_G2_MINI_ALU_nx433, L1_2_L2_3_G2_MINI_ALU_nx435, 
         L1_2_L2_3_G2_MINI_ALU_nx439, L1_2_L2_3_G2_MINI_ALU_nx441, 
         L1_2_L2_3_G2_MINI_ALU_nx443, L1_2_L2_3_G2_MINI_ALU_nx445, 
         L1_2_L2_3_G2_MINI_ALU_nx449, L1_2_L2_3_G2_MINI_ALU_nx451, 
         L1_2_L2_3_G2_MINI_ALU_nx453, L1_2_L2_3_G2_MINI_ALU_nx455, 
         L1_2_L2_3_G2_MINI_ALU_nx461, L1_2_L2_3_G2_MINI_ALU_nx463, 
         L1_2_L2_3_G2_MINI_ALU_nx467, L1_2_L2_3_G2_MINI_ALU_nx469, 
         L1_2_L2_3_G2_MINI_ALU_nx471, L1_2_L2_3_G2_MINI_ALU_nx475, 
         L1_2_L2_3_G2_MINI_ALU_nx477, L1_2_L2_3_G2_MINI_ALU_nx479, 
         L1_2_L2_3_G2_MINI_ALU_nx483, L1_2_L2_3_G2_MINI_ALU_nx485, 
         L1_2_L2_3_G2_MINI_ALU_nx487, L1_2_L2_3_G2_MINI_ALU_nx491, 
         L1_2_L2_3_G2_MINI_ALU_nx493, L1_2_L2_3_G2_MINI_ALU_nx495, 
         L1_2_L2_3_G2_MINI_ALU_nx499, L1_2_L2_3_G2_MINI_ALU_nx501, 
         L1_2_L2_3_G2_MINI_ALU_nx503, L1_2_L2_3_G2_MINI_ALU_nx507, 
         L1_2_L2_3_G2_MINI_ALU_nx509, L1_2_L2_3_G2_MINI_ALU_nx511, 
         L1_2_L2_3_G2_MINI_ALU_nx515, L1_2_L2_3_G2_MINI_ALU_nx517, 
         L1_2_L2_3_G2_MINI_ALU_nx529, L1_2_L2_3_G2_MINI_ALU_nx531, 
         L1_2_L2_3_G2_MINI_ALU_nx534, L1_2_L2_3_G2_MINI_ALU_nx537, 
         L1_2_L2_3_G2_MINI_ALU_nx540, L1_2_L2_3_G2_MINI_ALU_nx544, 
         L1_2_L2_3_G2_MINI_ALU_nx547, L1_2_L2_3_G2_MINI_ALU_nx551, 
         L1_2_L2_3_G2_MINI_ALU_nx554, L1_2_L2_3_G2_MINI_ALU_nx558, 
         L1_2_L2_3_G2_MINI_ALU_nx561, L1_2_L2_3_G2_MINI_ALU_nx565, 
         L1_2_L2_3_G2_MINI_ALU_nx568, 
         L1_2_L2_3_G2_MINI_ALU_WindowCellShiftedLeft_16, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_16, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_15, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_14, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_13, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_12, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_11, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_10, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_16, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_15, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_14, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_13, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_12, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_11, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_10, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_9, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_8, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_7, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_6, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_5, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_4, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_3, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_2, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_1, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_0, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_16, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_15, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_14, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_13, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_12, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_11, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_10, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_9, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_8, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_7, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_6, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_5, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_4, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_3, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_2, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_1, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_0, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_16, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_15, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_14, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_13, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_12, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_11, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_10, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_9, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_8, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_7, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_6, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_5, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_4, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_3, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_2, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_1, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_0, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx4, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx8, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx12, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx16, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx20, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx24, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx80, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx328, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx384, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642, 
         L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644, 
         L1_2_L2_4_G2_MINI_ALU_AddPToBoothOperand, 
         L1_2_L2_4_G2_MINI_ALU_BoothOperand_16, 
         L1_2_L2_4_G2_MINI_ALU_BoothOperand_15, 
         L1_2_L2_4_G2_MINI_ALU_BoothOperand_14, 
         L1_2_L2_4_G2_MINI_ALU_BoothOperand_13, 
         L1_2_L2_4_G2_MINI_ALU_BoothOperand_12, 
         L1_2_L2_4_G2_MINI_ALU_BoothOperand_11, 
         L1_2_L2_4_G2_MINI_ALU_BoothOperand_10, 
         L1_2_L2_4_G2_MINI_ALU_BoothOperand_9, 
         L1_2_L2_4_G2_MINI_ALU_BoothOperand_8, 
         L1_2_L2_4_G2_MINI_ALU_BoothOperand_7, 
         L1_2_L2_4_G2_MINI_ALU_BoothOperand_6, 
         L1_2_L2_4_G2_MINI_ALU_BoothOperand_5, 
         L1_2_L2_4_G2_MINI_ALU_BoothOperand_4, 
         L1_2_L2_4_G2_MINI_ALU_BoothOperand_3, 
         L1_2_L2_4_G2_MINI_ALU_BoothOperand_2, 
         L1_2_L2_4_G2_MINI_ALU_BoothOperand_1, 
         L1_2_L2_4_G2_MINI_ALU_BoothOperand_0, 
         L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_16, 
         L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_15, 
         L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_14, 
         L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_13, 
         L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_12, 
         L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_11, 
         L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_10, 
         L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_9, 
         L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_8, 
         L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_7, 
         L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_6, 
         L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_5, 
         L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_4, 
         L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_3, 
         L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_2, 
         L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_1, 
         L1_2_L2_4_G2_MINI_ALU_BoothP_16, L1_2_L2_4_G2_MINI_ALU_BoothP_15, 
         L1_2_L2_4_G2_MINI_ALU_BoothP_14, L1_2_L2_4_G2_MINI_ALU_BoothP_13, 
         L1_2_L2_4_G2_MINI_ALU_BoothP_12, L1_2_L2_4_G2_MINI_ALU_BoothP_11, 
         L1_2_L2_4_G2_MINI_ALU_BoothP_10, L1_2_L2_4_G2_MINI_ALU_BoothP_9, 
         L1_2_L2_4_G2_MINI_ALU_BoothP_8, L1_2_L2_4_G2_MINI_ALU_BoothP_7, 
         L1_2_L2_4_G2_MINI_ALU_BoothP_6, L1_2_L2_4_G2_MINI_ALU_BoothP_5, 
         L1_2_L2_4_G2_MINI_ALU_BoothP_4, L1_2_L2_4_G2_MINI_ALU_BoothP_3, 
         L1_2_L2_4_G2_MINI_ALU_BoothP_2, L1_2_L2_4_G2_MINI_ALU_BoothP_1, 
         L1_2_L2_4_G2_MINI_ALU_BoothP_0, L1_2_L2_4_G2_MINI_ALU_nx0, 
         L1_2_L2_4_G2_MINI_ALU_nx6, L1_2_L2_4_G2_MINI_ALU_nx12, 
         L1_2_L2_4_G2_MINI_ALU_nx18, L1_2_L2_4_G2_MINI_ALU_nx24, 
         L1_2_L2_4_G2_MINI_ALU_nx30, L1_2_L2_4_G2_MINI_ALU_nx40, 
         L1_2_L2_4_G2_MINI_ALU_nx44, L1_2_L2_4_G2_MINI_ALU_nx48, 
         L1_2_L2_4_G2_MINI_ALU_nx52, L1_2_L2_4_G2_MINI_ALU_nx56, 
         L1_2_L2_4_G2_MINI_ALU_nx62, L1_2_L2_4_G2_MINI_ALU_nx154, 
         L1_2_L2_4_G2_MINI_ALU_nx316, L1_2_L2_4_G2_MINI_ALU_nx336, 
         L1_2_L2_4_G2_MINI_ALU_nx356, L1_2_L2_4_G2_MINI_ALU_nx376, 
         L1_2_L2_4_G2_MINI_ALU_nx396, L1_2_L2_4_G2_MINI_ALU_nx416, 
         L1_2_L2_4_G2_MINI_ALU_nx436, L1_2_L2_4_G2_MINI_ALU_nx454, 
         L1_2_L2_4_G2_MINI_ALU_nx456, L1_2_L2_4_G2_MINI_ALU_nx379, 
         L1_2_L2_4_G2_MINI_ALU_nx381, L1_2_L2_4_G2_MINI_ALU_nx383, 
         L1_2_L2_4_G2_MINI_ALU_nx387, L1_2_L2_4_G2_MINI_ALU_nx389, 
         L1_2_L2_4_G2_MINI_ALU_nx391, L1_2_L2_4_G2_MINI_ALU_nx395, 
         L1_2_L2_4_G2_MINI_ALU_nx399, L1_2_L2_4_G2_MINI_ALU_nx401, 
         L1_2_L2_4_G2_MINI_ALU_nx403, L1_2_L2_4_G2_MINI_ALU_nx405, 
         L1_2_L2_4_G2_MINI_ALU_nx409, L1_2_L2_4_G2_MINI_ALU_nx411, 
         L1_2_L2_4_G2_MINI_ALU_nx413, L1_2_L2_4_G2_MINI_ALU_nx415, 
         L1_2_L2_4_G2_MINI_ALU_nx419, L1_2_L2_4_G2_MINI_ALU_nx421, 
         L1_2_L2_4_G2_MINI_ALU_nx423, L1_2_L2_4_G2_MINI_ALU_nx425, 
         L1_2_L2_4_G2_MINI_ALU_nx429, L1_2_L2_4_G2_MINI_ALU_nx431, 
         L1_2_L2_4_G2_MINI_ALU_nx433, L1_2_L2_4_G2_MINI_ALU_nx435, 
         L1_2_L2_4_G2_MINI_ALU_nx439, L1_2_L2_4_G2_MINI_ALU_nx441, 
         L1_2_L2_4_G2_MINI_ALU_nx443, L1_2_L2_4_G2_MINI_ALU_nx445, 
         L1_2_L2_4_G2_MINI_ALU_nx449, L1_2_L2_4_G2_MINI_ALU_nx451, 
         L1_2_L2_4_G2_MINI_ALU_nx453, L1_2_L2_4_G2_MINI_ALU_nx455, 
         L1_2_L2_4_G2_MINI_ALU_nx461, L1_2_L2_4_G2_MINI_ALU_nx463, 
         L1_2_L2_4_G2_MINI_ALU_nx467, L1_2_L2_4_G2_MINI_ALU_nx469, 
         L1_2_L2_4_G2_MINI_ALU_nx471, L1_2_L2_4_G2_MINI_ALU_nx475, 
         L1_2_L2_4_G2_MINI_ALU_nx477, L1_2_L2_4_G2_MINI_ALU_nx479, 
         L1_2_L2_4_G2_MINI_ALU_nx483, L1_2_L2_4_G2_MINI_ALU_nx485, 
         L1_2_L2_4_G2_MINI_ALU_nx487, L1_2_L2_4_G2_MINI_ALU_nx491, 
         L1_2_L2_4_G2_MINI_ALU_nx493, L1_2_L2_4_G2_MINI_ALU_nx495, 
         L1_2_L2_4_G2_MINI_ALU_nx499, L1_2_L2_4_G2_MINI_ALU_nx501, 
         L1_2_L2_4_G2_MINI_ALU_nx503, L1_2_L2_4_G2_MINI_ALU_nx507, 
         L1_2_L2_4_G2_MINI_ALU_nx509, L1_2_L2_4_G2_MINI_ALU_nx511, 
         L1_2_L2_4_G2_MINI_ALU_nx515, L1_2_L2_4_G2_MINI_ALU_nx517, 
         L1_2_L2_4_G2_MINI_ALU_nx529, L1_2_L2_4_G2_MINI_ALU_nx531, 
         L1_2_L2_4_G2_MINI_ALU_nx534, L1_2_L2_4_G2_MINI_ALU_nx537, 
         L1_2_L2_4_G2_MINI_ALU_nx540, L1_2_L2_4_G2_MINI_ALU_nx544, 
         L1_2_L2_4_G2_MINI_ALU_nx547, L1_2_L2_4_G2_MINI_ALU_nx551, 
         L1_2_L2_4_G2_MINI_ALU_nx554, L1_2_L2_4_G2_MINI_ALU_nx558, 
         L1_2_L2_4_G2_MINI_ALU_nx561, L1_2_L2_4_G2_MINI_ALU_nx565, 
         L1_2_L2_4_G2_MINI_ALU_nx568, 
         L1_2_L2_4_G2_MINI_ALU_WindowCellShiftedLeft_16, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_16, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_15, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_14, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_13, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_12, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_11, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_10, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_16, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_15, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_14, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_13, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_12, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_11, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_10, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_9, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_8, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_7, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_6, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_5, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_4, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_3, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_2, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_1, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_0, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_16, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_15, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_14, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_13, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_12, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_11, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_10, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_9, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_8, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_7, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_6, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_5, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_4, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_3, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_2, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_1, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_0, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_16, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_15, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_14, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_13, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_12, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_11, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_10, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_9, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_8, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_7, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_6, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_5, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_4, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_3, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_2, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_1, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_0, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_nx4, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_nx8, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_nx12, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_nx16, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_nx20, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_nx24, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_nx80, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_nx328, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_nx384, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642, 
         L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644, 
         L1_3_L2_0_G2_MINI_ALU_AddPToBoothOperand, 
         L1_3_L2_0_G2_MINI_ALU_BoothOperand_16, 
         L1_3_L2_0_G2_MINI_ALU_BoothOperand_15, 
         L1_3_L2_0_G2_MINI_ALU_BoothOperand_14, 
         L1_3_L2_0_G2_MINI_ALU_BoothOperand_13, 
         L1_3_L2_0_G2_MINI_ALU_BoothOperand_12, 
         L1_3_L2_0_G2_MINI_ALU_BoothOperand_11, 
         L1_3_L2_0_G2_MINI_ALU_BoothOperand_10, 
         L1_3_L2_0_G2_MINI_ALU_BoothOperand_9, 
         L1_3_L2_0_G2_MINI_ALU_BoothOperand_8, 
         L1_3_L2_0_G2_MINI_ALU_BoothOperand_7, 
         L1_3_L2_0_G2_MINI_ALU_BoothOperand_6, 
         L1_3_L2_0_G2_MINI_ALU_BoothOperand_5, 
         L1_3_L2_0_G2_MINI_ALU_BoothOperand_4, 
         L1_3_L2_0_G2_MINI_ALU_BoothOperand_3, 
         L1_3_L2_0_G2_MINI_ALU_BoothOperand_2, 
         L1_3_L2_0_G2_MINI_ALU_BoothOperand_1, 
         L1_3_L2_0_G2_MINI_ALU_BoothOperand_0, 
         L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_16, 
         L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_15, 
         L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_14, 
         L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_13, 
         L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_12, 
         L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_11, 
         L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_10, 
         L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_9, 
         L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_8, 
         L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_7, 
         L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_6, 
         L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_5, 
         L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_4, 
         L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_3, 
         L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_2, 
         L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_1, 
         L1_3_L2_0_G2_MINI_ALU_BoothP_16, L1_3_L2_0_G2_MINI_ALU_BoothP_15, 
         L1_3_L2_0_G2_MINI_ALU_BoothP_14, L1_3_L2_0_G2_MINI_ALU_BoothP_13, 
         L1_3_L2_0_G2_MINI_ALU_BoothP_12, L1_3_L2_0_G2_MINI_ALU_BoothP_11, 
         L1_3_L2_0_G2_MINI_ALU_BoothP_10, L1_3_L2_0_G2_MINI_ALU_BoothP_9, 
         L1_3_L2_0_G2_MINI_ALU_BoothP_8, L1_3_L2_0_G2_MINI_ALU_BoothP_7, 
         L1_3_L2_0_G2_MINI_ALU_BoothP_6, L1_3_L2_0_G2_MINI_ALU_BoothP_5, 
         L1_3_L2_0_G2_MINI_ALU_BoothP_4, L1_3_L2_0_G2_MINI_ALU_BoothP_3, 
         L1_3_L2_0_G2_MINI_ALU_BoothP_2, L1_3_L2_0_G2_MINI_ALU_BoothP_1, 
         L1_3_L2_0_G2_MINI_ALU_BoothP_0, L1_3_L2_0_G2_MINI_ALU_nx0, 
         L1_3_L2_0_G2_MINI_ALU_nx6, L1_3_L2_0_G2_MINI_ALU_nx12, 
         L1_3_L2_0_G2_MINI_ALU_nx18, L1_3_L2_0_G2_MINI_ALU_nx24, 
         L1_3_L2_0_G2_MINI_ALU_nx30, L1_3_L2_0_G2_MINI_ALU_nx40, 
         L1_3_L2_0_G2_MINI_ALU_nx44, L1_3_L2_0_G2_MINI_ALU_nx48, 
         L1_3_L2_0_G2_MINI_ALU_nx52, L1_3_L2_0_G2_MINI_ALU_nx56, 
         L1_3_L2_0_G2_MINI_ALU_nx62, L1_3_L2_0_G2_MINI_ALU_nx154, 
         L1_3_L2_0_G2_MINI_ALU_nx316, L1_3_L2_0_G2_MINI_ALU_nx336, 
         L1_3_L2_0_G2_MINI_ALU_nx356, L1_3_L2_0_G2_MINI_ALU_nx376, 
         L1_3_L2_0_G2_MINI_ALU_nx396, L1_3_L2_0_G2_MINI_ALU_nx416, 
         L1_3_L2_0_G2_MINI_ALU_nx436, L1_3_L2_0_G2_MINI_ALU_nx454, 
         L1_3_L2_0_G2_MINI_ALU_nx456, L1_3_L2_0_G2_MINI_ALU_nx379, 
         L1_3_L2_0_G2_MINI_ALU_nx381, L1_3_L2_0_G2_MINI_ALU_nx383, 
         L1_3_L2_0_G2_MINI_ALU_nx387, L1_3_L2_0_G2_MINI_ALU_nx389, 
         L1_3_L2_0_G2_MINI_ALU_nx391, L1_3_L2_0_G2_MINI_ALU_nx395, 
         L1_3_L2_0_G2_MINI_ALU_nx399, L1_3_L2_0_G2_MINI_ALU_nx401, 
         L1_3_L2_0_G2_MINI_ALU_nx403, L1_3_L2_0_G2_MINI_ALU_nx405, 
         L1_3_L2_0_G2_MINI_ALU_nx409, L1_3_L2_0_G2_MINI_ALU_nx411, 
         L1_3_L2_0_G2_MINI_ALU_nx413, L1_3_L2_0_G2_MINI_ALU_nx415, 
         L1_3_L2_0_G2_MINI_ALU_nx419, L1_3_L2_0_G2_MINI_ALU_nx421, 
         L1_3_L2_0_G2_MINI_ALU_nx423, L1_3_L2_0_G2_MINI_ALU_nx425, 
         L1_3_L2_0_G2_MINI_ALU_nx429, L1_3_L2_0_G2_MINI_ALU_nx431, 
         L1_3_L2_0_G2_MINI_ALU_nx433, L1_3_L2_0_G2_MINI_ALU_nx435, 
         L1_3_L2_0_G2_MINI_ALU_nx439, L1_3_L2_0_G2_MINI_ALU_nx441, 
         L1_3_L2_0_G2_MINI_ALU_nx443, L1_3_L2_0_G2_MINI_ALU_nx445, 
         L1_3_L2_0_G2_MINI_ALU_nx449, L1_3_L2_0_G2_MINI_ALU_nx451, 
         L1_3_L2_0_G2_MINI_ALU_nx453, L1_3_L2_0_G2_MINI_ALU_nx455, 
         L1_3_L2_0_G2_MINI_ALU_nx461, L1_3_L2_0_G2_MINI_ALU_nx463, 
         L1_3_L2_0_G2_MINI_ALU_nx467, L1_3_L2_0_G2_MINI_ALU_nx469, 
         L1_3_L2_0_G2_MINI_ALU_nx471, L1_3_L2_0_G2_MINI_ALU_nx475, 
         L1_3_L2_0_G2_MINI_ALU_nx477, L1_3_L2_0_G2_MINI_ALU_nx479, 
         L1_3_L2_0_G2_MINI_ALU_nx483, L1_3_L2_0_G2_MINI_ALU_nx485, 
         L1_3_L2_0_G2_MINI_ALU_nx487, L1_3_L2_0_G2_MINI_ALU_nx491, 
         L1_3_L2_0_G2_MINI_ALU_nx493, L1_3_L2_0_G2_MINI_ALU_nx495, 
         L1_3_L2_0_G2_MINI_ALU_nx499, L1_3_L2_0_G2_MINI_ALU_nx501, 
         L1_3_L2_0_G2_MINI_ALU_nx503, L1_3_L2_0_G2_MINI_ALU_nx507, 
         L1_3_L2_0_G2_MINI_ALU_nx509, L1_3_L2_0_G2_MINI_ALU_nx511, 
         L1_3_L2_0_G2_MINI_ALU_nx515, L1_3_L2_0_G2_MINI_ALU_nx517, 
         L1_3_L2_0_G2_MINI_ALU_nx529, L1_3_L2_0_G2_MINI_ALU_nx531, 
         L1_3_L2_0_G2_MINI_ALU_nx534, L1_3_L2_0_G2_MINI_ALU_nx537, 
         L1_3_L2_0_G2_MINI_ALU_nx540, L1_3_L2_0_G2_MINI_ALU_nx544, 
         L1_3_L2_0_G2_MINI_ALU_nx547, L1_3_L2_0_G2_MINI_ALU_nx551, 
         L1_3_L2_0_G2_MINI_ALU_nx554, L1_3_L2_0_G2_MINI_ALU_nx558, 
         L1_3_L2_0_G2_MINI_ALU_nx561, L1_3_L2_0_G2_MINI_ALU_nx565, 
         L1_3_L2_0_G2_MINI_ALU_nx568, 
         L1_3_L2_0_G2_MINI_ALU_WindowCellShiftedLeft_16, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_16, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_15, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_14, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_13, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_12, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_11, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_10, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_16, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_15, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_14, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_13, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_12, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_11, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_10, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_9, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_8, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_7, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_6, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_5, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_4, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_3, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_2, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_1, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_0, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_16, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_15, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_14, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_13, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_12, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_11, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_10, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_9, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_8, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_7, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_6, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_5, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_4, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_3, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_2, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_1, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_0, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_16, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_15, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_14, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_13, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_12, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_11, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_10, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_9, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_8, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_7, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_6, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_5, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_4, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_3, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_2, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_1, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_0, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_nx4, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_nx8, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_nx12, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_nx16, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_nx20, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_nx24, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_nx80, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_nx328, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_nx384, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642, 
         L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644, 
         L1_3_L2_1_G2_MINI_ALU_AddPToBoothOperand, 
         L1_3_L2_1_G2_MINI_ALU_BoothOperand_16, 
         L1_3_L2_1_G2_MINI_ALU_BoothOperand_15, 
         L1_3_L2_1_G2_MINI_ALU_BoothOperand_14, 
         L1_3_L2_1_G2_MINI_ALU_BoothOperand_13, 
         L1_3_L2_1_G2_MINI_ALU_BoothOperand_12, 
         L1_3_L2_1_G2_MINI_ALU_BoothOperand_11, 
         L1_3_L2_1_G2_MINI_ALU_BoothOperand_10, 
         L1_3_L2_1_G2_MINI_ALU_BoothOperand_9, 
         L1_3_L2_1_G2_MINI_ALU_BoothOperand_8, 
         L1_3_L2_1_G2_MINI_ALU_BoothOperand_7, 
         L1_3_L2_1_G2_MINI_ALU_BoothOperand_6, 
         L1_3_L2_1_G2_MINI_ALU_BoothOperand_5, 
         L1_3_L2_1_G2_MINI_ALU_BoothOperand_4, 
         L1_3_L2_1_G2_MINI_ALU_BoothOperand_3, 
         L1_3_L2_1_G2_MINI_ALU_BoothOperand_2, 
         L1_3_L2_1_G2_MINI_ALU_BoothOperand_1, 
         L1_3_L2_1_G2_MINI_ALU_BoothOperand_0, 
         L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_16, 
         L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_15, 
         L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_14, 
         L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_13, 
         L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_12, 
         L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_11, 
         L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_10, 
         L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_9, 
         L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_8, 
         L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_7, 
         L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_6, 
         L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_5, 
         L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_4, 
         L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_3, 
         L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_2, 
         L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_1, 
         L1_3_L2_1_G2_MINI_ALU_BoothP_16, L1_3_L2_1_G2_MINI_ALU_BoothP_15, 
         L1_3_L2_1_G2_MINI_ALU_BoothP_14, L1_3_L2_1_G2_MINI_ALU_BoothP_13, 
         L1_3_L2_1_G2_MINI_ALU_BoothP_12, L1_3_L2_1_G2_MINI_ALU_BoothP_11, 
         L1_3_L2_1_G2_MINI_ALU_BoothP_10, L1_3_L2_1_G2_MINI_ALU_BoothP_9, 
         L1_3_L2_1_G2_MINI_ALU_BoothP_8, L1_3_L2_1_G2_MINI_ALU_BoothP_7, 
         L1_3_L2_1_G2_MINI_ALU_BoothP_6, L1_3_L2_1_G2_MINI_ALU_BoothP_5, 
         L1_3_L2_1_G2_MINI_ALU_BoothP_4, L1_3_L2_1_G2_MINI_ALU_BoothP_3, 
         L1_3_L2_1_G2_MINI_ALU_BoothP_2, L1_3_L2_1_G2_MINI_ALU_BoothP_1, 
         L1_3_L2_1_G2_MINI_ALU_BoothP_0, L1_3_L2_1_G2_MINI_ALU_nx0, 
         L1_3_L2_1_G2_MINI_ALU_nx6, L1_3_L2_1_G2_MINI_ALU_nx12, 
         L1_3_L2_1_G2_MINI_ALU_nx18, L1_3_L2_1_G2_MINI_ALU_nx24, 
         L1_3_L2_1_G2_MINI_ALU_nx30, L1_3_L2_1_G2_MINI_ALU_nx40, 
         L1_3_L2_1_G2_MINI_ALU_nx44, L1_3_L2_1_G2_MINI_ALU_nx48, 
         L1_3_L2_1_G2_MINI_ALU_nx52, L1_3_L2_1_G2_MINI_ALU_nx56, 
         L1_3_L2_1_G2_MINI_ALU_nx62, L1_3_L2_1_G2_MINI_ALU_nx154, 
         L1_3_L2_1_G2_MINI_ALU_nx316, L1_3_L2_1_G2_MINI_ALU_nx336, 
         L1_3_L2_1_G2_MINI_ALU_nx356, L1_3_L2_1_G2_MINI_ALU_nx376, 
         L1_3_L2_1_G2_MINI_ALU_nx396, L1_3_L2_1_G2_MINI_ALU_nx416, 
         L1_3_L2_1_G2_MINI_ALU_nx436, L1_3_L2_1_G2_MINI_ALU_nx454, 
         L1_3_L2_1_G2_MINI_ALU_nx456, L1_3_L2_1_G2_MINI_ALU_nx379, 
         L1_3_L2_1_G2_MINI_ALU_nx381, L1_3_L2_1_G2_MINI_ALU_nx383, 
         L1_3_L2_1_G2_MINI_ALU_nx387, L1_3_L2_1_G2_MINI_ALU_nx389, 
         L1_3_L2_1_G2_MINI_ALU_nx391, L1_3_L2_1_G2_MINI_ALU_nx395, 
         L1_3_L2_1_G2_MINI_ALU_nx399, L1_3_L2_1_G2_MINI_ALU_nx401, 
         L1_3_L2_1_G2_MINI_ALU_nx403, L1_3_L2_1_G2_MINI_ALU_nx405, 
         L1_3_L2_1_G2_MINI_ALU_nx409, L1_3_L2_1_G2_MINI_ALU_nx411, 
         L1_3_L2_1_G2_MINI_ALU_nx413, L1_3_L2_1_G2_MINI_ALU_nx415, 
         L1_3_L2_1_G2_MINI_ALU_nx419, L1_3_L2_1_G2_MINI_ALU_nx421, 
         L1_3_L2_1_G2_MINI_ALU_nx423, L1_3_L2_1_G2_MINI_ALU_nx425, 
         L1_3_L2_1_G2_MINI_ALU_nx429, L1_3_L2_1_G2_MINI_ALU_nx431, 
         L1_3_L2_1_G2_MINI_ALU_nx433, L1_3_L2_1_G2_MINI_ALU_nx435, 
         L1_3_L2_1_G2_MINI_ALU_nx439, L1_3_L2_1_G2_MINI_ALU_nx441, 
         L1_3_L2_1_G2_MINI_ALU_nx443, L1_3_L2_1_G2_MINI_ALU_nx445, 
         L1_3_L2_1_G2_MINI_ALU_nx449, L1_3_L2_1_G2_MINI_ALU_nx451, 
         L1_3_L2_1_G2_MINI_ALU_nx453, L1_3_L2_1_G2_MINI_ALU_nx455, 
         L1_3_L2_1_G2_MINI_ALU_nx461, L1_3_L2_1_G2_MINI_ALU_nx463, 
         L1_3_L2_1_G2_MINI_ALU_nx467, L1_3_L2_1_G2_MINI_ALU_nx469, 
         L1_3_L2_1_G2_MINI_ALU_nx471, L1_3_L2_1_G2_MINI_ALU_nx475, 
         L1_3_L2_1_G2_MINI_ALU_nx477, L1_3_L2_1_G2_MINI_ALU_nx479, 
         L1_3_L2_1_G2_MINI_ALU_nx483, L1_3_L2_1_G2_MINI_ALU_nx485, 
         L1_3_L2_1_G2_MINI_ALU_nx487, L1_3_L2_1_G2_MINI_ALU_nx491, 
         L1_3_L2_1_G2_MINI_ALU_nx493, L1_3_L2_1_G2_MINI_ALU_nx495, 
         L1_3_L2_1_G2_MINI_ALU_nx499, L1_3_L2_1_G2_MINI_ALU_nx501, 
         L1_3_L2_1_G2_MINI_ALU_nx503, L1_3_L2_1_G2_MINI_ALU_nx507, 
         L1_3_L2_1_G2_MINI_ALU_nx509, L1_3_L2_1_G2_MINI_ALU_nx511, 
         L1_3_L2_1_G2_MINI_ALU_nx515, L1_3_L2_1_G2_MINI_ALU_nx517, 
         L1_3_L2_1_G2_MINI_ALU_nx529, L1_3_L2_1_G2_MINI_ALU_nx531, 
         L1_3_L2_1_G2_MINI_ALU_nx534, L1_3_L2_1_G2_MINI_ALU_nx537, 
         L1_3_L2_1_G2_MINI_ALU_nx540, L1_3_L2_1_G2_MINI_ALU_nx544, 
         L1_3_L2_1_G2_MINI_ALU_nx547, L1_3_L2_1_G2_MINI_ALU_nx551, 
         L1_3_L2_1_G2_MINI_ALU_nx554, L1_3_L2_1_G2_MINI_ALU_nx558, 
         L1_3_L2_1_G2_MINI_ALU_nx561, L1_3_L2_1_G2_MINI_ALU_nx565, 
         L1_3_L2_1_G2_MINI_ALU_nx568, 
         L1_3_L2_1_G2_MINI_ALU_WindowCellShiftedLeft_16, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_16, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_15, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_14, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_13, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_12, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_11, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_10, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_16, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_15, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_14, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_13, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_12, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_11, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_10, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_9, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_8, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_7, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_6, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_5, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_4, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_3, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_2, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_1, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_0, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_16, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_15, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_14, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_13, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_12, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_11, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_10, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_9, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_8, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_7, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_6, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_5, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_4, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_3, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_2, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_1, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_0, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_16, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_15, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_14, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_13, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_12, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_11, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_10, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_9, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_8, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_7, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_6, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_5, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_4, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_3, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_2, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_1, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_0, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_nx4, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_nx8, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_nx12, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_nx16, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_nx20, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_nx24, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_nx80, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_nx328, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_nx384, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642, 
         L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644, 
         L1_3_L2_2_G2_MINI_ALU_AddPToBoothOperand, 
         L1_3_L2_2_G2_MINI_ALU_BoothOperand_16, 
         L1_3_L2_2_G2_MINI_ALU_BoothOperand_15, 
         L1_3_L2_2_G2_MINI_ALU_BoothOperand_14, 
         L1_3_L2_2_G2_MINI_ALU_BoothOperand_13, 
         L1_3_L2_2_G2_MINI_ALU_BoothOperand_12, 
         L1_3_L2_2_G2_MINI_ALU_BoothOperand_11, 
         L1_3_L2_2_G2_MINI_ALU_BoothOperand_10, 
         L1_3_L2_2_G2_MINI_ALU_BoothOperand_9, 
         L1_3_L2_2_G2_MINI_ALU_BoothOperand_8, 
         L1_3_L2_2_G2_MINI_ALU_BoothOperand_7, 
         L1_3_L2_2_G2_MINI_ALU_BoothOperand_6, 
         L1_3_L2_2_G2_MINI_ALU_BoothOperand_5, 
         L1_3_L2_2_G2_MINI_ALU_BoothOperand_4, 
         L1_3_L2_2_G2_MINI_ALU_BoothOperand_3, 
         L1_3_L2_2_G2_MINI_ALU_BoothOperand_2, 
         L1_3_L2_2_G2_MINI_ALU_BoothOperand_1, 
         L1_3_L2_2_G2_MINI_ALU_BoothOperand_0, 
         L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_16, 
         L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_15, 
         L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_14, 
         L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_13, 
         L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_12, 
         L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_11, 
         L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_10, 
         L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_9, 
         L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_8, 
         L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_7, 
         L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_6, 
         L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_5, 
         L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_4, 
         L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_3, 
         L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_2, 
         L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_1, 
         L1_3_L2_2_G2_MINI_ALU_BoothP_16, L1_3_L2_2_G2_MINI_ALU_BoothP_15, 
         L1_3_L2_2_G2_MINI_ALU_BoothP_14, L1_3_L2_2_G2_MINI_ALU_BoothP_13, 
         L1_3_L2_2_G2_MINI_ALU_BoothP_12, L1_3_L2_2_G2_MINI_ALU_BoothP_11, 
         L1_3_L2_2_G2_MINI_ALU_BoothP_10, L1_3_L2_2_G2_MINI_ALU_BoothP_9, 
         L1_3_L2_2_G2_MINI_ALU_BoothP_8, L1_3_L2_2_G2_MINI_ALU_BoothP_7, 
         L1_3_L2_2_G2_MINI_ALU_BoothP_6, L1_3_L2_2_G2_MINI_ALU_BoothP_5, 
         L1_3_L2_2_G2_MINI_ALU_BoothP_4, L1_3_L2_2_G2_MINI_ALU_BoothP_3, 
         L1_3_L2_2_G2_MINI_ALU_BoothP_2, L1_3_L2_2_G2_MINI_ALU_BoothP_1, 
         L1_3_L2_2_G2_MINI_ALU_BoothP_0, L1_3_L2_2_G2_MINI_ALU_nx0, 
         L1_3_L2_2_G2_MINI_ALU_nx6, L1_3_L2_2_G2_MINI_ALU_nx12, 
         L1_3_L2_2_G2_MINI_ALU_nx18, L1_3_L2_2_G2_MINI_ALU_nx24, 
         L1_3_L2_2_G2_MINI_ALU_nx30, L1_3_L2_2_G2_MINI_ALU_nx40, 
         L1_3_L2_2_G2_MINI_ALU_nx44, L1_3_L2_2_G2_MINI_ALU_nx48, 
         L1_3_L2_2_G2_MINI_ALU_nx52, L1_3_L2_2_G2_MINI_ALU_nx56, 
         L1_3_L2_2_G2_MINI_ALU_nx62, L1_3_L2_2_G2_MINI_ALU_nx154, 
         L1_3_L2_2_G2_MINI_ALU_nx316, L1_3_L2_2_G2_MINI_ALU_nx336, 
         L1_3_L2_2_G2_MINI_ALU_nx356, L1_3_L2_2_G2_MINI_ALU_nx376, 
         L1_3_L2_2_G2_MINI_ALU_nx396, L1_3_L2_2_G2_MINI_ALU_nx416, 
         L1_3_L2_2_G2_MINI_ALU_nx436, L1_3_L2_2_G2_MINI_ALU_nx454, 
         L1_3_L2_2_G2_MINI_ALU_nx456, L1_3_L2_2_G2_MINI_ALU_nx379, 
         L1_3_L2_2_G2_MINI_ALU_nx381, L1_3_L2_2_G2_MINI_ALU_nx383, 
         L1_3_L2_2_G2_MINI_ALU_nx387, L1_3_L2_2_G2_MINI_ALU_nx389, 
         L1_3_L2_2_G2_MINI_ALU_nx391, L1_3_L2_2_G2_MINI_ALU_nx395, 
         L1_3_L2_2_G2_MINI_ALU_nx399, L1_3_L2_2_G2_MINI_ALU_nx401, 
         L1_3_L2_2_G2_MINI_ALU_nx403, L1_3_L2_2_G2_MINI_ALU_nx405, 
         L1_3_L2_2_G2_MINI_ALU_nx409, L1_3_L2_2_G2_MINI_ALU_nx411, 
         L1_3_L2_2_G2_MINI_ALU_nx413, L1_3_L2_2_G2_MINI_ALU_nx415, 
         L1_3_L2_2_G2_MINI_ALU_nx419, L1_3_L2_2_G2_MINI_ALU_nx421, 
         L1_3_L2_2_G2_MINI_ALU_nx423, L1_3_L2_2_G2_MINI_ALU_nx425, 
         L1_3_L2_2_G2_MINI_ALU_nx429, L1_3_L2_2_G2_MINI_ALU_nx431, 
         L1_3_L2_2_G2_MINI_ALU_nx433, L1_3_L2_2_G2_MINI_ALU_nx435, 
         L1_3_L2_2_G2_MINI_ALU_nx439, L1_3_L2_2_G2_MINI_ALU_nx441, 
         L1_3_L2_2_G2_MINI_ALU_nx443, L1_3_L2_2_G2_MINI_ALU_nx445, 
         L1_3_L2_2_G2_MINI_ALU_nx449, L1_3_L2_2_G2_MINI_ALU_nx451, 
         L1_3_L2_2_G2_MINI_ALU_nx453, L1_3_L2_2_G2_MINI_ALU_nx455, 
         L1_3_L2_2_G2_MINI_ALU_nx461, L1_3_L2_2_G2_MINI_ALU_nx463, 
         L1_3_L2_2_G2_MINI_ALU_nx467, L1_3_L2_2_G2_MINI_ALU_nx469, 
         L1_3_L2_2_G2_MINI_ALU_nx471, L1_3_L2_2_G2_MINI_ALU_nx475, 
         L1_3_L2_2_G2_MINI_ALU_nx477, L1_3_L2_2_G2_MINI_ALU_nx479, 
         L1_3_L2_2_G2_MINI_ALU_nx483, L1_3_L2_2_G2_MINI_ALU_nx485, 
         L1_3_L2_2_G2_MINI_ALU_nx487, L1_3_L2_2_G2_MINI_ALU_nx491, 
         L1_3_L2_2_G2_MINI_ALU_nx493, L1_3_L2_2_G2_MINI_ALU_nx495, 
         L1_3_L2_2_G2_MINI_ALU_nx499, L1_3_L2_2_G2_MINI_ALU_nx501, 
         L1_3_L2_2_G2_MINI_ALU_nx503, L1_3_L2_2_G2_MINI_ALU_nx507, 
         L1_3_L2_2_G2_MINI_ALU_nx509, L1_3_L2_2_G2_MINI_ALU_nx511, 
         L1_3_L2_2_G2_MINI_ALU_nx515, L1_3_L2_2_G2_MINI_ALU_nx517, 
         L1_3_L2_2_G2_MINI_ALU_nx529, L1_3_L2_2_G2_MINI_ALU_nx531, 
         L1_3_L2_2_G2_MINI_ALU_nx534, L1_3_L2_2_G2_MINI_ALU_nx537, 
         L1_3_L2_2_G2_MINI_ALU_nx540, L1_3_L2_2_G2_MINI_ALU_nx544, 
         L1_3_L2_2_G2_MINI_ALU_nx547, L1_3_L2_2_G2_MINI_ALU_nx551, 
         L1_3_L2_2_G2_MINI_ALU_nx554, L1_3_L2_2_G2_MINI_ALU_nx558, 
         L1_3_L2_2_G2_MINI_ALU_nx561, L1_3_L2_2_G2_MINI_ALU_nx565, 
         L1_3_L2_2_G2_MINI_ALU_nx568, 
         L1_3_L2_2_G2_MINI_ALU_WindowCellShiftedLeft_16, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_16, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_15, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_14, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_13, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_12, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_11, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_10, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_16, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_15, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_14, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_13, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_12, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_11, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_10, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_9, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_8, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_7, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_6, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_5, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_4, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_3, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_2, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_1, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_0, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_16, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_15, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_14, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_13, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_12, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_11, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_10, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_9, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_8, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_7, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_6, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_5, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_4, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_3, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_2, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_1, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_0, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_16, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_15, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_14, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_13, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_12, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_11, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_10, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_9, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_8, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_7, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_6, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_5, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_4, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_3, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_2, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_1, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_0, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_nx4, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_nx8, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_nx12, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_nx16, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_nx20, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_nx24, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_nx80, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_nx328, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_nx384, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642, 
         L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644, 
         L1_3_L2_3_G2_MINI_ALU_AddPToBoothOperand, 
         L1_3_L2_3_G2_MINI_ALU_BoothOperand_16, 
         L1_3_L2_3_G2_MINI_ALU_BoothOperand_15, 
         L1_3_L2_3_G2_MINI_ALU_BoothOperand_14, 
         L1_3_L2_3_G2_MINI_ALU_BoothOperand_13, 
         L1_3_L2_3_G2_MINI_ALU_BoothOperand_12, 
         L1_3_L2_3_G2_MINI_ALU_BoothOperand_11, 
         L1_3_L2_3_G2_MINI_ALU_BoothOperand_10, 
         L1_3_L2_3_G2_MINI_ALU_BoothOperand_9, 
         L1_3_L2_3_G2_MINI_ALU_BoothOperand_8, 
         L1_3_L2_3_G2_MINI_ALU_BoothOperand_7, 
         L1_3_L2_3_G2_MINI_ALU_BoothOperand_6, 
         L1_3_L2_3_G2_MINI_ALU_BoothOperand_5, 
         L1_3_L2_3_G2_MINI_ALU_BoothOperand_4, 
         L1_3_L2_3_G2_MINI_ALU_BoothOperand_3, 
         L1_3_L2_3_G2_MINI_ALU_BoothOperand_2, 
         L1_3_L2_3_G2_MINI_ALU_BoothOperand_1, 
         L1_3_L2_3_G2_MINI_ALU_BoothOperand_0, 
         L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_16, 
         L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_15, 
         L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_14, 
         L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_13, 
         L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_12, 
         L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_11, 
         L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_10, 
         L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_9, 
         L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_8, 
         L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_7, 
         L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_6, 
         L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_5, 
         L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_4, 
         L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_3, 
         L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_2, 
         L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_1, 
         L1_3_L2_3_G2_MINI_ALU_BoothP_16, L1_3_L2_3_G2_MINI_ALU_BoothP_15, 
         L1_3_L2_3_G2_MINI_ALU_BoothP_14, L1_3_L2_3_G2_MINI_ALU_BoothP_13, 
         L1_3_L2_3_G2_MINI_ALU_BoothP_12, L1_3_L2_3_G2_MINI_ALU_BoothP_11, 
         L1_3_L2_3_G2_MINI_ALU_BoothP_10, L1_3_L2_3_G2_MINI_ALU_BoothP_9, 
         L1_3_L2_3_G2_MINI_ALU_BoothP_8, L1_3_L2_3_G2_MINI_ALU_BoothP_7, 
         L1_3_L2_3_G2_MINI_ALU_BoothP_6, L1_3_L2_3_G2_MINI_ALU_BoothP_5, 
         L1_3_L2_3_G2_MINI_ALU_BoothP_4, L1_3_L2_3_G2_MINI_ALU_BoothP_3, 
         L1_3_L2_3_G2_MINI_ALU_BoothP_2, L1_3_L2_3_G2_MINI_ALU_BoothP_1, 
         L1_3_L2_3_G2_MINI_ALU_BoothP_0, L1_3_L2_3_G2_MINI_ALU_nx0, 
         L1_3_L2_3_G2_MINI_ALU_nx6, L1_3_L2_3_G2_MINI_ALU_nx12, 
         L1_3_L2_3_G2_MINI_ALU_nx18, L1_3_L2_3_G2_MINI_ALU_nx24, 
         L1_3_L2_3_G2_MINI_ALU_nx30, L1_3_L2_3_G2_MINI_ALU_nx40, 
         L1_3_L2_3_G2_MINI_ALU_nx44, L1_3_L2_3_G2_MINI_ALU_nx48, 
         L1_3_L2_3_G2_MINI_ALU_nx52, L1_3_L2_3_G2_MINI_ALU_nx56, 
         L1_3_L2_3_G2_MINI_ALU_nx62, L1_3_L2_3_G2_MINI_ALU_nx154, 
         L1_3_L2_3_G2_MINI_ALU_nx316, L1_3_L2_3_G2_MINI_ALU_nx336, 
         L1_3_L2_3_G2_MINI_ALU_nx356, L1_3_L2_3_G2_MINI_ALU_nx376, 
         L1_3_L2_3_G2_MINI_ALU_nx396, L1_3_L2_3_G2_MINI_ALU_nx416, 
         L1_3_L2_3_G2_MINI_ALU_nx436, L1_3_L2_3_G2_MINI_ALU_nx454, 
         L1_3_L2_3_G2_MINI_ALU_nx456, L1_3_L2_3_G2_MINI_ALU_nx379, 
         L1_3_L2_3_G2_MINI_ALU_nx381, L1_3_L2_3_G2_MINI_ALU_nx383, 
         L1_3_L2_3_G2_MINI_ALU_nx387, L1_3_L2_3_G2_MINI_ALU_nx389, 
         L1_3_L2_3_G2_MINI_ALU_nx391, L1_3_L2_3_G2_MINI_ALU_nx395, 
         L1_3_L2_3_G2_MINI_ALU_nx399, L1_3_L2_3_G2_MINI_ALU_nx401, 
         L1_3_L2_3_G2_MINI_ALU_nx403, L1_3_L2_3_G2_MINI_ALU_nx405, 
         L1_3_L2_3_G2_MINI_ALU_nx409, L1_3_L2_3_G2_MINI_ALU_nx411, 
         L1_3_L2_3_G2_MINI_ALU_nx413, L1_3_L2_3_G2_MINI_ALU_nx415, 
         L1_3_L2_3_G2_MINI_ALU_nx419, L1_3_L2_3_G2_MINI_ALU_nx421, 
         L1_3_L2_3_G2_MINI_ALU_nx423, L1_3_L2_3_G2_MINI_ALU_nx425, 
         L1_3_L2_3_G2_MINI_ALU_nx429, L1_3_L2_3_G2_MINI_ALU_nx431, 
         L1_3_L2_3_G2_MINI_ALU_nx433, L1_3_L2_3_G2_MINI_ALU_nx435, 
         L1_3_L2_3_G2_MINI_ALU_nx439, L1_3_L2_3_G2_MINI_ALU_nx441, 
         L1_3_L2_3_G2_MINI_ALU_nx443, L1_3_L2_3_G2_MINI_ALU_nx445, 
         L1_3_L2_3_G2_MINI_ALU_nx449, L1_3_L2_3_G2_MINI_ALU_nx451, 
         L1_3_L2_3_G2_MINI_ALU_nx453, L1_3_L2_3_G2_MINI_ALU_nx455, 
         L1_3_L2_3_G2_MINI_ALU_nx461, L1_3_L2_3_G2_MINI_ALU_nx463, 
         L1_3_L2_3_G2_MINI_ALU_nx467, L1_3_L2_3_G2_MINI_ALU_nx469, 
         L1_3_L2_3_G2_MINI_ALU_nx471, L1_3_L2_3_G2_MINI_ALU_nx475, 
         L1_3_L2_3_G2_MINI_ALU_nx477, L1_3_L2_3_G2_MINI_ALU_nx479, 
         L1_3_L2_3_G2_MINI_ALU_nx483, L1_3_L2_3_G2_MINI_ALU_nx485, 
         L1_3_L2_3_G2_MINI_ALU_nx487, L1_3_L2_3_G2_MINI_ALU_nx491, 
         L1_3_L2_3_G2_MINI_ALU_nx493, L1_3_L2_3_G2_MINI_ALU_nx495, 
         L1_3_L2_3_G2_MINI_ALU_nx499, L1_3_L2_3_G2_MINI_ALU_nx501, 
         L1_3_L2_3_G2_MINI_ALU_nx503, L1_3_L2_3_G2_MINI_ALU_nx507, 
         L1_3_L2_3_G2_MINI_ALU_nx509, L1_3_L2_3_G2_MINI_ALU_nx511, 
         L1_3_L2_3_G2_MINI_ALU_nx515, L1_3_L2_3_G2_MINI_ALU_nx517, 
         L1_3_L2_3_G2_MINI_ALU_nx529, L1_3_L2_3_G2_MINI_ALU_nx531, 
         L1_3_L2_3_G2_MINI_ALU_nx534, L1_3_L2_3_G2_MINI_ALU_nx537, 
         L1_3_L2_3_G2_MINI_ALU_nx540, L1_3_L2_3_G2_MINI_ALU_nx544, 
         L1_3_L2_3_G2_MINI_ALU_nx547, L1_3_L2_3_G2_MINI_ALU_nx551, 
         L1_3_L2_3_G2_MINI_ALU_nx554, L1_3_L2_3_G2_MINI_ALU_nx558, 
         L1_3_L2_3_G2_MINI_ALU_nx561, L1_3_L2_3_G2_MINI_ALU_nx565, 
         L1_3_L2_3_G2_MINI_ALU_nx568, 
         L1_3_L2_3_G2_MINI_ALU_WindowCellShiftedLeft_16, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_16, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_15, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_14, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_13, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_12, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_11, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_10, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_16, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_15, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_14, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_13, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_12, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_11, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_10, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_9, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_8, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_7, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_6, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_5, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_4, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_3, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_2, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_1, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_0, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_16, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_15, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_14, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_13, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_12, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_11, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_10, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_9, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_8, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_7, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_6, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_5, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_4, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_3, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_2, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_1, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_0, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_16, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_15, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_14, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_13, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_12, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_11, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_10, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_9, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_8, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_7, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_6, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_5, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_4, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_3, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_2, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_1, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_0, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx4, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx8, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx12, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx16, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx20, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx24, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx80, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx328, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx384, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642, 
         L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644, 
         L1_3_L2_4_G3_MINI_ALU_AddPToBoothOperand, 
         L1_3_L2_4_G3_MINI_ALU_BoothOperand_16, 
         L1_3_L2_4_G3_MINI_ALU_BoothOperand_15, 
         L1_3_L2_4_G3_MINI_ALU_BoothOperand_14, 
         L1_3_L2_4_G3_MINI_ALU_BoothOperand_13, 
         L1_3_L2_4_G3_MINI_ALU_BoothOperand_12, 
         L1_3_L2_4_G3_MINI_ALU_BoothOperand_11, 
         L1_3_L2_4_G3_MINI_ALU_BoothOperand_10, 
         L1_3_L2_4_G3_MINI_ALU_BoothOperand_9, 
         L1_3_L2_4_G3_MINI_ALU_BoothOperand_8, 
         L1_3_L2_4_G3_MINI_ALU_BoothOperand_7, 
         L1_3_L2_4_G3_MINI_ALU_BoothOperand_6, 
         L1_3_L2_4_G3_MINI_ALU_BoothOperand_5, 
         L1_3_L2_4_G3_MINI_ALU_BoothOperand_4, 
         L1_3_L2_4_G3_MINI_ALU_BoothOperand_3, 
         L1_3_L2_4_G3_MINI_ALU_BoothOperand_2, 
         L1_3_L2_4_G3_MINI_ALU_BoothOperand_1, 
         L1_3_L2_4_G3_MINI_ALU_BoothOperand_0, 
         L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_16, 
         L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_15, 
         L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_14, 
         L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_13, 
         L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_12, 
         L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_11, 
         L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_10, 
         L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_9, 
         L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_8, 
         L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_7, 
         L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_6, 
         L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_5, 
         L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_4, 
         L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_3, 
         L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_2, 
         L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_1, 
         L1_3_L2_4_G3_MINI_ALU_BoothP_16, L1_3_L2_4_G3_MINI_ALU_BoothP_15, 
         L1_3_L2_4_G3_MINI_ALU_BoothP_14, L1_3_L2_4_G3_MINI_ALU_BoothP_13, 
         L1_3_L2_4_G3_MINI_ALU_BoothP_12, L1_3_L2_4_G3_MINI_ALU_BoothP_11, 
         L1_3_L2_4_G3_MINI_ALU_BoothP_10, L1_3_L2_4_G3_MINI_ALU_BoothP_9, 
         L1_3_L2_4_G3_MINI_ALU_BoothP_8, L1_3_L2_4_G3_MINI_ALU_BoothP_7, 
         L1_3_L2_4_G3_MINI_ALU_BoothP_6, L1_3_L2_4_G3_MINI_ALU_BoothP_5, 
         L1_3_L2_4_G3_MINI_ALU_BoothP_4, L1_3_L2_4_G3_MINI_ALU_BoothP_3, 
         L1_3_L2_4_G3_MINI_ALU_BoothP_2, L1_3_L2_4_G3_MINI_ALU_BoothP_1, 
         L1_3_L2_4_G3_MINI_ALU_BoothP_0, L1_3_L2_4_G3_MINI_ALU_nx0, 
         L1_3_L2_4_G3_MINI_ALU_nx6, L1_3_L2_4_G3_MINI_ALU_nx12, 
         L1_3_L2_4_G3_MINI_ALU_nx18, L1_3_L2_4_G3_MINI_ALU_nx24, 
         L1_3_L2_4_G3_MINI_ALU_nx30, L1_3_L2_4_G3_MINI_ALU_nx40, 
         L1_3_L2_4_G3_MINI_ALU_nx44, L1_3_L2_4_G3_MINI_ALU_nx48, 
         L1_3_L2_4_G3_MINI_ALU_nx52, L1_3_L2_4_G3_MINI_ALU_nx56, 
         L1_3_L2_4_G3_MINI_ALU_nx62, L1_3_L2_4_G3_MINI_ALU_nx154, 
         L1_3_L2_4_G3_MINI_ALU_nx316, L1_3_L2_4_G3_MINI_ALU_nx336, 
         L1_3_L2_4_G3_MINI_ALU_nx356, L1_3_L2_4_G3_MINI_ALU_nx376, 
         L1_3_L2_4_G3_MINI_ALU_nx396, L1_3_L2_4_G3_MINI_ALU_nx416, 
         L1_3_L2_4_G3_MINI_ALU_nx436, L1_3_L2_4_G3_MINI_ALU_nx454, 
         L1_3_L2_4_G3_MINI_ALU_nx456, L1_3_L2_4_G3_MINI_ALU_nx379, 
         L1_3_L2_4_G3_MINI_ALU_nx381, L1_3_L2_4_G3_MINI_ALU_nx383, 
         L1_3_L2_4_G3_MINI_ALU_nx387, L1_3_L2_4_G3_MINI_ALU_nx389, 
         L1_3_L2_4_G3_MINI_ALU_nx391, L1_3_L2_4_G3_MINI_ALU_nx395, 
         L1_3_L2_4_G3_MINI_ALU_nx399, L1_3_L2_4_G3_MINI_ALU_nx401, 
         L1_3_L2_4_G3_MINI_ALU_nx403, L1_3_L2_4_G3_MINI_ALU_nx405, 
         L1_3_L2_4_G3_MINI_ALU_nx409, L1_3_L2_4_G3_MINI_ALU_nx411, 
         L1_3_L2_4_G3_MINI_ALU_nx413, L1_3_L2_4_G3_MINI_ALU_nx415, 
         L1_3_L2_4_G3_MINI_ALU_nx419, L1_3_L2_4_G3_MINI_ALU_nx421, 
         L1_3_L2_4_G3_MINI_ALU_nx423, L1_3_L2_4_G3_MINI_ALU_nx425, 
         L1_3_L2_4_G3_MINI_ALU_nx429, L1_3_L2_4_G3_MINI_ALU_nx431, 
         L1_3_L2_4_G3_MINI_ALU_nx433, L1_3_L2_4_G3_MINI_ALU_nx435, 
         L1_3_L2_4_G3_MINI_ALU_nx439, L1_3_L2_4_G3_MINI_ALU_nx441, 
         L1_3_L2_4_G3_MINI_ALU_nx443, L1_3_L2_4_G3_MINI_ALU_nx445, 
         L1_3_L2_4_G3_MINI_ALU_nx449, L1_3_L2_4_G3_MINI_ALU_nx451, 
         L1_3_L2_4_G3_MINI_ALU_nx453, L1_3_L2_4_G3_MINI_ALU_nx455, 
         L1_3_L2_4_G3_MINI_ALU_nx461, L1_3_L2_4_G3_MINI_ALU_nx463, 
         L1_3_L2_4_G3_MINI_ALU_nx467, L1_3_L2_4_G3_MINI_ALU_nx469, 
         L1_3_L2_4_G3_MINI_ALU_nx471, L1_3_L2_4_G3_MINI_ALU_nx475, 
         L1_3_L2_4_G3_MINI_ALU_nx477, L1_3_L2_4_G3_MINI_ALU_nx479, 
         L1_3_L2_4_G3_MINI_ALU_nx483, L1_3_L2_4_G3_MINI_ALU_nx485, 
         L1_3_L2_4_G3_MINI_ALU_nx487, L1_3_L2_4_G3_MINI_ALU_nx491, 
         L1_3_L2_4_G3_MINI_ALU_nx493, L1_3_L2_4_G3_MINI_ALU_nx495, 
         L1_3_L2_4_G3_MINI_ALU_nx499, L1_3_L2_4_G3_MINI_ALU_nx501, 
         L1_3_L2_4_G3_MINI_ALU_nx503, L1_3_L2_4_G3_MINI_ALU_nx507, 
         L1_3_L2_4_G3_MINI_ALU_nx509, L1_3_L2_4_G3_MINI_ALU_nx511, 
         L1_3_L2_4_G3_MINI_ALU_nx515, L1_3_L2_4_G3_MINI_ALU_nx517, 
         L1_3_L2_4_G3_MINI_ALU_nx529, L1_3_L2_4_G3_MINI_ALU_nx531, 
         L1_3_L2_4_G3_MINI_ALU_nx534, L1_3_L2_4_G3_MINI_ALU_nx537, 
         L1_3_L2_4_G3_MINI_ALU_nx540, L1_3_L2_4_G3_MINI_ALU_nx544, 
         L1_3_L2_4_G3_MINI_ALU_nx547, L1_3_L2_4_G3_MINI_ALU_nx551, 
         L1_3_L2_4_G3_MINI_ALU_nx554, L1_3_L2_4_G3_MINI_ALU_nx558, 
         L1_3_L2_4_G3_MINI_ALU_nx561, L1_3_L2_4_G3_MINI_ALU_nx565, 
         L1_3_L2_4_G3_MINI_ALU_nx568, 
         L1_3_L2_4_G3_MINI_ALU_WindowCellShiftedLeft_16, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_16, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_15, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_14, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_13, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_12, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_11, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_10, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_16, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_15, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_14, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_13, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_12, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_11, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_10, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_9, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_8, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_7, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_6, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_5, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_4, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_3, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_2, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_1, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_0, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_16, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_15, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_14, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_13, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_12, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_11, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_10, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_9, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_8, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_7, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_6, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_5, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_4, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_3, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_2, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_1, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_0, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_16, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_15, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_14, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_13, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_12, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_11, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_10, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_9, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_8, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_7, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_6, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_5, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_4, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_3, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_2, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_1, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_0, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_nx4, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_nx8, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_nx12, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_nx16, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_nx20, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_nx24, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_nx80, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_nx328, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_nx384, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642, 
         L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644, 
         L1_4_L2_0_G3_MINI_ALU_AddPToBoothOperand, 
         L1_4_L2_0_G3_MINI_ALU_BoothOperand_16, 
         L1_4_L2_0_G3_MINI_ALU_BoothOperand_15, 
         L1_4_L2_0_G3_MINI_ALU_BoothOperand_14, 
         L1_4_L2_0_G3_MINI_ALU_BoothOperand_13, 
         L1_4_L2_0_G3_MINI_ALU_BoothOperand_12, 
         L1_4_L2_0_G3_MINI_ALU_BoothOperand_11, 
         L1_4_L2_0_G3_MINI_ALU_BoothOperand_10, 
         L1_4_L2_0_G3_MINI_ALU_BoothOperand_9, 
         L1_4_L2_0_G3_MINI_ALU_BoothOperand_8, 
         L1_4_L2_0_G3_MINI_ALU_BoothOperand_7, 
         L1_4_L2_0_G3_MINI_ALU_BoothOperand_6, 
         L1_4_L2_0_G3_MINI_ALU_BoothOperand_5, 
         L1_4_L2_0_G3_MINI_ALU_BoothOperand_4, 
         L1_4_L2_0_G3_MINI_ALU_BoothOperand_3, 
         L1_4_L2_0_G3_MINI_ALU_BoothOperand_2, 
         L1_4_L2_0_G3_MINI_ALU_BoothOperand_1, 
         L1_4_L2_0_G3_MINI_ALU_BoothOperand_0, 
         L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_16, 
         L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_15, 
         L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_14, 
         L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_13, 
         L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_12, 
         L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_11, 
         L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_10, 
         L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_9, 
         L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_8, 
         L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_7, 
         L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_6, 
         L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_5, 
         L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_4, 
         L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_3, 
         L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_2, 
         L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_1, 
         L1_4_L2_0_G3_MINI_ALU_BoothP_16, L1_4_L2_0_G3_MINI_ALU_BoothP_15, 
         L1_4_L2_0_G3_MINI_ALU_BoothP_14, L1_4_L2_0_G3_MINI_ALU_BoothP_13, 
         L1_4_L2_0_G3_MINI_ALU_BoothP_12, L1_4_L2_0_G3_MINI_ALU_BoothP_11, 
         L1_4_L2_0_G3_MINI_ALU_BoothP_10, L1_4_L2_0_G3_MINI_ALU_BoothP_9, 
         L1_4_L2_0_G3_MINI_ALU_BoothP_8, L1_4_L2_0_G3_MINI_ALU_BoothP_7, 
         L1_4_L2_0_G3_MINI_ALU_BoothP_6, L1_4_L2_0_G3_MINI_ALU_BoothP_5, 
         L1_4_L2_0_G3_MINI_ALU_BoothP_4, L1_4_L2_0_G3_MINI_ALU_BoothP_3, 
         L1_4_L2_0_G3_MINI_ALU_BoothP_2, L1_4_L2_0_G3_MINI_ALU_BoothP_1, 
         L1_4_L2_0_G3_MINI_ALU_BoothP_0, L1_4_L2_0_G3_MINI_ALU_nx0, 
         L1_4_L2_0_G3_MINI_ALU_nx6, L1_4_L2_0_G3_MINI_ALU_nx12, 
         L1_4_L2_0_G3_MINI_ALU_nx18, L1_4_L2_0_G3_MINI_ALU_nx24, 
         L1_4_L2_0_G3_MINI_ALU_nx30, L1_4_L2_0_G3_MINI_ALU_nx40, 
         L1_4_L2_0_G3_MINI_ALU_nx44, L1_4_L2_0_G3_MINI_ALU_nx48, 
         L1_4_L2_0_G3_MINI_ALU_nx52, L1_4_L2_0_G3_MINI_ALU_nx56, 
         L1_4_L2_0_G3_MINI_ALU_nx62, L1_4_L2_0_G3_MINI_ALU_nx154, 
         L1_4_L2_0_G3_MINI_ALU_nx316, L1_4_L2_0_G3_MINI_ALU_nx336, 
         L1_4_L2_0_G3_MINI_ALU_nx356, L1_4_L2_0_G3_MINI_ALU_nx376, 
         L1_4_L2_0_G3_MINI_ALU_nx396, L1_4_L2_0_G3_MINI_ALU_nx416, 
         L1_4_L2_0_G3_MINI_ALU_nx436, L1_4_L2_0_G3_MINI_ALU_nx454, 
         L1_4_L2_0_G3_MINI_ALU_nx456, L1_4_L2_0_G3_MINI_ALU_nx379, 
         L1_4_L2_0_G3_MINI_ALU_nx381, L1_4_L2_0_G3_MINI_ALU_nx383, 
         L1_4_L2_0_G3_MINI_ALU_nx387, L1_4_L2_0_G3_MINI_ALU_nx389, 
         L1_4_L2_0_G3_MINI_ALU_nx391, L1_4_L2_0_G3_MINI_ALU_nx395, 
         L1_4_L2_0_G3_MINI_ALU_nx399, L1_4_L2_0_G3_MINI_ALU_nx401, 
         L1_4_L2_0_G3_MINI_ALU_nx403, L1_4_L2_0_G3_MINI_ALU_nx405, 
         L1_4_L2_0_G3_MINI_ALU_nx409, L1_4_L2_0_G3_MINI_ALU_nx411, 
         L1_4_L2_0_G3_MINI_ALU_nx413, L1_4_L2_0_G3_MINI_ALU_nx415, 
         L1_4_L2_0_G3_MINI_ALU_nx419, L1_4_L2_0_G3_MINI_ALU_nx421, 
         L1_4_L2_0_G3_MINI_ALU_nx423, L1_4_L2_0_G3_MINI_ALU_nx425, 
         L1_4_L2_0_G3_MINI_ALU_nx429, L1_4_L2_0_G3_MINI_ALU_nx431, 
         L1_4_L2_0_G3_MINI_ALU_nx433, L1_4_L2_0_G3_MINI_ALU_nx435, 
         L1_4_L2_0_G3_MINI_ALU_nx439, L1_4_L2_0_G3_MINI_ALU_nx441, 
         L1_4_L2_0_G3_MINI_ALU_nx443, L1_4_L2_0_G3_MINI_ALU_nx445, 
         L1_4_L2_0_G3_MINI_ALU_nx449, L1_4_L2_0_G3_MINI_ALU_nx451, 
         L1_4_L2_0_G3_MINI_ALU_nx453, L1_4_L2_0_G3_MINI_ALU_nx455, 
         L1_4_L2_0_G3_MINI_ALU_nx461, L1_4_L2_0_G3_MINI_ALU_nx463, 
         L1_4_L2_0_G3_MINI_ALU_nx467, L1_4_L2_0_G3_MINI_ALU_nx469, 
         L1_4_L2_0_G3_MINI_ALU_nx471, L1_4_L2_0_G3_MINI_ALU_nx475, 
         L1_4_L2_0_G3_MINI_ALU_nx477, L1_4_L2_0_G3_MINI_ALU_nx479, 
         L1_4_L2_0_G3_MINI_ALU_nx483, L1_4_L2_0_G3_MINI_ALU_nx485, 
         L1_4_L2_0_G3_MINI_ALU_nx487, L1_4_L2_0_G3_MINI_ALU_nx491, 
         L1_4_L2_0_G3_MINI_ALU_nx493, L1_4_L2_0_G3_MINI_ALU_nx495, 
         L1_4_L2_0_G3_MINI_ALU_nx499, L1_4_L2_0_G3_MINI_ALU_nx501, 
         L1_4_L2_0_G3_MINI_ALU_nx503, L1_4_L2_0_G3_MINI_ALU_nx507, 
         L1_4_L2_0_G3_MINI_ALU_nx509, L1_4_L2_0_G3_MINI_ALU_nx511, 
         L1_4_L2_0_G3_MINI_ALU_nx515, L1_4_L2_0_G3_MINI_ALU_nx517, 
         L1_4_L2_0_G3_MINI_ALU_nx529, L1_4_L2_0_G3_MINI_ALU_nx531, 
         L1_4_L2_0_G3_MINI_ALU_nx534, L1_4_L2_0_G3_MINI_ALU_nx537, 
         L1_4_L2_0_G3_MINI_ALU_nx540, L1_4_L2_0_G3_MINI_ALU_nx544, 
         L1_4_L2_0_G3_MINI_ALU_nx547, L1_4_L2_0_G3_MINI_ALU_nx551, 
         L1_4_L2_0_G3_MINI_ALU_nx554, L1_4_L2_0_G3_MINI_ALU_nx558, 
         L1_4_L2_0_G3_MINI_ALU_nx561, L1_4_L2_0_G3_MINI_ALU_nx565, 
         L1_4_L2_0_G3_MINI_ALU_nx568, 
         L1_4_L2_0_G3_MINI_ALU_WindowCellShiftedLeft_16, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_16, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_15, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_14, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_13, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_12, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_11, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_10, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_16, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_15, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_14, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_13, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_12, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_11, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_10, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_9, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_8, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_7, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_6, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_5, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_4, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_3, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_2, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_1, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_0, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_16, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_15, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_14, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_13, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_12, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_11, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_10, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_9, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_8, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_7, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_6, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_5, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_4, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_3, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_2, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_1, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_0, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_16, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_15, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_14, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_13, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_12, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_11, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_10, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_9, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_8, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_7, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_6, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_5, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_4, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_3, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_2, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_1, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_0, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_nx4, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_nx8, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_nx12, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_nx16, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_nx20, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_nx24, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_nx80, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_nx328, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_nx384, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642, 
         L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644, 
         L1_4_L2_1_G3_MINI_ALU_AddPToBoothOperand, 
         L1_4_L2_1_G3_MINI_ALU_BoothOperand_16, 
         L1_4_L2_1_G3_MINI_ALU_BoothOperand_15, 
         L1_4_L2_1_G3_MINI_ALU_BoothOperand_14, 
         L1_4_L2_1_G3_MINI_ALU_BoothOperand_13, 
         L1_4_L2_1_G3_MINI_ALU_BoothOperand_12, 
         L1_4_L2_1_G3_MINI_ALU_BoothOperand_11, 
         L1_4_L2_1_G3_MINI_ALU_BoothOperand_10, 
         L1_4_L2_1_G3_MINI_ALU_BoothOperand_9, 
         L1_4_L2_1_G3_MINI_ALU_BoothOperand_8, 
         L1_4_L2_1_G3_MINI_ALU_BoothOperand_7, 
         L1_4_L2_1_G3_MINI_ALU_BoothOperand_6, 
         L1_4_L2_1_G3_MINI_ALU_BoothOperand_5, 
         L1_4_L2_1_G3_MINI_ALU_BoothOperand_4, 
         L1_4_L2_1_G3_MINI_ALU_BoothOperand_3, 
         L1_4_L2_1_G3_MINI_ALU_BoothOperand_2, 
         L1_4_L2_1_G3_MINI_ALU_BoothOperand_1, 
         L1_4_L2_1_G3_MINI_ALU_BoothOperand_0, 
         L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_16, 
         L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_15, 
         L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_14, 
         L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_13, 
         L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_12, 
         L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_11, 
         L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_10, 
         L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_9, 
         L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_8, 
         L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_7, 
         L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_6, 
         L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_5, 
         L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_4, 
         L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_3, 
         L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_2, 
         L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_1, 
         L1_4_L2_1_G3_MINI_ALU_BoothP_16, L1_4_L2_1_G3_MINI_ALU_BoothP_15, 
         L1_4_L2_1_G3_MINI_ALU_BoothP_14, L1_4_L2_1_G3_MINI_ALU_BoothP_13, 
         L1_4_L2_1_G3_MINI_ALU_BoothP_12, L1_4_L2_1_G3_MINI_ALU_BoothP_11, 
         L1_4_L2_1_G3_MINI_ALU_BoothP_10, L1_4_L2_1_G3_MINI_ALU_BoothP_9, 
         L1_4_L2_1_G3_MINI_ALU_BoothP_8, L1_4_L2_1_G3_MINI_ALU_BoothP_7, 
         L1_4_L2_1_G3_MINI_ALU_BoothP_6, L1_4_L2_1_G3_MINI_ALU_BoothP_5, 
         L1_4_L2_1_G3_MINI_ALU_BoothP_4, L1_4_L2_1_G3_MINI_ALU_BoothP_3, 
         L1_4_L2_1_G3_MINI_ALU_BoothP_2, L1_4_L2_1_G3_MINI_ALU_BoothP_1, 
         L1_4_L2_1_G3_MINI_ALU_BoothP_0, L1_4_L2_1_G3_MINI_ALU_nx0, 
         L1_4_L2_1_G3_MINI_ALU_nx6, L1_4_L2_1_G3_MINI_ALU_nx12, 
         L1_4_L2_1_G3_MINI_ALU_nx18, L1_4_L2_1_G3_MINI_ALU_nx24, 
         L1_4_L2_1_G3_MINI_ALU_nx30, L1_4_L2_1_G3_MINI_ALU_nx40, 
         L1_4_L2_1_G3_MINI_ALU_nx44, L1_4_L2_1_G3_MINI_ALU_nx48, 
         L1_4_L2_1_G3_MINI_ALU_nx52, L1_4_L2_1_G3_MINI_ALU_nx56, 
         L1_4_L2_1_G3_MINI_ALU_nx62, L1_4_L2_1_G3_MINI_ALU_nx154, 
         L1_4_L2_1_G3_MINI_ALU_nx316, L1_4_L2_1_G3_MINI_ALU_nx336, 
         L1_4_L2_1_G3_MINI_ALU_nx356, L1_4_L2_1_G3_MINI_ALU_nx376, 
         L1_4_L2_1_G3_MINI_ALU_nx396, L1_4_L2_1_G3_MINI_ALU_nx416, 
         L1_4_L2_1_G3_MINI_ALU_nx436, L1_4_L2_1_G3_MINI_ALU_nx454, 
         L1_4_L2_1_G3_MINI_ALU_nx456, L1_4_L2_1_G3_MINI_ALU_nx379, 
         L1_4_L2_1_G3_MINI_ALU_nx381, L1_4_L2_1_G3_MINI_ALU_nx383, 
         L1_4_L2_1_G3_MINI_ALU_nx387, L1_4_L2_1_G3_MINI_ALU_nx389, 
         L1_4_L2_1_G3_MINI_ALU_nx391, L1_4_L2_1_G3_MINI_ALU_nx395, 
         L1_4_L2_1_G3_MINI_ALU_nx399, L1_4_L2_1_G3_MINI_ALU_nx401, 
         L1_4_L2_1_G3_MINI_ALU_nx403, L1_4_L2_1_G3_MINI_ALU_nx405, 
         L1_4_L2_1_G3_MINI_ALU_nx409, L1_4_L2_1_G3_MINI_ALU_nx411, 
         L1_4_L2_1_G3_MINI_ALU_nx413, L1_4_L2_1_G3_MINI_ALU_nx415, 
         L1_4_L2_1_G3_MINI_ALU_nx419, L1_4_L2_1_G3_MINI_ALU_nx421, 
         L1_4_L2_1_G3_MINI_ALU_nx423, L1_4_L2_1_G3_MINI_ALU_nx425, 
         L1_4_L2_1_G3_MINI_ALU_nx429, L1_4_L2_1_G3_MINI_ALU_nx431, 
         L1_4_L2_1_G3_MINI_ALU_nx433, L1_4_L2_1_G3_MINI_ALU_nx435, 
         L1_4_L2_1_G3_MINI_ALU_nx439, L1_4_L2_1_G3_MINI_ALU_nx441, 
         L1_4_L2_1_G3_MINI_ALU_nx443, L1_4_L2_1_G3_MINI_ALU_nx445, 
         L1_4_L2_1_G3_MINI_ALU_nx449, L1_4_L2_1_G3_MINI_ALU_nx451, 
         L1_4_L2_1_G3_MINI_ALU_nx453, L1_4_L2_1_G3_MINI_ALU_nx455, 
         L1_4_L2_1_G3_MINI_ALU_nx461, L1_4_L2_1_G3_MINI_ALU_nx463, 
         L1_4_L2_1_G3_MINI_ALU_nx467, L1_4_L2_1_G3_MINI_ALU_nx469, 
         L1_4_L2_1_G3_MINI_ALU_nx471, L1_4_L2_1_G3_MINI_ALU_nx475, 
         L1_4_L2_1_G3_MINI_ALU_nx477, L1_4_L2_1_G3_MINI_ALU_nx479, 
         L1_4_L2_1_G3_MINI_ALU_nx483, L1_4_L2_1_G3_MINI_ALU_nx485, 
         L1_4_L2_1_G3_MINI_ALU_nx487, L1_4_L2_1_G3_MINI_ALU_nx491, 
         L1_4_L2_1_G3_MINI_ALU_nx493, L1_4_L2_1_G3_MINI_ALU_nx495, 
         L1_4_L2_1_G3_MINI_ALU_nx499, L1_4_L2_1_G3_MINI_ALU_nx501, 
         L1_4_L2_1_G3_MINI_ALU_nx503, L1_4_L2_1_G3_MINI_ALU_nx507, 
         L1_4_L2_1_G3_MINI_ALU_nx509, L1_4_L2_1_G3_MINI_ALU_nx511, 
         L1_4_L2_1_G3_MINI_ALU_nx515, L1_4_L2_1_G3_MINI_ALU_nx517, 
         L1_4_L2_1_G3_MINI_ALU_nx529, L1_4_L2_1_G3_MINI_ALU_nx531, 
         L1_4_L2_1_G3_MINI_ALU_nx534, L1_4_L2_1_G3_MINI_ALU_nx537, 
         L1_4_L2_1_G3_MINI_ALU_nx540, L1_4_L2_1_G3_MINI_ALU_nx544, 
         L1_4_L2_1_G3_MINI_ALU_nx547, L1_4_L2_1_G3_MINI_ALU_nx551, 
         L1_4_L2_1_G3_MINI_ALU_nx554, L1_4_L2_1_G3_MINI_ALU_nx558, 
         L1_4_L2_1_G3_MINI_ALU_nx561, L1_4_L2_1_G3_MINI_ALU_nx565, 
         L1_4_L2_1_G3_MINI_ALU_nx568, 
         L1_4_L2_1_G3_MINI_ALU_WindowCellShiftedLeft_16, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_16, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_15, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_14, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_13, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_12, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_11, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_10, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_16, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_15, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_14, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_13, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_12, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_11, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_10, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_9, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_8, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_7, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_6, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_5, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_4, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_3, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_2, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_1, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_0, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_16, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_15, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_14, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_13, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_12, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_11, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_10, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_9, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_8, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_7, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_6, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_5, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_4, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_3, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_2, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_1, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_0, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_16, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_15, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_14, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_13, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_12, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_11, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_10, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_9, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_8, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_7, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_6, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_5, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_4, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_3, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_2, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_1, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_0, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_nx4, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_nx8, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_nx12, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_nx16, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_nx20, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_nx24, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_nx80, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_nx328, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_nx384, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642, 
         L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644, 
         L1_4_L2_2_G4_MINI_ALU_AddPToBoothOperand, 
         L1_4_L2_2_G4_MINI_ALU_BoothOperand_16, 
         L1_4_L2_2_G4_MINI_ALU_BoothOperand_15, 
         L1_4_L2_2_G4_MINI_ALU_BoothOperand_14, 
         L1_4_L2_2_G4_MINI_ALU_BoothOperand_13, 
         L1_4_L2_2_G4_MINI_ALU_BoothOperand_12, 
         L1_4_L2_2_G4_MINI_ALU_BoothOperand_11, 
         L1_4_L2_2_G4_MINI_ALU_BoothOperand_10, 
         L1_4_L2_2_G4_MINI_ALU_BoothOperand_9, 
         L1_4_L2_2_G4_MINI_ALU_BoothOperand_8, 
         L1_4_L2_2_G4_MINI_ALU_BoothOperand_7, 
         L1_4_L2_2_G4_MINI_ALU_BoothOperand_6, 
         L1_4_L2_2_G4_MINI_ALU_BoothOperand_5, 
         L1_4_L2_2_G4_MINI_ALU_BoothOperand_4, 
         L1_4_L2_2_G4_MINI_ALU_BoothOperand_3, 
         L1_4_L2_2_G4_MINI_ALU_BoothOperand_2, 
         L1_4_L2_2_G4_MINI_ALU_BoothOperand_1, 
         L1_4_L2_2_G4_MINI_ALU_BoothOperand_0, 
         L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_16, 
         L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_15, 
         L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_14, 
         L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_13, 
         L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_12, 
         L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_11, 
         L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_10, 
         L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_9, 
         L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_8, 
         L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_7, 
         L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_6, 
         L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_5, 
         L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_4, 
         L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_3, 
         L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_2, 
         L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_1, 
         L1_4_L2_2_G4_MINI_ALU_BoothP_16, L1_4_L2_2_G4_MINI_ALU_BoothP_15, 
         L1_4_L2_2_G4_MINI_ALU_BoothP_14, L1_4_L2_2_G4_MINI_ALU_BoothP_13, 
         L1_4_L2_2_G4_MINI_ALU_BoothP_12, L1_4_L2_2_G4_MINI_ALU_BoothP_11, 
         L1_4_L2_2_G4_MINI_ALU_BoothP_10, L1_4_L2_2_G4_MINI_ALU_BoothP_9, 
         L1_4_L2_2_G4_MINI_ALU_BoothP_8, L1_4_L2_2_G4_MINI_ALU_BoothP_7, 
         L1_4_L2_2_G4_MINI_ALU_BoothP_6, L1_4_L2_2_G4_MINI_ALU_BoothP_5, 
         L1_4_L2_2_G4_MINI_ALU_BoothP_4, L1_4_L2_2_G4_MINI_ALU_BoothP_3, 
         L1_4_L2_2_G4_MINI_ALU_BoothP_2, L1_4_L2_2_G4_MINI_ALU_BoothP_1, 
         L1_4_L2_2_G4_MINI_ALU_BoothP_0, L1_4_L2_2_G4_MINI_ALU_nx0, 
         L1_4_L2_2_G4_MINI_ALU_nx6, L1_4_L2_2_G4_MINI_ALU_nx12, 
         L1_4_L2_2_G4_MINI_ALU_nx18, L1_4_L2_2_G4_MINI_ALU_nx24, 
         L1_4_L2_2_G4_MINI_ALU_nx30, L1_4_L2_2_G4_MINI_ALU_nx40, 
         L1_4_L2_2_G4_MINI_ALU_nx44, L1_4_L2_2_G4_MINI_ALU_nx48, 
         L1_4_L2_2_G4_MINI_ALU_nx52, L1_4_L2_2_G4_MINI_ALU_nx56, 
         L1_4_L2_2_G4_MINI_ALU_nx62, L1_4_L2_2_G4_MINI_ALU_nx154, 
         L1_4_L2_2_G4_MINI_ALU_nx316, L1_4_L2_2_G4_MINI_ALU_nx336, 
         L1_4_L2_2_G4_MINI_ALU_nx356, L1_4_L2_2_G4_MINI_ALU_nx376, 
         L1_4_L2_2_G4_MINI_ALU_nx396, L1_4_L2_2_G4_MINI_ALU_nx416, 
         L1_4_L2_2_G4_MINI_ALU_nx436, L1_4_L2_2_G4_MINI_ALU_nx454, 
         L1_4_L2_2_G4_MINI_ALU_nx456, L1_4_L2_2_G4_MINI_ALU_nx379, 
         L1_4_L2_2_G4_MINI_ALU_nx381, L1_4_L2_2_G4_MINI_ALU_nx383, 
         L1_4_L2_2_G4_MINI_ALU_nx387, L1_4_L2_2_G4_MINI_ALU_nx389, 
         L1_4_L2_2_G4_MINI_ALU_nx391, L1_4_L2_2_G4_MINI_ALU_nx395, 
         L1_4_L2_2_G4_MINI_ALU_nx399, L1_4_L2_2_G4_MINI_ALU_nx401, 
         L1_4_L2_2_G4_MINI_ALU_nx403, L1_4_L2_2_G4_MINI_ALU_nx405, 
         L1_4_L2_2_G4_MINI_ALU_nx409, L1_4_L2_2_G4_MINI_ALU_nx411, 
         L1_4_L2_2_G4_MINI_ALU_nx413, L1_4_L2_2_G4_MINI_ALU_nx415, 
         L1_4_L2_2_G4_MINI_ALU_nx419, L1_4_L2_2_G4_MINI_ALU_nx421, 
         L1_4_L2_2_G4_MINI_ALU_nx423, L1_4_L2_2_G4_MINI_ALU_nx425, 
         L1_4_L2_2_G4_MINI_ALU_nx429, L1_4_L2_2_G4_MINI_ALU_nx431, 
         L1_4_L2_2_G4_MINI_ALU_nx433, L1_4_L2_2_G4_MINI_ALU_nx435, 
         L1_4_L2_2_G4_MINI_ALU_nx439, L1_4_L2_2_G4_MINI_ALU_nx441, 
         L1_4_L2_2_G4_MINI_ALU_nx443, L1_4_L2_2_G4_MINI_ALU_nx445, 
         L1_4_L2_2_G4_MINI_ALU_nx449, L1_4_L2_2_G4_MINI_ALU_nx451, 
         L1_4_L2_2_G4_MINI_ALU_nx453, L1_4_L2_2_G4_MINI_ALU_nx455, 
         L1_4_L2_2_G4_MINI_ALU_nx461, L1_4_L2_2_G4_MINI_ALU_nx463, 
         L1_4_L2_2_G4_MINI_ALU_nx467, L1_4_L2_2_G4_MINI_ALU_nx469, 
         L1_4_L2_2_G4_MINI_ALU_nx471, L1_4_L2_2_G4_MINI_ALU_nx475, 
         L1_4_L2_2_G4_MINI_ALU_nx477, L1_4_L2_2_G4_MINI_ALU_nx479, 
         L1_4_L2_2_G4_MINI_ALU_nx483, L1_4_L2_2_G4_MINI_ALU_nx485, 
         L1_4_L2_2_G4_MINI_ALU_nx487, L1_4_L2_2_G4_MINI_ALU_nx491, 
         L1_4_L2_2_G4_MINI_ALU_nx493, L1_4_L2_2_G4_MINI_ALU_nx495, 
         L1_4_L2_2_G4_MINI_ALU_nx499, L1_4_L2_2_G4_MINI_ALU_nx501, 
         L1_4_L2_2_G4_MINI_ALU_nx503, L1_4_L2_2_G4_MINI_ALU_nx507, 
         L1_4_L2_2_G4_MINI_ALU_nx509, L1_4_L2_2_G4_MINI_ALU_nx511, 
         L1_4_L2_2_G4_MINI_ALU_nx515, L1_4_L2_2_G4_MINI_ALU_nx517, 
         L1_4_L2_2_G4_MINI_ALU_nx529, L1_4_L2_2_G4_MINI_ALU_nx531, 
         L1_4_L2_2_G4_MINI_ALU_nx534, L1_4_L2_2_G4_MINI_ALU_nx537, 
         L1_4_L2_2_G4_MINI_ALU_nx540, L1_4_L2_2_G4_MINI_ALU_nx544, 
         L1_4_L2_2_G4_MINI_ALU_nx547, L1_4_L2_2_G4_MINI_ALU_nx551, 
         L1_4_L2_2_G4_MINI_ALU_nx554, L1_4_L2_2_G4_MINI_ALU_nx558, 
         L1_4_L2_2_G4_MINI_ALU_nx561, L1_4_L2_2_G4_MINI_ALU_nx565, 
         L1_4_L2_2_G4_MINI_ALU_nx568, 
         L1_4_L2_2_G4_MINI_ALU_WindowCellShiftedLeft_16, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDin_16, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDin_15, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDin_14, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDin_13, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDin_12, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDin_11, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDin_10, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_16, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_15, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_14, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_13, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_12, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_11, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_10, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_9, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_8, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_7, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_6, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_5, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_4, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_3, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_2, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_1, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_0, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_16, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_15, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_14, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_13, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_12, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_11, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_10, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_9, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_8, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_7, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_6, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_5, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_4, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_3, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_2, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_1, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_0, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_16, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_15, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_14, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_13, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_12, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_11, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_10, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_9, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_8, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_7, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_6, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_5, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_4, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_3, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_2, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_1, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_0, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_nx4, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_nx8, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_nx12, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_nx16, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_nx20, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_nx24, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_nx80, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_nx328, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_nx384, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642, 
         L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644, 
         L1_4_L2_3_G5_MINI_ALU_AddPToBoothOperand, 
         L1_4_L2_3_G5_MINI_ALU_BoothOperand_16, 
         L1_4_L2_3_G5_MINI_ALU_BoothOperand_15, 
         L1_4_L2_3_G5_MINI_ALU_BoothOperand_14, 
         L1_4_L2_3_G5_MINI_ALU_BoothOperand_13, 
         L1_4_L2_3_G5_MINI_ALU_BoothOperand_12, 
         L1_4_L2_3_G5_MINI_ALU_BoothOperand_11, 
         L1_4_L2_3_G5_MINI_ALU_BoothOperand_10, 
         L1_4_L2_3_G5_MINI_ALU_BoothOperand_9, 
         L1_4_L2_3_G5_MINI_ALU_BoothOperand_8, 
         L1_4_L2_3_G5_MINI_ALU_BoothOperand_7, 
         L1_4_L2_3_G5_MINI_ALU_BoothOperand_6, 
         L1_4_L2_3_G5_MINI_ALU_BoothOperand_5, 
         L1_4_L2_3_G5_MINI_ALU_BoothOperand_4, 
         L1_4_L2_3_G5_MINI_ALU_BoothOperand_3, 
         L1_4_L2_3_G5_MINI_ALU_BoothOperand_2, 
         L1_4_L2_3_G5_MINI_ALU_BoothOperand_1, 
         L1_4_L2_3_G5_MINI_ALU_BoothOperand_0, 
         L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_16, 
         L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_15, 
         L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_14, 
         L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_13, 
         L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_12, 
         L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_11, 
         L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_10, 
         L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_9, 
         L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_8, 
         L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_7, 
         L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_6, 
         L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_5, 
         L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_4, 
         L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_3, 
         L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_2, 
         L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_1, 
         L1_4_L2_3_G5_MINI_ALU_BoothP_16, L1_4_L2_3_G5_MINI_ALU_BoothP_15, 
         L1_4_L2_3_G5_MINI_ALU_BoothP_14, L1_4_L2_3_G5_MINI_ALU_BoothP_13, 
         L1_4_L2_3_G5_MINI_ALU_BoothP_12, L1_4_L2_3_G5_MINI_ALU_BoothP_11, 
         L1_4_L2_3_G5_MINI_ALU_BoothP_10, L1_4_L2_3_G5_MINI_ALU_BoothP_9, 
         L1_4_L2_3_G5_MINI_ALU_BoothP_8, L1_4_L2_3_G5_MINI_ALU_BoothP_7, 
         L1_4_L2_3_G5_MINI_ALU_BoothP_6, L1_4_L2_3_G5_MINI_ALU_BoothP_5, 
         L1_4_L2_3_G5_MINI_ALU_BoothP_4, L1_4_L2_3_G5_MINI_ALU_BoothP_3, 
         L1_4_L2_3_G5_MINI_ALU_BoothP_2, L1_4_L2_3_G5_MINI_ALU_BoothP_1, 
         L1_4_L2_3_G5_MINI_ALU_BoothP_0, L1_4_L2_3_G5_MINI_ALU_nx0, 
         L1_4_L2_3_G5_MINI_ALU_nx6, L1_4_L2_3_G5_MINI_ALU_nx12, 
         L1_4_L2_3_G5_MINI_ALU_nx18, L1_4_L2_3_G5_MINI_ALU_nx24, 
         L1_4_L2_3_G5_MINI_ALU_nx30, L1_4_L2_3_G5_MINI_ALU_nx40, 
         L1_4_L2_3_G5_MINI_ALU_nx44, L1_4_L2_3_G5_MINI_ALU_nx48, 
         L1_4_L2_3_G5_MINI_ALU_nx52, L1_4_L2_3_G5_MINI_ALU_nx56, 
         L1_4_L2_3_G5_MINI_ALU_nx62, L1_4_L2_3_G5_MINI_ALU_nx154, 
         L1_4_L2_3_G5_MINI_ALU_nx316, L1_4_L2_3_G5_MINI_ALU_nx336, 
         L1_4_L2_3_G5_MINI_ALU_nx356, L1_4_L2_3_G5_MINI_ALU_nx376, 
         L1_4_L2_3_G5_MINI_ALU_nx396, L1_4_L2_3_G5_MINI_ALU_nx416, 
         L1_4_L2_3_G5_MINI_ALU_nx436, L1_4_L2_3_G5_MINI_ALU_nx454, 
         L1_4_L2_3_G5_MINI_ALU_nx456, L1_4_L2_3_G5_MINI_ALU_nx379, 
         L1_4_L2_3_G5_MINI_ALU_nx381, L1_4_L2_3_G5_MINI_ALU_nx383, 
         L1_4_L2_3_G5_MINI_ALU_nx387, L1_4_L2_3_G5_MINI_ALU_nx389, 
         L1_4_L2_3_G5_MINI_ALU_nx391, L1_4_L2_3_G5_MINI_ALU_nx395, 
         L1_4_L2_3_G5_MINI_ALU_nx399, L1_4_L2_3_G5_MINI_ALU_nx401, 
         L1_4_L2_3_G5_MINI_ALU_nx403, L1_4_L2_3_G5_MINI_ALU_nx405, 
         L1_4_L2_3_G5_MINI_ALU_nx409, L1_4_L2_3_G5_MINI_ALU_nx411, 
         L1_4_L2_3_G5_MINI_ALU_nx413, L1_4_L2_3_G5_MINI_ALU_nx415, 
         L1_4_L2_3_G5_MINI_ALU_nx419, L1_4_L2_3_G5_MINI_ALU_nx421, 
         L1_4_L2_3_G5_MINI_ALU_nx423, L1_4_L2_3_G5_MINI_ALU_nx425, 
         L1_4_L2_3_G5_MINI_ALU_nx429, L1_4_L2_3_G5_MINI_ALU_nx431, 
         L1_4_L2_3_G5_MINI_ALU_nx433, L1_4_L2_3_G5_MINI_ALU_nx435, 
         L1_4_L2_3_G5_MINI_ALU_nx439, L1_4_L2_3_G5_MINI_ALU_nx441, 
         L1_4_L2_3_G5_MINI_ALU_nx443, L1_4_L2_3_G5_MINI_ALU_nx445, 
         L1_4_L2_3_G5_MINI_ALU_nx449, L1_4_L2_3_G5_MINI_ALU_nx451, 
         L1_4_L2_3_G5_MINI_ALU_nx453, L1_4_L2_3_G5_MINI_ALU_nx455, 
         L1_4_L2_3_G5_MINI_ALU_nx461, L1_4_L2_3_G5_MINI_ALU_nx463, 
         L1_4_L2_3_G5_MINI_ALU_nx467, L1_4_L2_3_G5_MINI_ALU_nx469, 
         L1_4_L2_3_G5_MINI_ALU_nx471, L1_4_L2_3_G5_MINI_ALU_nx475, 
         L1_4_L2_3_G5_MINI_ALU_nx477, L1_4_L2_3_G5_MINI_ALU_nx479, 
         L1_4_L2_3_G5_MINI_ALU_nx483, L1_4_L2_3_G5_MINI_ALU_nx485, 
         L1_4_L2_3_G5_MINI_ALU_nx487, L1_4_L2_3_G5_MINI_ALU_nx491, 
         L1_4_L2_3_G5_MINI_ALU_nx493, L1_4_L2_3_G5_MINI_ALU_nx495, 
         L1_4_L2_3_G5_MINI_ALU_nx499, L1_4_L2_3_G5_MINI_ALU_nx501, 
         L1_4_L2_3_G5_MINI_ALU_nx503, L1_4_L2_3_G5_MINI_ALU_nx507, 
         L1_4_L2_3_G5_MINI_ALU_nx509, L1_4_L2_3_G5_MINI_ALU_nx511, 
         L1_4_L2_3_G5_MINI_ALU_nx515, L1_4_L2_3_G5_MINI_ALU_nx517, 
         L1_4_L2_3_G5_MINI_ALU_nx529, L1_4_L2_3_G5_MINI_ALU_nx531, 
         L1_4_L2_3_G5_MINI_ALU_nx534, L1_4_L2_3_G5_MINI_ALU_nx537, 
         L1_4_L2_3_G5_MINI_ALU_nx540, L1_4_L2_3_G5_MINI_ALU_nx544, 
         L1_4_L2_3_G5_MINI_ALU_nx547, L1_4_L2_3_G5_MINI_ALU_nx551, 
         L1_4_L2_3_G5_MINI_ALU_nx554, L1_4_L2_3_G5_MINI_ALU_nx558, 
         L1_4_L2_3_G5_MINI_ALU_nx561, L1_4_L2_3_G5_MINI_ALU_nx565, 
         L1_4_L2_3_G5_MINI_ALU_nx568, 
         L1_4_L2_3_G5_MINI_ALU_WindowCellShiftedLeft_16, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_16, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_15, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_14, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_13, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_12, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_11, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_10, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_16, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_15, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_14, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_13, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_12, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_11, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_10, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_9, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_8, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_7, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_6, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_5, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_4, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_3, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_2, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_1, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_0, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_16, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_15, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_14, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_13, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_12, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_11, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_10, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_9, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_8, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_7, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_6, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_5, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_4, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_3, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_2, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_1, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_0, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_16, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_15, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_14, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_13, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_12, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_11, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_10, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_9, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_8, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_7, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_6, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_5, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_4, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_3, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_2, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_1, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_0, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_nx4, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_nx8, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_nx12, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_nx16, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_nx20, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_nx24, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_nx80, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_nx328, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_nx384, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642, 
         L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644, 
         L1_4_L2_4_G5_MINI_ALU_AddPToBoothOperand, 
         L1_4_L2_4_G5_MINI_ALU_BoothOperand_16, 
         L1_4_L2_4_G5_MINI_ALU_BoothOperand_15, 
         L1_4_L2_4_G5_MINI_ALU_BoothOperand_14, 
         L1_4_L2_4_G5_MINI_ALU_BoothOperand_13, 
         L1_4_L2_4_G5_MINI_ALU_BoothOperand_12, 
         L1_4_L2_4_G5_MINI_ALU_BoothOperand_11, 
         L1_4_L2_4_G5_MINI_ALU_BoothOperand_10, 
         L1_4_L2_4_G5_MINI_ALU_BoothOperand_9, 
         L1_4_L2_4_G5_MINI_ALU_BoothOperand_8, 
         L1_4_L2_4_G5_MINI_ALU_BoothOperand_7, 
         L1_4_L2_4_G5_MINI_ALU_BoothOperand_6, 
         L1_4_L2_4_G5_MINI_ALU_BoothOperand_5, 
         L1_4_L2_4_G5_MINI_ALU_BoothOperand_4, 
         L1_4_L2_4_G5_MINI_ALU_BoothOperand_3, 
         L1_4_L2_4_G5_MINI_ALU_BoothOperand_2, 
         L1_4_L2_4_G5_MINI_ALU_BoothOperand_1, 
         L1_4_L2_4_G5_MINI_ALU_BoothOperand_0, 
         L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_16, 
         L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_15, 
         L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_14, 
         L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_13, 
         L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_12, 
         L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_11, 
         L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_10, 
         L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_9, 
         L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_8, 
         L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_7, 
         L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_6, 
         L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_5, 
         L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_4, 
         L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_3, 
         L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_2, 
         L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_1, 
         L1_4_L2_4_G5_MINI_ALU_BoothP_16, L1_4_L2_4_G5_MINI_ALU_BoothP_15, 
         L1_4_L2_4_G5_MINI_ALU_BoothP_14, L1_4_L2_4_G5_MINI_ALU_BoothP_13, 
         L1_4_L2_4_G5_MINI_ALU_BoothP_12, L1_4_L2_4_G5_MINI_ALU_BoothP_11, 
         L1_4_L2_4_G5_MINI_ALU_BoothP_10, L1_4_L2_4_G5_MINI_ALU_BoothP_9, 
         L1_4_L2_4_G5_MINI_ALU_BoothP_8, L1_4_L2_4_G5_MINI_ALU_BoothP_7, 
         L1_4_L2_4_G5_MINI_ALU_BoothP_6, L1_4_L2_4_G5_MINI_ALU_BoothP_5, 
         L1_4_L2_4_G5_MINI_ALU_BoothP_4, L1_4_L2_4_G5_MINI_ALU_BoothP_3, 
         L1_4_L2_4_G5_MINI_ALU_BoothP_2, L1_4_L2_4_G5_MINI_ALU_BoothP_1, 
         L1_4_L2_4_G5_MINI_ALU_BoothP_0, L1_4_L2_4_G5_MINI_ALU_nx0, 
         L1_4_L2_4_G5_MINI_ALU_nx6, L1_4_L2_4_G5_MINI_ALU_nx12, 
         L1_4_L2_4_G5_MINI_ALU_nx18, L1_4_L2_4_G5_MINI_ALU_nx24, 
         L1_4_L2_4_G5_MINI_ALU_nx30, L1_4_L2_4_G5_MINI_ALU_nx40, 
         L1_4_L2_4_G5_MINI_ALU_nx44, L1_4_L2_4_G5_MINI_ALU_nx48, 
         L1_4_L2_4_G5_MINI_ALU_nx52, L1_4_L2_4_G5_MINI_ALU_nx56, 
         L1_4_L2_4_G5_MINI_ALU_nx62, L1_4_L2_4_G5_MINI_ALU_nx154, 
         L1_4_L2_4_G5_MINI_ALU_nx316, L1_4_L2_4_G5_MINI_ALU_nx336, 
         L1_4_L2_4_G5_MINI_ALU_nx356, L1_4_L2_4_G5_MINI_ALU_nx376, 
         L1_4_L2_4_G5_MINI_ALU_nx396, L1_4_L2_4_G5_MINI_ALU_nx416, 
         L1_4_L2_4_G5_MINI_ALU_nx436, L1_4_L2_4_G5_MINI_ALU_nx454, 
         L1_4_L2_4_G5_MINI_ALU_nx456, L1_4_L2_4_G5_MINI_ALU_nx379, 
         L1_4_L2_4_G5_MINI_ALU_nx381, L1_4_L2_4_G5_MINI_ALU_nx383, 
         L1_4_L2_4_G5_MINI_ALU_nx387, L1_4_L2_4_G5_MINI_ALU_nx389, 
         L1_4_L2_4_G5_MINI_ALU_nx391, L1_4_L2_4_G5_MINI_ALU_nx395, 
         L1_4_L2_4_G5_MINI_ALU_nx399, L1_4_L2_4_G5_MINI_ALU_nx401, 
         L1_4_L2_4_G5_MINI_ALU_nx403, L1_4_L2_4_G5_MINI_ALU_nx405, 
         L1_4_L2_4_G5_MINI_ALU_nx409, L1_4_L2_4_G5_MINI_ALU_nx411, 
         L1_4_L2_4_G5_MINI_ALU_nx413, L1_4_L2_4_G5_MINI_ALU_nx415, 
         L1_4_L2_4_G5_MINI_ALU_nx419, L1_4_L2_4_G5_MINI_ALU_nx421, 
         L1_4_L2_4_G5_MINI_ALU_nx423, L1_4_L2_4_G5_MINI_ALU_nx425, 
         L1_4_L2_4_G5_MINI_ALU_nx429, L1_4_L2_4_G5_MINI_ALU_nx431, 
         L1_4_L2_4_G5_MINI_ALU_nx433, L1_4_L2_4_G5_MINI_ALU_nx435, 
         L1_4_L2_4_G5_MINI_ALU_nx439, L1_4_L2_4_G5_MINI_ALU_nx441, 
         L1_4_L2_4_G5_MINI_ALU_nx443, L1_4_L2_4_G5_MINI_ALU_nx445, 
         L1_4_L2_4_G5_MINI_ALU_nx449, L1_4_L2_4_G5_MINI_ALU_nx451, 
         L1_4_L2_4_G5_MINI_ALU_nx453, L1_4_L2_4_G5_MINI_ALU_nx455, 
         L1_4_L2_4_G5_MINI_ALU_nx461, L1_4_L2_4_G5_MINI_ALU_nx463, 
         L1_4_L2_4_G5_MINI_ALU_nx467, L1_4_L2_4_G5_MINI_ALU_nx469, 
         L1_4_L2_4_G5_MINI_ALU_nx471, L1_4_L2_4_G5_MINI_ALU_nx475, 
         L1_4_L2_4_G5_MINI_ALU_nx477, L1_4_L2_4_G5_MINI_ALU_nx479, 
         L1_4_L2_4_G5_MINI_ALU_nx483, L1_4_L2_4_G5_MINI_ALU_nx485, 
         L1_4_L2_4_G5_MINI_ALU_nx487, L1_4_L2_4_G5_MINI_ALU_nx491, 
         L1_4_L2_4_G5_MINI_ALU_nx493, L1_4_L2_4_G5_MINI_ALU_nx495, 
         L1_4_L2_4_G5_MINI_ALU_nx499, L1_4_L2_4_G5_MINI_ALU_nx501, 
         L1_4_L2_4_G5_MINI_ALU_nx503, L1_4_L2_4_G5_MINI_ALU_nx507, 
         L1_4_L2_4_G5_MINI_ALU_nx509, L1_4_L2_4_G5_MINI_ALU_nx511, 
         L1_4_L2_4_G5_MINI_ALU_nx515, L1_4_L2_4_G5_MINI_ALU_nx517, 
         L1_4_L2_4_G5_MINI_ALU_nx529, L1_4_L2_4_G5_MINI_ALU_nx531, 
         L1_4_L2_4_G5_MINI_ALU_nx534, L1_4_L2_4_G5_MINI_ALU_nx537, 
         L1_4_L2_4_G5_MINI_ALU_nx540, L1_4_L2_4_G5_MINI_ALU_nx544, 
         L1_4_L2_4_G5_MINI_ALU_nx547, L1_4_L2_4_G5_MINI_ALU_nx551, 
         L1_4_L2_4_G5_MINI_ALU_nx554, L1_4_L2_4_G5_MINI_ALU_nx558, 
         L1_4_L2_4_G5_MINI_ALU_nx561, L1_4_L2_4_G5_MINI_ALU_nx565, 
         L1_4_L2_4_G5_MINI_ALU_nx568, 
         L1_4_L2_4_G5_MINI_ALU_WindowCellShiftedLeft_16, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_16, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_15, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_14, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_13, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_12, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_11, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_10, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_16, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_15, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_14, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_13, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_12, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_11, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_10, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_9, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_8, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_7, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_6, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_5, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_4, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_3, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_2, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_1, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_0, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_16, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_15, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_14, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_13, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_12, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_11, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_10, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_9, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_8, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_7, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_6, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_5, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_4, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_3, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_2, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_1, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_0, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_16, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_15, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_14, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_13, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_12, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_11, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_10, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_9, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_8, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_7, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_6, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_5, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_4, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_3, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_2, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_1, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_0, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_nx4, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_nx8, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_nx12, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_nx16, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_nx20, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_nx24, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_nx80, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_nx328, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_nx384, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642, 
         L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644, nx1336, nx1338, 
         nx1340, nx1342, nx1344, nx1346, nx1348, nx1350, nx1352, nx1354, nx1356, 
         nx1358, nx1360, nx1362, nx1364, nx1366, nx1368, nx1370, nx1372, nx1374, 
         nx1376, nx1378, nx1380, nx1382, nx1384, nx1386, nx1388, nx1390, nx1392, 
         nx1394, nx1396, nx1398, nx1400, nx1402, nx1404, nx1406, nx1408, nx1410, 
         nx1412, nx1414, nx1416, nx1418, nx1420, nx1422, nx1424, nx1426, nx1428, 
         nx1430, nx1432, nx1434, nx1436, nx1438, nx1440, nx1442, nx1444, nx1446, 
         nx1448, nx1450, nx1452, nx1454, nx1456, nx1458, nx1460, nx1462, nx1464, 
         nx1466, nx1468, nx1470, nx1472, nx1474, nx1476, nx1478, nx1480, nx1482, 
         nx1484, nx1486, nx1488, nx1490, nx1492, nx1494, nx1496, nx1498, nx1500, 
         nx1502, nx1504, nx1506, nx1508, nx1510, nx1512, nx1514, nx1516, nx1520, 
         nx1522, nx1524, nx1526, nx1528, nx1530, nx1532, nx1534, nx1536, nx1538, 
         nx1540, nx1542, nx1544, nx1546, nx1548, nx1550, nx1552, nx1554, nx1556, 
         nx1558, nx1560, nx1562, nx1564, nx1566, nx1568, nx1570, nx1572, nx1574, 
         nx1576, nx1578, nx1580, nx1582, nx1584, nx1586, nx1588, nx1590, nx1592, 
         nx1594, nx1596, nx1598, nx1600, nx1602, nx1604, nx1606, nx1608, nx1610, 
         nx1612, nx1614, nx1616, nx1618, nx1620, nx1622, nx1624, nx1626, nx1628, 
         nx1630, nx1632, nx1634, nx1636, nx1638, nx1640, nx1642, nx1644, nx1646, 
         nx1648, nx1650, nx1652, nx1654, nx1656, nx1658, nx1660, nx1662, nx1664, 
         nx1666, nx1668, nx1670, nx1672, nx1674, nx1676, nx1678, nx1680, nx1682, 
         nx1684, nx1686, nx1688, nx1690, nx1692, nx1694, nx1696, nx1698, nx1700, 
         nx1702, nx1704, nx1706, nx1708, nx1710, nx1712, nx1714, nx1716, nx1718, 
         nx1720, nx1722, nx1724, nx1726, nx1728, nx1730, nx1732, nx1734, nx1736, 
         nx1738, nx1740, nx1742, nx1744, nx1746, nx1748, nx1750, nx1752, nx1754, 
         nx1756, nx1758, nx1760, nx1762, nx1764, nx1768, nx1770, nx1772, nx1774, 
         nx1776, nx1778, nx1780, nx1782, nx1784, nx1786, nx1788, nx1790, nx1792, 
         nx1794, nx1796, nx1798, nx1800, nx1802, nx1804, nx1806, nx1808, nx1810, 
         nx1812, nx1814, nx1816, nx1818, nx1820, nx1822, nx1824, nx1826, nx1828, 
         nx1830, nx1832, nx1834, nx1836, nx1838, nx1840, nx1842, nx1844, nx1846, 
         nx1848, nx1850, nx1852, nx1854, nx1856, nx1858, nx1860, nx1862, nx1864, 
         nx1866, nx1868, nx1870, nx1872, nx1874, nx1876, nx1878, nx1880, nx1882, 
         nx1884, nx1886, nx1888, nx1890, nx1892, nx1894, nx1896, nx1898, nx1900, 
         nx1902, nx1904, nx1906, nx1908, nx1910, nx1912, nx1914, nx1916, nx1918, 
         nx1920, nx1922, nx1924, nx1926, nx1928, nx1930, nx1932, nx1934, nx1936, 
         nx1938, nx1940, nx1942, nx1944, nx1946, nx1948, nx1950, nx1952, nx1954, 
         nx1956, nx1958, nx1960, nx1962, nx1964, nx1966, nx1968, nx1970, nx1972, 
         nx1974, nx1976, nx1978, nx1980, nx1982, nx1984, nx1986, nx1988, nx1990, 
         nx1992, nx1994, nx1996, nx1998, nx2000, nx2002, nx2004, nx2006, nx2008, 
         nx2010, nx2012, nx2016, nx2018, nx2020, nx2022, nx2024, nx2026, nx2028, 
         nx2030, nx2032, nx2034, nx2036, nx2038, nx2040, nx2042, nx2044, nx2046, 
         nx2048, nx2050, nx2052, nx2054, nx2056, nx2058, nx2060, nx2062, nx2064, 
         nx2066, nx2068, nx2070, nx2072, nx2074, nx2076, nx2078, nx2080, nx2082, 
         nx2084, nx2086, nx2088, nx2090, nx2092, nx2094, nx2096, nx2098, nx2100, 
         nx2102, nx2104, nx2106, nx2108, nx2110, nx2112, nx2114, nx2116, nx2118, 
         nx2120, nx2122, nx2124, nx2126, nx2128, nx2130, nx2132, nx2134, nx2136, 
         nx2138, nx2140, nx2142, nx2144, nx2146, nx2148, nx2150, nx2152, nx2154, 
         nx2156, nx2158, nx2160, nx2162, nx2164, nx2166, nx2168, nx2170, nx2172, 
         nx2174, nx2176, nx2178, nx2180, nx2182, nx2184, nx2186, nx2188, nx2190, 
         nx2192, nx2194, nx2196, nx2198, nx2200, nx2202, nx2204, nx2206, nx2208, 
         nx2210, nx2212, nx2214, nx2216, nx2218, nx2220, nx2222, nx2224, nx2226, 
         nx2228, nx2230, nx2232, nx2234, nx2236, nx2238, nx2240, nx2242, nx2244, 
         nx2246, nx2248, nx2250, nx2252, nx2254, nx2256, nx2258, nx2260, nx2264, 
         nx2266, nx2268, nx2270, nx2272, nx2274, nx2276, nx2278, nx2280, nx2282, 
         nx2284, nx2286, nx2288, nx2290, nx2292, nx2294, nx2296, nx2298, nx2300, 
         nx2302, nx2304, nx2306, nx2308, nx2310, nx2312, nx2314, nx2316, nx2318, 
         nx2320, nx2322, nx2324, nx2326, nx2328, nx2330, nx2332, nx2334, nx2336, 
         nx2338, nx2340, nx2342, nx2344, nx2346, nx2348, nx2350, nx2352, nx2354, 
         nx2356, nx2358, nx2360, nx2362, nx2364, nx2366, nx2368, nx2370, nx2372, 
         nx2374, nx2376, nx2378, nx2380, nx2382, nx2384, nx2386, nx2388, nx2390, 
         nx2392, nx2394, nx2396, nx2398, nx2400, nx2402, nx2404, nx2406, nx2408, 
         nx2410, nx2412, nx2414, nx2416, nx2418, nx2420, nx2422, nx2424, nx2426, 
         nx2428, nx2430, nx2432, nx2434, nx2436, nx2438, nx2440, nx2442, nx2444, 
         nx2446, nx2448, nx2450, nx2452, nx2454, nx2456, nx2458, nx2460, nx2462, 
         nx2464, nx2466, nx2468, nx2470, nx2472, nx2474, nx2476, nx2478, nx2480, 
         nx2482, nx2484, nx2486, nx2488, nx2490, nx2492, nx2494, nx2496, nx2498, 
         nx2500, nx2502, nx2504, nx2506, nx2508, nx2512, nx2514, nx2516, nx2518, 
         nx2520, nx2522, nx2524, nx2526, nx2528, nx2530, nx2532, nx2534, nx2536, 
         nx2538, nx2540, nx2542, nx2544, nx2546, nx2548, nx2550, nx2552, nx2554, 
         nx2556, nx2558, nx2560, nx2562, nx2564, nx2566, nx2568, nx2570, nx2572, 
         nx2574, nx2576, nx2578, nx2580, nx2582, nx2584, nx2586, nx2588, nx2590, 
         nx2592, nx2594, nx2596, nx2598, nx2600, nx2602, nx2604, nx2606, nx2608, 
         nx2610, nx2612, nx2614, nx2616, nx2618, nx2620, nx2622, nx2624, nx2626, 
         nx2628, nx2630, nx2632, nx2634, nx2636, nx2638, nx2640, nx2642, nx2644, 
         nx2646, nx2648, nx2650, nx2652, nx2654, nx2656, nx2658, nx2660, nx2662, 
         nx2664, nx2666, nx2668, nx2670, nx2672, nx2674, nx2676, nx2678, nx2680, 
         nx2682, nx2684, nx2686, nx2688, nx2690, nx2692, nx2694, nx2696, nx2698, 
         nx2700, nx2702, nx2704, nx2706, nx2708, nx2710, nx2712, nx2714, nx2716, 
         nx2718, nx2720, nx2722, nx2724, nx2726, nx2728, nx2730, nx2732, nx2734, 
         nx2736, nx2738, nx2740, nx2742, nx2744, nx2746, nx2748, nx2750, nx2752, 
         nx2754, nx2756, nx2760, nx2762, nx2764, nx2766, nx2768, nx2770, nx2772, 
         nx2774, nx2776, nx2778, nx2780, nx2782, nx2784, nx2786, nx2788, nx2790, 
         nx2792, nx2794, nx2796, nx2798, nx2800, nx2802, nx2804, nx2806, nx2808, 
         nx2810, nx2812, nx2814, nx2816, nx2818, nx2820, nx2822, nx2824, nx2826, 
         nx2828, nx2830, nx2832, nx2834, nx2836, nx2838, nx2840, nx2842, nx2844, 
         nx2846, nx2848, nx2850, nx2852, nx2854, nx2856, nx2858, nx2860, nx2862, 
         nx2864, nx2866, nx2868, nx2870, nx2872, nx2874, nx2876, nx2878, nx2880, 
         nx2882, nx2884, nx2886, nx2888, nx2890, nx2892, nx2894, nx2896, nx2898, 
         nx2900, nx2902, nx2904, nx2906, nx2908, nx2910, nx2912, nx2914, nx2916, 
         nx2918, nx2920, nx2922, nx2924, nx2926, nx2928, nx2930, nx2932, nx2934, 
         nx2936, nx2938, nx2940, nx2942, nx2944, nx2946, nx2948, nx2950, nx2952, 
         nx2954, nx2956, nx2958, nx2960, nx2962, nx2964, nx2966, nx2968, nx2970, 
         nx2972, nx2974, nx2976, nx2978, nx2980, nx2982, nx2984, nx2986, nx2988, 
         nx2990, nx2992, nx2994, nx2996, nx2998, nx3000, nx3002, nx3004, nx3008, 
         nx3010, nx3012, nx3014, nx3016, nx3018, nx3020, nx3022, nx3024, nx3026, 
         nx3028, nx3030, nx3032, nx3034, nx3036, nx3038, nx3040, nx3042, nx3044, 
         nx3046, nx3048, nx3050, nx3052, nx3054, nx3056, nx3058, nx3060, nx3062, 
         nx3064, nx3066, nx3068, nx3070, nx3072, nx3074, nx3076, nx3078, nx3080, 
         nx3082, nx3084, nx3086, nx3088, nx3090, nx3092, nx3094, nx3096, nx3098, 
         nx3100, nx3102, nx3104, nx3106, nx3108, nx3110, nx3112, nx3114, nx3116, 
         nx3118, nx3120, nx3122, nx3124, nx3126, nx3128, nx3130, nx3132, nx3134, 
         nx3136, nx3138, nx3140, nx3142, nx3144, nx3146, nx3148, nx3150, nx3152, 
         nx3154, nx3156, nx3158, nx3160, nx3162, nx3164, nx3166, nx3168, nx3170, 
         nx3172, nx3174, nx3176, nx3178, nx3180, nx3182, nx3184, nx3186, nx3188, 
         nx3190, nx3192, nx3194, nx3196, nx3198, nx3200, nx3202, nx3204, nx3206, 
         nx3208, nx3210, nx3212, nx3214, nx3216, nx3218, nx3220, nx3222, nx3224, 
         nx3226, nx3228, nx3230, nx3232, nx3234, nx3236, nx3238, nx3240, nx3242, 
         nx3244, nx3246, nx3248, nx3250, nx3252, nx3256, nx3258, nx3260, nx3262, 
         nx3264, nx3266, nx3268, nx3270, nx3272, nx3274, nx3276, nx3278, nx3280, 
         nx3282, nx3284, nx3286, nx3288, nx3290, nx3292, nx3294, nx3296, nx3298, 
         nx3300, nx3302, nx3304, nx3306, nx3308, nx3310, nx3312, nx3314, nx3316, 
         nx3318, nx3320, nx3322, nx3324, nx3326, nx3328, nx3330, nx3332, nx3334, 
         nx3336, nx3338, nx3340, nx3342, nx3344, nx3346, nx3348, nx3350, nx3352, 
         nx3354, nx3356, nx3358, nx3360, nx3362, nx3364, nx3366, nx3368, nx3370, 
         nx3372, nx3374, nx3376, nx3378, nx3380, nx3382, nx3384, nx3386, nx3388, 
         nx3390, nx3392, nx3394, nx3396, nx3398, nx3400, nx3402, nx3404, nx3406, 
         nx3408, nx3410, nx3412, nx3414, nx3416, nx3418, nx3420, nx3422, nx3424, 
         nx3426, nx3428, nx3430, nx3432, nx3434, nx3436, nx3438, nx3440, nx3442, 
         nx3444, nx3446, nx3448, nx3450, nx3452, nx3454, nx3456, nx3458, nx3460, 
         nx3462, nx3464, nx3466, nx3468, nx3470, nx3472, nx3474, nx3476, nx3478, 
         nx3480, nx3482, nx3484, nx3486, nx3488, nx3490, nx3492, nx3494, nx3496, 
         nx3498, nx3500, nx3504, nx3506, nx3508, nx3510, nx3512, nx3514, nx3516, 
         nx3518, nx3520, nx3522, nx3524, nx3526, nx3528, nx3530, nx3532, nx3534, 
         nx3536, nx3538, nx3540, nx3542, nx3544, nx3546, nx3548, nx3550, nx3552, 
         nx3554, nx3556, nx3558, nx3560, nx3562, nx3564, nx3566, nx3568, nx3570, 
         nx3572, nx3574, nx3576, nx3578, nx3580, nx3582, nx3584, nx3586, nx3588, 
         nx3590, nx3592, nx3594, nx3596, nx3598, nx3600, nx3602, nx3604, nx3606, 
         nx3608, nx3610, nx3612, nx3614, nx3616, nx3618, nx3620, nx3622, nx3624, 
         nx3626, nx3628, nx3630, nx3632, nx3634, nx3636, nx3638, nx3640, nx3642, 
         nx3644, nx3646, nx3648, nx3650, nx3652, nx3654, nx3656, nx3658, nx3660, 
         nx3662, nx3664, nx3666, nx3668, nx3670, nx3672, nx3674, nx3676, nx3678, 
         nx3680, nx3682, nx3684, nx3686, nx3688, nx3690, nx3692, nx3694, nx3696, 
         nx3698, nx3700, nx3702, nx3704, nx3706, nx3708, nx3710, nx3712, nx3714, 
         nx3716, nx3718, nx3720, nx3722, nx3724, nx3726, nx3728, nx3730, nx3732, 
         nx3734, nx3736, nx3738, nx3740, nx3742, nx3744, nx3746, nx3748, nx3752, 
         nx3754, nx3756, nx3758, nx3760, nx3762, nx3764, nx3766, nx3768, nx3770, 
         nx3772, nx3774, nx3776, nx3778, nx3780, nx3782, nx3784, nx3786, nx3788, 
         nx3790, nx3792, nx3794, nx3796, nx3798, nx3800, nx3802, nx3804, nx3806, 
         nx3808, nx3810, nx3812, nx3814, nx3816, nx3818, nx3820, nx3822, nx3824, 
         nx3826, nx3828, nx3830, nx3832, nx3834, nx3836, nx3838, nx3840, nx3842, 
         nx3844, nx3846, nx3848, nx3850, nx3852, nx3854, nx3856, nx3858, nx3860, 
         nx3862, nx3864, nx3866, nx3868, nx3870, nx3872, nx3874, nx3876, nx3878, 
         nx3880, nx3882, nx3884, nx3886, nx3888, nx3890, nx3892, nx3894, nx3896, 
         nx3898, nx3900, nx3902, nx3904, nx3906, nx3908, nx3910, nx3912, nx3914, 
         nx3916, nx3918, nx3920, nx3922, nx3924, nx3926, nx3928, nx3930, nx3932, 
         nx3934, nx3936, nx3938, nx3940, nx3942, nx3944, nx3946, nx3948, nx3950, 
         nx3952, nx3954, nx3956, nx3958, nx3960, nx3962, nx3964, nx3966, nx3968, 
         nx3970, nx3972, nx3974, nx3976, nx3978, nx3980, nx3982, nx3984, nx3986, 
         nx3988, nx3990, nx3992, nx3994, nx3996, nx4000, nx4002, nx4004, nx4006, 
         nx4008, nx4010, nx4012, nx4014, nx4016, nx4018, nx4020, nx4022, nx4024, 
         nx4026, nx4028, nx4030, nx4032, nx4034, nx4036, nx4038, nx4040, nx4042, 
         nx4044, nx4046, nx4048, nx4050, nx4052, nx4054, nx4056, nx4058, nx4060, 
         nx4062, nx4064, nx4066, nx4068, nx4070, nx4072, nx4074, nx4076, nx4078, 
         nx4080, nx4082, nx4084, nx4086, nx4088, nx4090, nx4092, nx4094, nx4096, 
         nx4098, nx4100, nx4102, nx4104, nx4106, nx4108, nx4110, nx4112, nx4114, 
         nx4116, nx4118, nx4120, nx4122, nx4124, nx4126, nx4128, nx4130, nx4132, 
         nx4134, nx4136, nx4138, nx4140, nx4142, nx4144, nx4146, nx4148, nx4150, 
         nx4152, nx4154, nx4156, nx4158, nx4160, nx4162, nx4164, nx4166, nx4168, 
         nx4170, nx4172, nx4174, nx4176, nx4178, nx4180, nx4182, nx4184, nx4186, 
         nx4188, nx4190, nx4192, nx4194, nx4196, nx4198, nx4200, nx4202, nx4204, 
         nx4206, nx4208, nx4210, nx4212, nx4214, nx4216, nx4218, nx4220, nx4222, 
         nx4224, nx4226, nx4228, nx4230, nx4232, nx4234, nx4236, nx4238, nx4240, 
         nx4242, nx4244, nx4248, nx4250, nx4252, nx4254, nx4256, nx4258, nx4260, 
         nx4262, nx4264, nx4266, nx4268, nx4270, nx4272, nx4274, nx4276, nx4278, 
         nx4280, nx4282, nx4284, nx4286, nx4288, nx4290, nx4292, nx4294, nx4296, 
         nx4298, nx4300, nx4302, nx4304, nx4306, nx4308, nx4310, nx4312, nx4314, 
         nx4316, nx4318, nx4320, nx4322, nx4324, nx4326, nx4328, nx4330, nx4332, 
         nx4334, nx4336, nx4338, nx4340, nx4342, nx4344, nx4346, nx4348, nx4350, 
         nx4352, nx4354, nx4356, nx4358, nx4360, nx4362, nx4364, nx4366, nx4368, 
         nx4370, nx4372, nx4374, nx4376, nx4378, nx4380, nx4382, nx4384, nx4386, 
         nx4388, nx4390, nx4392, nx4394, nx4396, nx4398, nx4400, nx4402, nx4404, 
         nx4406, nx4408, nx4410, nx4412, nx4414, nx4416, nx4418, nx4420, nx4422, 
         nx4424, nx4426, nx4428, nx4430, nx4432, nx4434, nx4436, nx4438, nx4440, 
         nx4442, nx4444, nx4446, nx4448, nx4450, nx4452, nx4454, nx4456, nx4458, 
         nx4460, nx4462, nx4464, nx4466, nx4468, nx4470, nx4472, nx4474, nx4476, 
         nx4478, nx4480, nx4482, nx4484, nx4486, nx4488, nx4490, nx4492, nx4496, 
         nx4498, nx4500, nx4502, nx4504, nx4506, nx4508, nx4510, nx4512, nx4514, 
         nx4516, nx4518, nx4520, nx4522, nx4524, nx4526, nx4528, nx4530, nx4532, 
         nx4534, nx4536, nx4538, nx4540, nx4542, nx4544, nx4546, nx4548, nx4550, 
         nx4552, nx4554, nx4556, nx4558, nx4560, nx4562, nx4564, nx4566, nx4568, 
         nx4570, nx4572, nx4574, nx4576, nx4578, nx4580, nx4582, nx4584, nx4586, 
         nx4588, nx4590, nx4592, nx4594, nx4596, nx4598, nx4600, nx4602, nx4604, 
         nx4606, nx4608, nx4610, nx4612, nx4614, nx4616, nx4618, nx4620, nx4622, 
         nx4624, nx4626, nx4628, nx4630, nx4632, nx4634, nx4636, nx4638, nx4640, 
         nx4642, nx4644, nx4646, nx4648, nx4650, nx4652, nx4654, nx4656, nx4658, 
         nx4660, nx4662, nx4664, nx4666, nx4668, nx4670, nx4672, nx4674, nx4676, 
         nx4678, nx4680, nx4682, nx4684, nx4686, nx4688, nx4690, nx4692, nx4694, 
         nx4696, nx4698, nx4700, nx4702, nx4704, nx4706, nx4708, nx4710, nx4712, 
         nx4714, nx4716, nx4718, nx4720, nx4722, nx4724, nx4726, nx4728, nx4730, 
         nx4732, nx4734, nx4736, nx4738, nx4740, nx4744, nx4746, nx4748, nx4750, 
         nx4752, nx4754, nx4756, nx4758, nx4760, nx4762, nx4764, nx4766, nx4768, 
         nx4770, nx4772, nx4774, nx4776, nx4778, nx4780, nx4782, nx4784, nx4786, 
         nx4788, nx4790, nx4792, nx4794, nx4796, nx4798, nx4800, nx4802, nx4804, 
         nx4806, nx4808, nx4810, nx4812, nx4814, nx4816, nx4818, nx4820, nx4822, 
         nx4824, nx4826, nx4828, nx4830, nx4832, nx4834, nx4836, nx4838, nx4840, 
         nx4842, nx4844, nx4846, nx4848, nx4850, nx4852, nx4854, nx4856, nx4858, 
         nx4860, nx4862, nx4864, nx4866, nx4868, nx4870, nx4872, nx4874, nx4876, 
         nx4878, nx4880, nx4882, nx4884, nx4886, nx4888, nx4890, nx4892, nx4894, 
         nx4896, nx4898, nx4900, nx4902, nx4904, nx4906, nx4908, nx4910, nx4912, 
         nx4914, nx4916, nx4918, nx4920, nx4922, nx4924, nx4926, nx4928, nx4930, 
         nx4932, nx4934, nx4936, nx4938, nx4940, nx4942, nx4944, nx4946, nx4948, 
         nx4950, nx4952, nx4954, nx4956, nx4958, nx4960, nx4962, nx4964, nx4966, 
         nx4968, nx4970, nx4972, nx4974, nx4976, nx4978, nx4980, nx4982, nx4984, 
         nx4986, nx4988, nx4992, nx4994, nx4996, nx4998, nx5000, nx5002, nx5004, 
         nx5006, nx5008, nx5010, nx5012, nx5014, nx5016, nx5018, nx5020, nx5022, 
         nx5024, nx5026, nx5028, nx5030, nx5032, nx5034, nx5036, nx5038, nx5040, 
         nx5042, nx5044, nx5046, nx5048, nx5050, nx5052, nx5054, nx5056, nx5058, 
         nx5060, nx5062, nx5064, nx5066, nx5068, nx5070, nx5072, nx5074, nx5076, 
         nx5078, nx5080, nx5082, nx5084, nx5086, nx5088, nx5090, nx5092, nx5094, 
         nx5096, nx5098, nx5100, nx5102, nx5104, nx5106, nx5108, nx5110, nx5112, 
         nx5114, nx5116, nx5118, nx5120, nx5122, nx5124, nx5126, nx5128, nx5130, 
         nx5132, nx5134, nx5136, nx5138, nx5140, nx5142, nx5144, nx5146, nx5148, 
         nx5150, nx5152, nx5154, nx5156, nx5158, nx5160, nx5162, nx5164, nx5166, 
         nx5168, nx5170, nx5172, nx5174, nx5176, nx5178, nx5180, nx5182, nx5184, 
         nx5186, nx5188, nx5190, nx5192, nx5194, nx5196, nx5198, nx5200, nx5202, 
         nx5204, nx5206, nx5208, nx5210, nx5212, nx5214, nx5216, nx5218, nx5220, 
         nx5222, nx5224, nx5226, nx5228, nx5230, nx5232, nx5234, nx5236, nx5240, 
         nx5242, nx5244, nx5246, nx5248, nx5250, nx5252, nx5254, nx5256, nx5258, 
         nx5260, nx5262, nx5264, nx5266, nx5268, nx5270, nx5272, nx5274, nx5276, 
         nx5278, nx5280, nx5282, nx5284, nx5286, nx5288, nx5290, nx5292, nx5294, 
         nx5296, nx5298, nx5300, nx5302, nx5304, nx5306, nx5308, nx5310, nx5312, 
         nx5314, nx5316, nx5318, nx5320, nx5322, nx5324, nx5326, nx5328, nx5330, 
         nx5332, nx5334, nx5336, nx5338, nx5340, nx5342, nx5344, nx5346, nx5348, 
         nx5350, nx5352, nx5354, nx5356, nx5358, nx5360, nx5362, nx5364, nx5366, 
         nx5368, nx5370, nx5372, nx5374, nx5376, nx5378, nx5380, nx5382, nx5384, 
         nx5386, nx5388, nx5390, nx5392, nx5394, nx5396, nx5398, nx5400, nx5402, 
         nx5404, nx5406, nx5408, nx5410, nx5412, nx5414, nx5416, nx5418, nx5420, 
         nx5422, nx5424, nx5426, nx5428, nx5430, nx5432, nx5434, nx5436, nx5438, 
         nx5440, nx5442, nx5444, nx5446, nx5448, nx5450, nx5452, nx5454, nx5456, 
         nx5458, nx5460, nx5462, nx5464, nx5466, nx5468, nx5470, nx5472, nx5474, 
         nx5476, nx5478, nx5480, nx5482, nx5484, nx5488, nx5490, nx5492, nx5494, 
         nx5496, nx5498, nx5500, nx5502, nx5504, nx5506, nx5508, nx5510, nx5512, 
         nx5514, nx5516, nx5518, nx5520, nx5522, nx5524, nx5526, nx5528, nx5530, 
         nx5532, nx5534, nx5536, nx5538, nx5540, nx5542, nx5544, nx5546, nx5548, 
         nx5550, nx5552, nx5554, nx5556, nx5558, nx5560, nx5562, nx5564, nx5566, 
         nx5568, nx5570, nx5572, nx5574, nx5576, nx5578, nx5580, nx5582, nx5584, 
         nx5586, nx5588, nx5590, nx5592, nx5594, nx5596, nx5598, nx5600, nx5602, 
         nx5604, nx5606, nx5608, nx5610, nx5612, nx5614, nx5616, nx5618, nx5620, 
         nx5622, nx5624, nx5626, nx5628, nx5630, nx5632, nx5634, nx5636, nx5638, 
         nx5640, nx5642, nx5644, nx5646, nx5648, nx5650, nx5652, nx5654, nx5656, 
         nx5658, nx5660, nx5662, nx5664, nx5666, nx5668, nx5670, nx5672, nx5674, 
         nx5676, nx5678, nx5680, nx5682, nx5684, nx5686, nx5688, nx5690, nx5692, 
         nx5694, nx5696, nx5698, nx5700, nx5702, nx5704, nx5706, nx5708, nx5710, 
         nx5712, nx5714, nx5716, nx5718, nx5720, nx5722, nx5724, nx5726, nx5728, 
         nx5730, nx5732, nx5736, nx5738, nx5740, nx5742, nx5744, nx5746, nx5748, 
         nx5750, nx5752, nx5754, nx5756, nx5758, nx5760, nx5762, nx5764, nx5766, 
         nx5768, nx5770, nx5772, nx5774, nx5776, nx5778, nx5780, nx5782, nx5784, 
         nx5786, nx5788, nx5790, nx5792, nx5794, nx5796, nx5798, nx5800, nx5802, 
         nx5804, nx5806, nx5808, nx5810, nx5812, nx5814, nx5816, nx5818, nx5820, 
         nx5822, nx5824, nx5826, nx5828, nx5830, nx5832, nx5834, nx5836, nx5838, 
         nx5840, nx5842, nx5844, nx5846, nx5848, nx5850, nx5852, nx5854, nx5856, 
         nx5858, nx5860, nx5862, nx5864, nx5866, nx5868, nx5870, nx5872, nx5874, 
         nx5876, nx5878, nx5880, nx5882, nx5884, nx5886, nx5888, nx5890, nx5892, 
         nx5894, nx5896, nx5898, nx5900, nx5902, nx5904, nx5906, nx5908, nx5910, 
         nx5912, nx5914, nx5916, nx5918, nx5920, nx5922, nx5924, nx5926, nx5928, 
         nx5930, nx5932, nx5934, nx5936, nx5938, nx5940, nx5942, nx5944, nx5946, 
         nx5948, nx5950, nx5952, nx5954, nx5956, nx5958, nx5960, nx5962, nx5964, 
         nx5966, nx5968, nx5970, nx5972, nx5974, nx5976, nx5978, nx5980, nx5984, 
         nx5986, nx5988, nx5990, nx5992, nx5994, nx5996, nx5998, nx6000, nx6002, 
         nx6004, nx6006, nx6008, nx6010, nx6012, nx6014, nx6016, nx6018, nx6020, 
         nx6022, nx6024, nx6026, nx6028, nx6030, nx6032, nx6034, nx6036, nx6038, 
         nx6040, nx6042, nx6044, nx6046, nx6048, nx6050, nx6052, nx6054, nx6056, 
         nx6058, nx6060, nx6062, nx6064, nx6066, nx6068, nx6070, nx6072, nx6074, 
         nx6076, nx6078, nx6080, nx6082, nx6084, nx6086, nx6088, nx6090, nx6092, 
         nx6094, nx6096, nx6098, nx6100, nx6102, nx6104, nx6106, nx6108, nx6110, 
         nx6112, nx6114, nx6116, nx6118, nx6120, nx6122, nx6124, nx6126, nx6128, 
         nx6130, nx6132, nx6134, nx6136, nx6138, nx6140, nx6142, nx6144, nx6146, 
         nx6148, nx6150, nx6152, nx6154, nx6156, nx6158, nx6160, nx6162, nx6164, 
         nx6166, nx6168, nx6170, nx6172, nx6174, nx6176, nx6178, nx6180, nx6182, 
         nx6184, nx6186, nx6188, nx6190, nx6192, nx6194, nx6196, nx6198, nx6200, 
         nx6202, nx6204, nx6206, nx6208, nx6210, nx6212, nx6214, nx6216, nx6218, 
         nx6220, nx6222, nx6224, nx6226, nx6228, nx6232, nx6234, nx6236, nx6238, 
         nx6240, nx6242, nx6244, nx6246, nx6248, nx6250, nx6252, nx6254, nx6256, 
         nx6258, nx6260, nx6262, nx6264, nx6266, nx6268, nx6270, nx6272, nx6274, 
         nx6276, nx6278, nx6280, nx6282, nx6284, nx6286, nx6288, nx6290, nx6292, 
         nx6294, nx6296, nx6298, nx6300, nx6302, nx6304, nx6306, nx6308, nx6310, 
         nx6312, nx6314, nx6316, nx6318, nx6320, nx6322, nx6324, nx6326, nx6328, 
         nx6330, nx6332, nx6334, nx6336, nx6338, nx6340, nx6342, nx6344, nx6346, 
         nx6348, nx6350, nx6352, nx6354, nx6356, nx6358, nx6360, nx6362, nx6364, 
         nx6366, nx6368, nx6370, nx6372, nx6374, nx6376, nx6378, nx6380, nx6382, 
         nx6384, nx6386, nx6388, nx6390, nx6392, nx6394, nx6396, nx6398, nx6400, 
         nx6402, nx6404, nx6406, nx6408, nx6410, nx6412, nx6414, nx6416, nx6418, 
         nx6420, nx6422, nx6424, nx6426, nx6428, nx6430, nx6432, nx6434, nx6436, 
         nx6438, nx6440, nx6442, nx6444, nx6446, nx6448, nx6450, nx6452, nx6454, 
         nx6456, nx6458, nx6460, nx6462, nx6464, nx6466, nx6468, nx6470, nx6472, 
         nx6474, nx6476, nx6480, nx6482, nx6484, nx6486, nx6488, nx6490, nx6492, 
         nx6494, nx6496, nx6498, nx6500, nx6502, nx6504, nx6506, nx6508, nx6510, 
         nx6512, nx6514, nx6516, nx6518, nx6520, nx6522, nx6524, nx6526, nx6528, 
         nx6530, nx6532, nx6534, nx6536, nx6538, nx6540, nx6542, nx6544, nx6546, 
         nx6548, nx6550, nx6552, nx6554, nx6556, nx6558, nx6560, nx6562, nx6564, 
         nx6566, nx6568, nx6570, nx6572, nx6574, nx6576, nx6578, nx6580, nx6582, 
         nx6584, nx6586, nx6588, nx6590, nx6592, nx6594, nx6596, nx6598, nx6600, 
         nx6602, nx6604, nx6606, nx6608, nx6610, nx6612, nx6614, nx6616, nx6618, 
         nx6620, nx6622, nx6624, nx6626, nx6628, nx6630, nx6632, nx6634, nx6636, 
         nx6638, nx6640, nx6642, nx6644, nx6646, nx6648, nx6650, nx6652, nx6654, 
         nx6656, nx6658, nx6660, nx6662, nx6664, nx6666, nx6668, nx6670, nx6672, 
         nx6674, nx6676, nx6678, nx6680, nx6682, nx6684, nx6686, nx6688, nx6690, 
         nx6692, nx6694, nx6696, nx6698, nx6700, nx6702, nx6704, nx6706, nx6708, 
         nx6710, nx6712, nx6714, nx6716, nx6718, nx6720, nx6722, nx6724, nx6728, 
         nx6730, nx6732, nx6734, nx6736, nx6738, nx6740, nx6742, nx6744, nx6746, 
         nx6748, nx6750, nx6752, nx6754, nx6756, nx6758, nx6760, nx6762, nx6764, 
         nx6766, nx6768, nx6770, nx6772, nx6774, nx6776, nx6778, nx6780, nx6782, 
         nx6784, nx6786, nx6788, nx6790, nx6792, nx6794, nx6796, nx6798, nx6800, 
         nx6802, nx6804, nx6806, nx6808, nx6810, nx6812, nx6814, nx6816, nx6818, 
         nx6820, nx6822, nx6824, nx6826, nx6828, nx6830, nx6832, nx6834, nx6836, 
         nx6838, nx6840, nx6842, nx6844, nx6846, nx6848, nx6850, nx6852, nx6854, 
         nx6856, nx6858, nx6860, nx6862, nx6864, nx6866, nx6868, nx6870, nx6872, 
         nx6874, nx6876, nx6878, nx6880, nx6882, nx6884, nx6886, nx6888, nx6890, 
         nx6892, nx6894, nx6896, nx6898, nx6900, nx6902, nx6904, nx6906, nx6908, 
         nx6910, nx6912, nx6914, nx6916, nx6918, nx6920, nx6922, nx6924, nx6926, 
         nx6928, nx6930, nx6932, nx6934, nx6936, nx6938, nx6940, nx6942, nx6944, 
         nx6946, nx6948, nx6950, nx6952, nx6954, nx6956, nx6958, nx6960, nx6962, 
         nx6964, nx6966, nx6968, nx6970, nx6972, nx6976, nx6978, nx6980, nx6982, 
         nx6984, nx6986, nx6988, nx6990, nx6992, nx6994, nx6996, nx6998, nx7000, 
         nx7002, nx7004, nx7006, nx7008, nx7010, nx7012, nx7014, nx7016, nx7018, 
         nx7020, nx7022, nx7024, nx7026, nx7028, nx7030, nx7032, nx7034, nx7036, 
         nx7038, nx7040, nx7042, nx7044, nx7046, nx7048, nx7050, nx7052, nx7054, 
         nx7056, nx7058, nx7060, nx7062, nx7064, nx7066, nx7068, nx7070, nx7072, 
         nx7074, nx7076, nx7078, nx7080, nx7082, nx7084, nx7086, nx7088, nx7090, 
         nx7092, nx7094, nx7096, nx7098, nx7100, nx7102, nx7104, nx7106, nx7108, 
         nx7110, nx7112, nx7114, nx7116, nx7118, nx7120, nx7122, nx7124, nx7126, 
         nx7128, nx7130, nx7132, nx7134, nx7136, nx7138, nx7140, nx7142, nx7144, 
         nx7146, nx7148, nx7150, nx7152, nx7154, nx7156, nx7158, nx7160, nx7162, 
         nx7164, nx7166, nx7168, nx7170, nx7172, nx7174, nx7176, nx7178, nx7180, 
         nx7182, nx7184, nx7186, nx7188, nx7190, nx7192, nx7194, nx7196, nx7198, 
         nx7200, nx7202, nx7204, nx7206, nx7208, nx7210, nx7212, nx7214, nx7216, 
         nx7218, nx7220, nx7224, nx7226, nx7228, nx7230, nx7232, nx7234, nx7236, 
         nx7238, nx7240, nx7242, nx7244, nx7246, nx7248, nx7250, nx7252, nx7254, 
         nx7256, nx7258, nx7260, nx7262, nx7264, nx7266, nx7268, nx7270, nx7272, 
         nx7274, nx7276, nx7278, nx7280, nx7282, nx7284, nx7286, nx7288, nx7290, 
         nx7292, nx7294, nx7296, nx7298, nx7300, nx7302, nx7304, nx7306, nx7308, 
         nx7310, nx7312, nx7314, nx7316, nx7318, nx7320, nx7322, nx7324, nx7326, 
         nx7328, nx7330, nx7332, nx7334, nx7336, nx7338, nx7340, nx7342, nx7344, 
         nx7346, nx7348, nx7350, nx7352, nx7354, nx7356, nx7358, nx7360, nx7362, 
         nx7364, nx7366, nx7368, nx7370, nx7372, nx7374, nx7376, nx7378, nx7380, 
         nx7382, nx7384, nx7386, nx7388, nx7390, nx7392, nx7394, nx7396, nx7398, 
         nx7400, nx7402, nx7404, nx7406, nx7408, nx7410, nx7412, nx7414, nx7416, 
         nx7418, nx7420, nx7422, nx7424, nx7426, nx7428, nx7430, nx7432, nx7434, 
         nx7436, nx7438, nx7440, nx7442, nx7444, nx7446, nx7448, nx7450, nx7452, 
         nx7454, nx7456, nx7458, nx7460, nx7462, nx7464, nx7466, nx7468, nx7472, 
         nx7474, nx7476, nx7478, nx7480, nx7482, nx7484, nx7486, nx7488, nx7490, 
         nx7492, nx7494, nx7496, nx7498, nx7500, nx7502, nx7504, nx7506, nx7508, 
         nx7510, nx7512, nx7514, nx7516, nx7518, nx7520, nx7522, nx7524, nx7526, 
         nx7528, nx7530, nx7532, nx7534, nx7536, nx7538, nx7540, nx7542, nx7544, 
         nx7546, nx7548, nx7550, nx7552, nx7554, nx7556, nx7558, nx7560, nx7562, 
         nx7564, nx7566, nx7568, nx7570, nx7572, nx7574, nx7576, nx7578, nx7580, 
         nx7582, nx7584, nx7586, nx7588, nx7590, nx7592, nx7594, nx7596, nx7598, 
         nx7600, nx7602, nx7604, nx7606, nx7608, nx7610, nx7612, nx7614, nx7616, 
         nx7618, nx7620, nx7622, nx7624, nx7626, nx7628, nx7630, nx7632, nx7634, 
         nx7636, nx7638, nx7640, nx7642, nx7644, nx7646, nx7648, nx7650, nx7652, 
         nx7654, nx7656, nx7658, nx7660, nx7662, nx7664, nx7666, nx7668, nx7670, 
         nx7672, nx7674, nx7676, nx7678, nx7680, nx7682, nx7684, nx7686, nx7688, 
         nx7690, nx7692, nx7694, nx7696, nx7698, nx7700, nx7702, nx7704, nx7706, 
         nx7708, nx7710, nx7712, nx7714, nx7716, nx7718, nx7720, nx7722, nx7724, 
         nx7726, nx7728, nx7730, nx7732, nx7734, nx7736, nx7738, nx7740, nx7742, 
         nx7744, nx7746, nx7748, nx7750, nx7752, nx7754, nx7756, nx7758, nx7760, 
         nx7762, nx7764, nx7766, nx7768, nx7770, nx7772, nx7774, nx7776, nx7778, 
         nx7780, nx7782, nx7784, nx7786, nx7788, nx7790, nx7792, nx7794, nx7796, 
         nx7798, nx7800, nx7802, nx7804, nx7806, nx7808, nx7810, nx7812, nx7814, 
         nx7816, nx7818, nx7820, nx7822, nx7824, nx7826, nx7828, nx7830, nx7832, 
         nx7834, nx7836, nx7838, nx7840, nx7842, nx7844, nx7846, nx7848, nx7850, 
         nx7852, nx7854, nx7856, nx7858, nx7860, nx7862, nx7864, nx7866, nx7868, 
         nx7870, nx7872, nx7874, nx7876, nx7878, nx7880, nx7882, nx7884, nx7886, 
         nx7888, nx7890, nx7892, nx7894, nx7896, nx7898, nx7900, nx7902, nx7904, 
         nx7906, nx7908, nx7910, nx7912, nx7914, nx7916, nx7918, nx7920, nx7922, 
         nx7924, nx7926, nx7928, nx7930, nx7932, nx7934, nx7936, nx7938, nx7940, 
         nx7942, nx7944, nx7946, nx7948, nx7950, nx7952, nx7954, nx7956, nx7958, 
         nx7960, nx7962, nx7964, nx7966, nx7968, nx7970, nx7972, nx7974, nx7976, 
         nx7978, nx7980, nx7982, nx7984, nx7986, nx7988, nx7990, nx7992, nx7994, 
         nx7996, nx7998, nx8000, nx8002, nx8004, nx8006, nx8008, nx8010, nx8012, 
         nx8014, nx8016, nx8018, nx8020, nx8022, nx8024, nx8026, nx8028, nx8030, 
         nx8032, nx8034, nx8036, nx8038, nx8040, nx8042, nx8044, nx8046, nx8048, 
         nx8050, nx8052, nx8054, nx8056, nx8058, nx8060, nx8062, nx8064, nx8066, 
         nx8068, nx8070, nx8072, nx8074, nx8076, nx8078, nx8080, nx8082, nx8084, 
         nx8086, nx8088, nx8090, nx8092, nx8094, nx8096, nx8098, nx8100, nx8102, 
         nx8104, nx8106, nx8108, nx8110, nx8112, nx8114, nx8116, nx8118, nx8120, 
         nx8122, nx8124, nx8126, nx8128, nx8130, nx8132, nx8134, nx8136, nx8138, 
         nx8140, nx8142, nx8144, nx8146, nx8148, nx8150, nx8152, nx8154, nx8156, 
         nx8158, nx8160, nx8162, nx8164, nx8166, nx8168, nx8170, nx8172, nx8174, 
         nx8176, nx8178, nx8180, nx8182, nx8184, nx8186, nx8188, nx8190, nx8192, 
         nx8194, nx8196, nx8198, nx8200, nx8202, nx8204, nx8206, nx8208, nx8210, 
         nx8212, nx8214, nx8216, nx8218, nx8220, nx8222, nx8224, nx8226, nx8228, 
         nx8230, nx8232, nx8234, nx8236, nx8238, nx8240, nx8242, nx8244, nx8246, 
         nx8248, nx8250, nx8252, nx8254, nx8256, nx8258, nx8260, nx8262, nx8264, 
         nx8266, nx8268, nx8270, nx8272, nx8274, nx8276, nx8278, nx8280, nx8282, 
         nx8284, nx8286, nx8288, nx8290, nx8292, nx8294, nx8296, nx8298, nx8300, 
         nx8302, nx8304, nx8306, nx8308, nx8310, nx8312, nx8314, nx8316, nx8318, 
         nx8320, nx8322, nx8324, nx8326, nx8328, nx8330, nx8332, nx8334, nx8336, 
         nx8338, nx8340, nx8342, nx8344, nx8346, nx8348, nx8350, nx8352, nx8354, 
         nx8356, nx8358, nx8360, nx8362, nx8364, nx8366, nx8368, nx8370, nx8372, 
         nx8374, nx8376, nx8378, nx8380, nx8382, nx8384, nx8386, nx8388, nx8390, 
         nx8392, nx8394, nx8396, nx8398, nx8400, nx8402, nx8404, nx8406, nx8408, 
         nx8410, nx8412, nx8414, nx8416, nx8418, nx8420, nx8422, nx8424, nx8426, 
         nx8428, nx8430, nx8432, nx8434, nx8436, nx8438, nx8440, nx8442, nx8444, 
         nx8446, nx8448, nx8450, nx8452, nx8454, nx8456, nx8458, nx8460, nx8462, 
         nx8464, nx8466, nx8468, nx8470, nx8472, nx8474, nx8476, nx8478, nx8480, 
         nx8482, nx8484, nx8486, nx8488, nx8490, nx8492, nx8494, nx8496, nx8498, 
         nx8500, nx8502, nx8504, nx8506, nx8508, nx8510, nx8512, nx8514, nx8516, 
         nx8518, nx8520, nx8522, nx8524, nx8526, nx8528, nx8530, nx8532, nx8534, 
         nx8536, nx8538, nx8540, nx8542, nx8544, nx8546, nx8548, nx8550, nx8552, 
         nx8554, nx8556, nx8558, nx8560, nx8562, nx8564, nx8566, nx8568, nx8570, 
         nx8572, nx8574, nx8576, nx8578, nx8580, nx8582, nx8584, nx8586, nx8588, 
         nx8590, nx8592, nx8594, nx8596, nx8598, nx8600, nx8602, nx8604, nx8606, 
         nx8608, nx8610, nx8612, nx8614, nx8616, nx8618, nx8620, nx8622, nx8624, 
         nx8626, nx8628, nx8630, nx8632, nx8634, nx8636, nx8638, nx8640, nx8642, 
         nx8644, nx8646, nx8648, nx8650, nx8652, nx8654, nx8656, nx8658, nx8660, 
         nx8662, nx8664, nx8666, nx8668, nx8670, nx8672, nx8674, nx8676, nx8678, 
         nx8680, nx8682, nx8684, nx8686, nx8688, nx8690, nx8692, nx8694, nx8696, 
         nx8698, nx8700, nx8702, nx8704, nx8706, nx8708, nx8710, nx8712, nx8714, 
         nx8716, nx8718, nx8720, nx8722, nx8724, nx8726, nx8728, nx8730, nx8732, 
         nx8734, nx8736, nx8738, nx8740, nx8742, nx8744;
    wire [1278:0] \$dummy ;




    nor02ii ix87 (.Y (CalculatingBooth), .A0 (nx990), .A1 (nx78)) ;
    nor04 ix991 (.Y (nx990), .A0 (CounterOut_0), .A1 (CounterOut_1), .A2 (
          CounterOut_2), .A3 (CounterOut_3)) ;
    nand04 ix79 (.Y (nx78), .A0 (CounterOut_0), .A1 (nx993), .A2 (nx995), .A3 (
           CounterOut_3)) ;
    inv01 ix994 (.Y (nx993), .A (CounterOut_1)) ;
    inv01 ix996 (.Y (nx995), .A (CounterOut_2)) ;
    or02 ix89 (.Y (CounterRST), .A0 (RST), .A1 (Start)) ;
    nor02ii ix999 (.Y (CounterEN), .A0 (Instr), .A1 (nx78)) ;
    oai21 ix29 (.Y (Result[0]), .A0 (nx1001), .A1 (Instr), .B0 (nx1003)) ;
    inv01 ix1002 (.Y (nx1001), .A (L5Results_1__0)) ;
    aoi32 ix1004 (.Y (nx1003), .A0 (L5Results_1__5), .A1 (FilterSize), .A2 (
          Instr), .B0 (L5Results_1__3), .B1 (nx22)) ;
    nor02ii ix23 (.Y (nx22), .A0 (FilterSize), .A1 (Instr)) ;
    oai21 ix41 (.Y (Result[1]), .A0 (nx1007), .A1 (Instr), .B0 (nx1009)) ;
    inv01 ix1008 (.Y (nx1007), .A (L5Results_1__1)) ;
    aoi32 ix1010 (.Y (nx1009), .A0 (L5Results_1__6), .A1 (FilterSize), .A2 (
          Instr), .B0 (L5Results_1__4), .B1 (nx22)) ;
    oai21 ix53 (.Y (Result[2]), .A0 (nx1012), .A1 (Instr), .B0 (nx1014)) ;
    inv01 ix1013 (.Y (nx1012), .A (L5Results_1__2)) ;
    aoi32 ix1015 (.Y (nx1014), .A0 (L5Results_1__7), .A1 (FilterSize), .A2 (
          Instr), .B0 (L5Results_1__5), .B1 (nx22)) ;
    nor02ii ix3 (.Y (Result[5]), .A0 (Instr), .A1 (L5Results_1__5)) ;
    nor02ii ix7 (.Y (Result[6]), .A0 (Instr), .A1 (L5Results_1__6)) ;
    nor02ii ix11 (.Y (Result[7]), .A0 (Instr), .A1 (L5Results_1__7)) ;
    inv01 ix93 (.Y (Done), .A (CounterEN)) ;
    inv01 ix1042 (.Y (nx1043), .A (CalculatingBooth)) ;
    inv02 ix1044 (.Y (CalculatingBooth_dup_1084), .A (nx1043)) ;
    inv02 ix1046 (.Y (CalculatingBooth_dup_1119), .A (nx1043)) ;
    inv02 ix1048 (.Y (CalculatingBooth_dup_1162), .A (nx1043)) ;
    inv01 ix1050 (.Y (CalculatingBooth_dup_1253), .A (nx1043)) ;
    dffr ACCELERATOR_COUNTER_reg_Dout_0 (.Q (CounterOut_0), .QB (\$dummy [0]), .D (
         ACCELERATOR_COUNTER_nx81), .CLK (CLK), .R (CounterRST)) ;
    dffr ACCELERATOR_COUNTER_reg_Dout_1 (.Q (CounterOut_1), .QB (\$dummy [1]), .D (
         ACCELERATOR_COUNTER_nx91), .CLK (CLK), .R (CounterRST)) ;
    xor2 ACCELERATOR_COUNTER_ix7 (.Y (ACCELERATOR_COUNTER_nx6), .A0 (
         CounterOut_1), .A1 (CounterOut_0)) ;
    dffr ACCELERATOR_COUNTER_reg_Dout_2 (.Q (CounterOut_2), .QB (\$dummy [2]), .D (
         ACCELERATOR_COUNTER_nx101), .CLK (CLK), .R (CounterRST)) ;
    xnor2 ACCELERATOR_COUNTER_ix13 (.Y (ACCELERATOR_COUNTER_nx12), .A0 (
          CounterOut_2), .A1 (ACCELERATOR_COUNTER_nx133)) ;
    nand02 ACCELERATOR_COUNTER_ix134 (.Y (ACCELERATOR_COUNTER_nx133), .A0 (
           CounterOut_1), .A1 (CounterOut_0)) ;
    dffr ACCELERATOR_COUNTER_reg_Dout_3 (.Q (CounterOut_3), .QB (\$dummy [3]), .D (
         ACCELERATOR_COUNTER_nx111), .CLK (CLK), .R (CounterRST)) ;
    xnor2 ACCELERATOR_COUNTER_ix19 (.Y (ACCELERATOR_COUNTER_nx18), .A0 (
          CounterOut_3), .A1 (ACCELERATOR_COUNTER_nx139)) ;
    nand03 ACCELERATOR_COUNTER_ix140 (.Y (ACCELERATOR_COUNTER_nx139), .A0 (
           CounterOut_2), .A1 (CounterOut_1), .A2 (CounterOut_0)) ;
    xor2 L1_0_L2_0_G1_MINI_ALU_ix83 (.Y (L1Results_0__0), .A0 (
         L1SecondOperands_0__0), .A1 (L1FirstOperands_0__0)) ;
    xnor2 L1_0_L2_0_G1_MINI_ALU_ix380 (.Y (L1_0_L2_0_G1_MINI_ALU_nx379), .A0 (
          L1_0_L2_0_G1_MINI_ALU_nx381), .A1 (L1_0_L2_0_G1_MINI_ALU_nx383)) ;
    nand02 L1_0_L2_0_G1_MINI_ALU_ix382 (.Y (L1_0_L2_0_G1_MINI_ALU_nx381), .A0 (
           L1_0_L2_0_G1_MINI_ALU_BoothOperand_0), .A1 (nx7562)) ;
    xnor2 L1_0_L2_0_G1_MINI_ALU_ix384 (.Y (L1_0_L2_0_G1_MINI_ALU_nx383), .A0 (
          L1_0_L2_0_G1_MINI_ALU_BoothOperand_1), .A1 (
          L1_0_L2_0_G1_MINI_ALU_BoothP_1)) ;
    inv01 L1_0_L2_0_G1_MINI_ALU_ix388 (.Y (L1_0_L2_0_G1_MINI_ALU_nx387), .A (
          L1_0_L2_0_G1_MINI_ALU_BoothP_2)) ;
    xnor2 L1_0_L2_0_G1_MINI_ALU_ix390 (.Y (L1_0_L2_0_G1_MINI_ALU_nx389), .A0 (
          L1_0_L2_0_G1_MINI_ALU_nx391), .A1 (L1_0_L2_0_G1_MINI_ALU_nx395)) ;
    aoi32 L1_0_L2_0_G1_MINI_ALU_ix392 (.Y (L1_0_L2_0_G1_MINI_ALU_nx391), .A0 (
          L1_0_L2_0_G1_MINI_ALU_BoothOperand_0), .A1 (nx7562), .A2 (
          L1_0_L2_0_G1_MINI_ALU_nx154), .B0 (L1_0_L2_0_G1_MINI_ALU_BoothP_1), .B1 (
          L1_0_L2_0_G1_MINI_ALU_BoothOperand_1)) ;
    xnor2 L1_0_L2_0_G1_MINI_ALU_ix396 (.Y (L1_0_L2_0_G1_MINI_ALU_nx395), .A0 (
          L1_0_L2_0_G1_MINI_ALU_BoothOperand_2), .A1 (
          L1_0_L2_0_G1_MINI_ALU_BoothP_2)) ;
    inv01 L1_0_L2_0_G1_MINI_ALU_ix400 (.Y (L1_0_L2_0_G1_MINI_ALU_nx399), .A (
          L1_0_L2_0_G1_MINI_ALU_BoothP_3)) ;
    xnor2 L1_0_L2_0_G1_MINI_ALU_ix402 (.Y (L1_0_L2_0_G1_MINI_ALU_nx401), .A0 (
          L1_0_L2_0_G1_MINI_ALU_nx403), .A1 (L1_0_L2_0_G1_MINI_ALU_nx405)) ;
    xnor2 L1_0_L2_0_G1_MINI_ALU_ix406 (.Y (L1_0_L2_0_G1_MINI_ALU_nx405), .A0 (
          L1_0_L2_0_G1_MINI_ALU_BoothOperand_3), .A1 (
          L1_0_L2_0_G1_MINI_ALU_BoothP_3)) ;
    inv01 L1_0_L2_0_G1_MINI_ALU_ix410 (.Y (L1_0_L2_0_G1_MINI_ALU_nx409), .A (
          L1_0_L2_0_G1_MINI_ALU_BoothP_4)) ;
    xnor2 L1_0_L2_0_G1_MINI_ALU_ix412 (.Y (L1_0_L2_0_G1_MINI_ALU_nx411), .A0 (
          L1_0_L2_0_G1_MINI_ALU_nx413), .A1 (L1_0_L2_0_G1_MINI_ALU_nx415)) ;
    xnor2 L1_0_L2_0_G1_MINI_ALU_ix416 (.Y (L1_0_L2_0_G1_MINI_ALU_nx415), .A0 (
          L1_0_L2_0_G1_MINI_ALU_BoothOperand_4), .A1 (
          L1_0_L2_0_G1_MINI_ALU_BoothP_4)) ;
    inv01 L1_0_L2_0_G1_MINI_ALU_ix420 (.Y (L1_0_L2_0_G1_MINI_ALU_nx419), .A (
          L1_0_L2_0_G1_MINI_ALU_BoothP_5)) ;
    xnor2 L1_0_L2_0_G1_MINI_ALU_ix422 (.Y (L1_0_L2_0_G1_MINI_ALU_nx421), .A0 (
          L1_0_L2_0_G1_MINI_ALU_nx423), .A1 (L1_0_L2_0_G1_MINI_ALU_nx425)) ;
    xnor2 L1_0_L2_0_G1_MINI_ALU_ix426 (.Y (L1_0_L2_0_G1_MINI_ALU_nx425), .A0 (
          L1_0_L2_0_G1_MINI_ALU_BoothOperand_5), .A1 (
          L1_0_L2_0_G1_MINI_ALU_BoothP_5)) ;
    inv01 L1_0_L2_0_G1_MINI_ALU_ix430 (.Y (L1_0_L2_0_G1_MINI_ALU_nx429), .A (
          L1_0_L2_0_G1_MINI_ALU_BoothP_6)) ;
    xnor2 L1_0_L2_0_G1_MINI_ALU_ix432 (.Y (L1_0_L2_0_G1_MINI_ALU_nx431), .A0 (
          L1_0_L2_0_G1_MINI_ALU_nx433), .A1 (L1_0_L2_0_G1_MINI_ALU_nx435)) ;
    xnor2 L1_0_L2_0_G1_MINI_ALU_ix436 (.Y (L1_0_L2_0_G1_MINI_ALU_nx435), .A0 (
          L1_0_L2_0_G1_MINI_ALU_BoothOperand_6), .A1 (
          L1_0_L2_0_G1_MINI_ALU_BoothP_6)) ;
    inv01 L1_0_L2_0_G1_MINI_ALU_ix440 (.Y (L1_0_L2_0_G1_MINI_ALU_nx439), .A (
          L1_0_L2_0_G1_MINI_ALU_BoothP_7)) ;
    xnor2 L1_0_L2_0_G1_MINI_ALU_ix442 (.Y (L1_0_L2_0_G1_MINI_ALU_nx441), .A0 (
          L1_0_L2_0_G1_MINI_ALU_nx443), .A1 (L1_0_L2_0_G1_MINI_ALU_nx445)) ;
    xnor2 L1_0_L2_0_G1_MINI_ALU_ix446 (.Y (L1_0_L2_0_G1_MINI_ALU_nx445), .A0 (
          L1_0_L2_0_G1_MINI_ALU_BoothOperand_7), .A1 (
          L1_0_L2_0_G1_MINI_ALU_BoothP_7)) ;
    inv01 L1_0_L2_0_G1_MINI_ALU_ix450 (.Y (L1_0_L2_0_G1_MINI_ALU_nx449), .A (
          L1_0_L2_0_G1_MINI_ALU_BoothP_8)) ;
    xnor2 L1_0_L2_0_G1_MINI_ALU_ix452 (.Y (L1_0_L2_0_G1_MINI_ALU_nx451), .A0 (
          L1_0_L2_0_G1_MINI_ALU_nx453), .A1 (L1_0_L2_0_G1_MINI_ALU_nx455)) ;
    xnor2 L1_0_L2_0_G1_MINI_ALU_ix456 (.Y (L1_0_L2_0_G1_MINI_ALU_nx455), .A0 (
          L1_0_L2_0_G1_MINI_ALU_BoothOperand_8), .A1 (
          L1_0_L2_0_G1_MINI_ALU_BoothP_8)) ;
    xor2 L1_0_L2_0_G1_MINI_ALU_ix317 (.Y (L1_0_L2_0_G1_MINI_ALU_nx316), .A0 (
         L1_0_L2_0_G1_MINI_ALU_nx461), .A1 (L1_0_L2_0_G1_MINI_ALU_nx463)) ;
    xnor2 L1_0_L2_0_G1_MINI_ALU_ix464 (.Y (L1_0_L2_0_G1_MINI_ALU_nx463), .A0 (
          L1_0_L2_0_G1_MINI_ALU_BoothOperand_9), .A1 (
          L1_0_L2_0_G1_MINI_ALU_BoothP_9)) ;
    xor2 L1_0_L2_0_G1_MINI_ALU_ix337 (.Y (L1_0_L2_0_G1_MINI_ALU_nx336), .A0 (
         L1_0_L2_0_G1_MINI_ALU_nx467), .A1 (L1_0_L2_0_G1_MINI_ALU_nx471)) ;
    inv01 L1_0_L2_0_G1_MINI_ALU_ix470 (.Y (L1_0_L2_0_G1_MINI_ALU_nx469), .A (
          L1_0_L2_0_G1_MINI_ALU_BoothP_9)) ;
    xnor2 L1_0_L2_0_G1_MINI_ALU_ix472 (.Y (L1_0_L2_0_G1_MINI_ALU_nx471), .A0 (
          L1_0_L2_0_G1_MINI_ALU_BoothOperand_10), .A1 (
          L1_0_L2_0_G1_MINI_ALU_BoothP_10)) ;
    xor2 L1_0_L2_0_G1_MINI_ALU_ix357 (.Y (L1_0_L2_0_G1_MINI_ALU_nx356), .A0 (
         L1_0_L2_0_G1_MINI_ALU_nx475), .A1 (L1_0_L2_0_G1_MINI_ALU_nx479)) ;
    inv01 L1_0_L2_0_G1_MINI_ALU_ix478 (.Y (L1_0_L2_0_G1_MINI_ALU_nx477), .A (
          L1_0_L2_0_G1_MINI_ALU_BoothP_10)) ;
    xnor2 L1_0_L2_0_G1_MINI_ALU_ix480 (.Y (L1_0_L2_0_G1_MINI_ALU_nx479), .A0 (
          L1_0_L2_0_G1_MINI_ALU_BoothOperand_11), .A1 (
          L1_0_L2_0_G1_MINI_ALU_BoothP_11)) ;
    xor2 L1_0_L2_0_G1_MINI_ALU_ix377 (.Y (L1_0_L2_0_G1_MINI_ALU_nx376), .A0 (
         L1_0_L2_0_G1_MINI_ALU_nx483), .A1 (L1_0_L2_0_G1_MINI_ALU_nx487)) ;
    inv01 L1_0_L2_0_G1_MINI_ALU_ix486 (.Y (L1_0_L2_0_G1_MINI_ALU_nx485), .A (
          L1_0_L2_0_G1_MINI_ALU_BoothP_11)) ;
    xnor2 L1_0_L2_0_G1_MINI_ALU_ix488 (.Y (L1_0_L2_0_G1_MINI_ALU_nx487), .A0 (
          L1_0_L2_0_G1_MINI_ALU_BoothOperand_12), .A1 (
          L1_0_L2_0_G1_MINI_ALU_BoothP_12)) ;
    xor2 L1_0_L2_0_G1_MINI_ALU_ix397 (.Y (L1_0_L2_0_G1_MINI_ALU_nx396), .A0 (
         L1_0_L2_0_G1_MINI_ALU_nx491), .A1 (L1_0_L2_0_G1_MINI_ALU_nx495)) ;
    inv01 L1_0_L2_0_G1_MINI_ALU_ix494 (.Y (L1_0_L2_0_G1_MINI_ALU_nx493), .A (
          L1_0_L2_0_G1_MINI_ALU_BoothP_12)) ;
    xnor2 L1_0_L2_0_G1_MINI_ALU_ix496 (.Y (L1_0_L2_0_G1_MINI_ALU_nx495), .A0 (
          L1_0_L2_0_G1_MINI_ALU_BoothOperand_13), .A1 (
          L1_0_L2_0_G1_MINI_ALU_BoothP_13)) ;
    xor2 L1_0_L2_0_G1_MINI_ALU_ix417 (.Y (L1_0_L2_0_G1_MINI_ALU_nx416), .A0 (
         L1_0_L2_0_G1_MINI_ALU_nx499), .A1 (L1_0_L2_0_G1_MINI_ALU_nx503)) ;
    inv01 L1_0_L2_0_G1_MINI_ALU_ix502 (.Y (L1_0_L2_0_G1_MINI_ALU_nx501), .A (
          L1_0_L2_0_G1_MINI_ALU_BoothP_13)) ;
    xnor2 L1_0_L2_0_G1_MINI_ALU_ix504 (.Y (L1_0_L2_0_G1_MINI_ALU_nx503), .A0 (
          L1_0_L2_0_G1_MINI_ALU_BoothOperand_14), .A1 (
          L1_0_L2_0_G1_MINI_ALU_BoothP_14)) ;
    xor2 L1_0_L2_0_G1_MINI_ALU_ix437 (.Y (L1_0_L2_0_G1_MINI_ALU_nx436), .A0 (
         L1_0_L2_0_G1_MINI_ALU_nx507), .A1 (L1_0_L2_0_G1_MINI_ALU_nx511)) ;
    inv01 L1_0_L2_0_G1_MINI_ALU_ix510 (.Y (L1_0_L2_0_G1_MINI_ALU_nx509), .A (
          L1_0_L2_0_G1_MINI_ALU_BoothP_14)) ;
    xnor2 L1_0_L2_0_G1_MINI_ALU_ix512 (.Y (L1_0_L2_0_G1_MINI_ALU_nx511), .A0 (
          L1_0_L2_0_G1_MINI_ALU_BoothOperand_15), .A1 (
          L1_0_L2_0_G1_MINI_ALU_BoothP_15)) ;
    xnor2 L1_0_L2_0_G1_MINI_ALU_ix457 (.Y (L1_0_L2_0_G1_MINI_ALU_nx456), .A0 (
          L1_0_L2_0_G1_MINI_ALU_nx515), .A1 (L1_0_L2_0_G1_MINI_ALU_nx454)) ;
    inv01 L1_0_L2_0_G1_MINI_ALU_ix518 (.Y (L1_0_L2_0_G1_MINI_ALU_nx517), .A (
          L1_0_L2_0_G1_MINI_ALU_BoothP_15)) ;
    xor2 L1_0_L2_0_G1_MINI_ALU_ix455 (.Y (L1_0_L2_0_G1_MINI_ALU_nx454), .A0 (
         L1_0_L2_0_G1_MINI_ALU_BoothOperand_16), .A1 (
         L1_0_L2_0_G1_MINI_ALU_BoothP_16)) ;
    mux21_ni L1_0_L2_0_G1_MINI_ALU_ix91 (.Y (L1SecondOperands_0__0), .A0 (
             L1_0_L2_0_G1_MINI_ALU_BoothP_1), .A1 (WindowDin_0__0__0), .S0 (
             Instr)) ;
    mux21_ni L1_0_L2_0_G1_MINI_ALU_ix99 (.Y (L1SecondOperands_0__1), .A0 (
             L1_0_L2_0_G1_MINI_ALU_BoothP_2), .A1 (WindowDin_0__0__1), .S0 (
             Instr)) ;
    mux21_ni L1_0_L2_0_G1_MINI_ALU_ix107 (.Y (L1SecondOperands_0__2), .A0 (
             L1_0_L2_0_G1_MINI_ALU_BoothP_3), .A1 (WindowDin_0__0__2), .S0 (
             Instr)) ;
    mux21_ni L1_0_L2_0_G1_MINI_ALU_ix115 (.Y (L1SecondOperands_0__3), .A0 (
             L1_0_L2_0_G1_MINI_ALU_BoothP_4), .A1 (WindowDin_0__0__3), .S0 (
             Instr)) ;
    mux21_ni L1_0_L2_0_G1_MINI_ALU_ix123 (.Y (L1SecondOperands_0__4), .A0 (
             L1_0_L2_0_G1_MINI_ALU_BoothP_5), .A1 (WindowDin_0__0__4), .S0 (
             Instr)) ;
    mux21_ni L1_0_L2_0_G1_MINI_ALU_ix131 (.Y (L1SecondOperands_0__5), .A0 (
             L1_0_L2_0_G1_MINI_ALU_BoothP_6), .A1 (WindowDin_0__0__5), .S0 (
             Instr)) ;
    mux21_ni L1_0_L2_0_G1_MINI_ALU_ix139 (.Y (L1SecondOperands_0__6), .A0 (
             L1_0_L2_0_G1_MINI_ALU_BoothP_7), .A1 (WindowDin_0__0__6), .S0 (
             Instr)) ;
    mux21_ni L1_0_L2_0_G1_MINI_ALU_ix147 (.Y (L1SecondOperands_0__7), .A0 (
             L1_0_L2_0_G1_MINI_ALU_BoothP_8), .A1 (WindowDin_0__0__7), .S0 (
             Instr)) ;
    xor2 L1_0_L2_0_G1_MINI_ALU_ix77 (.Y (L1Results_0__1), .A0 (
         L1_0_L2_0_G1_MINI_ALU_nx529), .A1 (L1_0_L2_0_G1_MINI_ALU_nx531)) ;
    nand02 L1_0_L2_0_G1_MINI_ALU_ix530 (.Y (L1_0_L2_0_G1_MINI_ALU_nx529), .A0 (
           L1SecondOperands_0__0), .A1 (L1FirstOperands_0__0)) ;
    xnor2 L1_0_L2_0_G1_MINI_ALU_ix532 (.Y (L1_0_L2_0_G1_MINI_ALU_nx531), .A0 (
          L1SecondOperands_0__1), .A1 (L1FirstOperands_0__1)) ;
    xor2 L1_0_L2_0_G1_MINI_ALU_ix75 (.Y (L1Results_0__2), .A0 (
         L1_0_L2_0_G1_MINI_ALU_nx534), .A1 (L1_0_L2_0_G1_MINI_ALU_nx537)) ;
    aoi32 L1_0_L2_0_G1_MINI_ALU_ix535 (.Y (L1_0_L2_0_G1_MINI_ALU_nx534), .A0 (
          L1SecondOperands_0__0), .A1 (L1FirstOperands_0__0), .A2 (
          L1_0_L2_0_G1_MINI_ALU_nx30), .B0 (L1FirstOperands_0__1), .B1 (
          L1SecondOperands_0__1)) ;
    xnor2 L1_0_L2_0_G1_MINI_ALU_ix538 (.Y (L1_0_L2_0_G1_MINI_ALU_nx537), .A0 (
          L1SecondOperands_0__2), .A1 (L1FirstOperands_0__2)) ;
    xor2 L1_0_L2_0_G1_MINI_ALU_ix73 (.Y (L1Results_0__3), .A0 (
         L1_0_L2_0_G1_MINI_ALU_nx540), .A1 (L1_0_L2_0_G1_MINI_ALU_nx544)) ;
    aoi22 L1_0_L2_0_G1_MINI_ALU_ix541 (.Y (L1_0_L2_0_G1_MINI_ALU_nx540), .A0 (
          L1FirstOperands_0__2), .A1 (L1SecondOperands_0__2), .B0 (
          L1_0_L2_0_G1_MINI_ALU_nx40), .B1 (L1_0_L2_0_G1_MINI_ALU_nx24)) ;
    xnor2 L1_0_L2_0_G1_MINI_ALU_ix545 (.Y (L1_0_L2_0_G1_MINI_ALU_nx544), .A0 (
          L1SecondOperands_0__3), .A1 (L1FirstOperands_0__3)) ;
    xor2 L1_0_L2_0_G1_MINI_ALU_ix71 (.Y (L1Results_0__4), .A0 (
         L1_0_L2_0_G1_MINI_ALU_nx547), .A1 (L1_0_L2_0_G1_MINI_ALU_nx551)) ;
    aoi22 L1_0_L2_0_G1_MINI_ALU_ix548 (.Y (L1_0_L2_0_G1_MINI_ALU_nx547), .A0 (
          L1FirstOperands_0__3), .A1 (L1SecondOperands_0__3), .B0 (
          L1_0_L2_0_G1_MINI_ALU_nx44), .B1 (L1_0_L2_0_G1_MINI_ALU_nx18)) ;
    xnor2 L1_0_L2_0_G1_MINI_ALU_ix552 (.Y (L1_0_L2_0_G1_MINI_ALU_nx551), .A0 (
          L1SecondOperands_0__4), .A1 (L1FirstOperands_0__4)) ;
    xor2 L1_0_L2_0_G1_MINI_ALU_ix69 (.Y (L1Results_0__5), .A0 (
         L1_0_L2_0_G1_MINI_ALU_nx554), .A1 (L1_0_L2_0_G1_MINI_ALU_nx558)) ;
    aoi22 L1_0_L2_0_G1_MINI_ALU_ix555 (.Y (L1_0_L2_0_G1_MINI_ALU_nx554), .A0 (
          L1FirstOperands_0__4), .A1 (L1SecondOperands_0__4), .B0 (
          L1_0_L2_0_G1_MINI_ALU_nx48), .B1 (L1_0_L2_0_G1_MINI_ALU_nx12)) ;
    xnor2 L1_0_L2_0_G1_MINI_ALU_ix559 (.Y (L1_0_L2_0_G1_MINI_ALU_nx558), .A0 (
          L1SecondOperands_0__5), .A1 (L1FirstOperands_0__5)) ;
    xor2 L1_0_L2_0_G1_MINI_ALU_ix67 (.Y (L1Results_0__6), .A0 (
         L1_0_L2_0_G1_MINI_ALU_nx561), .A1 (L1_0_L2_0_G1_MINI_ALU_nx565)) ;
    aoi22 L1_0_L2_0_G1_MINI_ALU_ix562 (.Y (L1_0_L2_0_G1_MINI_ALU_nx561), .A0 (
          L1FirstOperands_0__5), .A1 (L1SecondOperands_0__5), .B0 (
          L1_0_L2_0_G1_MINI_ALU_nx52), .B1 (L1_0_L2_0_G1_MINI_ALU_nx6)) ;
    xnor2 L1_0_L2_0_G1_MINI_ALU_ix566 (.Y (L1_0_L2_0_G1_MINI_ALU_nx565), .A0 (
          L1SecondOperands_0__6), .A1 (L1FirstOperands_0__6)) ;
    xnor2 L1_0_L2_0_G1_MINI_ALU_ix65 (.Y (L1Results_0__7), .A0 (
          L1_0_L2_0_G1_MINI_ALU_nx568), .A1 (L1_0_L2_0_G1_MINI_ALU_nx62)) ;
    aoi22 L1_0_L2_0_G1_MINI_ALU_ix569 (.Y (L1_0_L2_0_G1_MINI_ALU_nx568), .A0 (
          L1FirstOperands_0__6), .A1 (L1SecondOperands_0__6), .B0 (
          L1_0_L2_0_G1_MINI_ALU_nx56), .B1 (L1_0_L2_0_G1_MINI_ALU_nx0)) ;
    xor2 L1_0_L2_0_G1_MINI_ALU_ix63 (.Y (L1_0_L2_0_G1_MINI_ALU_nx62), .A0 (
         L1SecondOperands_0__7), .A1 (L1FirstOperands_0__7)) ;
    inv01 L1_0_L2_0_G1_MINI_ALU_ix155 (.Y (L1_0_L2_0_G1_MINI_ALU_nx154), .A (
          L1_0_L2_0_G1_MINI_ALU_nx383)) ;
    inv01 L1_0_L2_0_G1_MINI_ALU_ix57 (.Y (L1_0_L2_0_G1_MINI_ALU_nx56), .A (
          L1_0_L2_0_G1_MINI_ALU_nx561)) ;
    inv01 L1_0_L2_0_G1_MINI_ALU_ix53 (.Y (L1_0_L2_0_G1_MINI_ALU_nx52), .A (
          L1_0_L2_0_G1_MINI_ALU_nx554)) ;
    inv01 L1_0_L2_0_G1_MINI_ALU_ix49 (.Y (L1_0_L2_0_G1_MINI_ALU_nx48), .A (
          L1_0_L2_0_G1_MINI_ALU_nx547)) ;
    inv01 L1_0_L2_0_G1_MINI_ALU_ix45 (.Y (L1_0_L2_0_G1_MINI_ALU_nx44), .A (
          L1_0_L2_0_G1_MINI_ALU_nx540)) ;
    inv01 L1_0_L2_0_G1_MINI_ALU_ix41 (.Y (L1_0_L2_0_G1_MINI_ALU_nx40), .A (
          L1_0_L2_0_G1_MINI_ALU_nx534)) ;
    inv01 L1_0_L2_0_G1_MINI_ALU_ix31 (.Y (L1_0_L2_0_G1_MINI_ALU_nx30), .A (
          L1_0_L2_0_G1_MINI_ALU_nx531)) ;
    inv01 L1_0_L2_0_G1_MINI_ALU_ix25 (.Y (L1_0_L2_0_G1_MINI_ALU_nx24), .A (
          L1_0_L2_0_G1_MINI_ALU_nx537)) ;
    inv01 L1_0_L2_0_G1_MINI_ALU_ix19 (.Y (L1_0_L2_0_G1_MINI_ALU_nx18), .A (
          L1_0_L2_0_G1_MINI_ALU_nx544)) ;
    inv01 L1_0_L2_0_G1_MINI_ALU_ix13 (.Y (L1_0_L2_0_G1_MINI_ALU_nx12), .A (
          L1_0_L2_0_G1_MINI_ALU_nx551)) ;
    inv01 L1_0_L2_0_G1_MINI_ALU_ix7 (.Y (L1_0_L2_0_G1_MINI_ALU_nx6), .A (
          L1_0_L2_0_G1_MINI_ALU_nx558)) ;
    inv01 L1_0_L2_0_G1_MINI_ALU_ix1 (.Y (L1_0_L2_0_G1_MINI_ALU_nx0), .A (
          L1_0_L2_0_G1_MINI_ALU_nx565)) ;
    fake_gnd L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix216 (.Y (
             L1_0_L2_0_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    nor02ii L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix81 (.Y (
            L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx80), .A0 (Instr), .A1 (Start)) ;
    aoi21 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix77 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_10), .A0 (
          FilterDin_0__0__1), .A1 (FilterDin_0__0__0), .B0 (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx4)) ;
    nor02_2x L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix5 (.Y (
             L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx4), .A0 (FilterDin_0__0__0), .A1 (
             FilterDin_0__0__1)) ;
    aoi21 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix67 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_11), .A0 (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx328), .A1 (FilterDin_0__0__2), .B0 (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx8)) ;
    nor03_2x L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix9 (.Y (
             L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx8), .A0 (FilterDin_0__0__2), .A1 (
             FilterDin_0__0__0), .A2 (FilterDin_0__0__1)) ;
    xnor2 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix59 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_12), .A0 (
          FilterDin_0__0__3), .A1 (L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx8)) ;
    xnor2 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix51 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_13), .A0 (
          FilterDin_0__0__4), .A1 (L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx12)) ;
    nor04 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix13 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx12), .A0 (FilterDin_0__0__3), .A1 (
          FilterDin_0__0__2), .A2 (FilterDin_0__0__0), .A3 (FilterDin_0__0__1)
          ) ;
    xnor2 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix43 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_14), .A0 (
          FilterDin_0__0__5), .A1 (L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx16)) ;
    nor02ii L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix17 (.Y (
            L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx16), .A0 (FilterDin_0__0__4), .A1 (
            L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx12)) ;
    xnor2 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix35 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_15), .A0 (
          FilterDin_0__0__6), .A1 (L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx20)) ;
    nor02ii L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix21 (.Y (
            L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx20), .A0 (FilterDin_0__0__5), .A1 (
            L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx16)) ;
    xnor2 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix27 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_16), .A0 (
          FilterDin_0__0__7), .A1 (L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx24)) ;
    nor02ii L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix25 (.Y (
            L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx24), .A0 (FilterDin_0__0__6), .A1 (
            L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx20)) ;
    inv01 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix329 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx328), .A (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx4)) ;
    inv02 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix383 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx384), .A (
          L1_0_L2_0_G1_MINI_ALU_BoothP_0)) ;
    dff L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_0 (.Q (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_0), .QB (\$dummy [4]), .D (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .CLK (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    inv01 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix565 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx564), .A (RST)) ;
    nor02_2x L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix567 (.Y (
             L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566), .A0 (RST), .A1 (
             L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644)) ;
    dff L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_1 (.Q (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_1), .QB (\$dummy [5]), .D (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .CLK (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_2 (.Q (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_2), .QB (\$dummy [6]), .D (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .CLK (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_3 (.Q (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_3), .QB (\$dummy [7]), .D (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .CLK (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_4 (.Q (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_4), .QB (\$dummy [8]), .D (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .CLK (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_5 (.Q (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_5), .QB (\$dummy [9]), .D (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .CLK (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_6 (.Q (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_6), .QB (\$dummy [10]), .D (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .CLK (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_7 (.Q (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_7), .QB (\$dummy [11]), .D (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .CLK (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_8 (.Q (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_8), .QB (\$dummy [12]), .D (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .CLK (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_9 (.Q (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_9), .QB (\$dummy [13]), .D (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .CLK (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_10 (.Q (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_10), .QB (\$dummy [14]), 
        .D (L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .CLK (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_11 (.Q (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_11), .QB (\$dummy [15]), 
        .D (L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .CLK (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_12 (.Q (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_12), .QB (\$dummy [16]), 
        .D (L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .CLK (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_13 (.Q (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_13), .QB (\$dummy [17]), 
        .D (L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .CLK (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_14 (.Q (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_14), .QB (\$dummy [18]), 
        .D (L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .CLK (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_15 (.Q (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_15), .QB (\$dummy [19]), 
        .D (L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .CLK (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_16 (.Q (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_16), .QB (\$dummy [20]), 
        .D (L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .CLK (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    inv02 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix623 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624), .A (CLK)) ;
    inv02 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix625 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626), .A (CLK)) ;
    inv02 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix627 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628), .A (CLK)) ;
    inv02 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix643 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644), .A (nx7618)) ;
    dff L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_0 (.Q (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_0), .QB (\$dummy [21]), .D (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .CLK (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    nor02_2x L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix567 (.Y (
             L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566), .A0 (RST), .A1 (
             L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644)) ;
    dff L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_1 (.Q (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_1), .QB (\$dummy [22]), .D (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .CLK (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_2 (.Q (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_2), .QB (\$dummy [23]), .D (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .CLK (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_3 (.Q (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_3), .QB (\$dummy [24]), .D (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .CLK (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_4 (.Q (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_4), .QB (\$dummy [25]), .D (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .CLK (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_5 (.Q (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_5), .QB (\$dummy [26]), .D (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .CLK (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_6 (.Q (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_6), .QB (\$dummy [27]), .D (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .CLK (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_7 (.Q (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_7), .QB (\$dummy [28]), .D (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .CLK (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_8 (.Q (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_8), .QB (\$dummy [29]), .D (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .CLK (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_9 (.Q (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_9), .QB (\$dummy [30]), .D (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .CLK (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_10 (.Q (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_10), .QB (\$dummy [31]), 
        .D (L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .CLK (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_11 (.Q (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_11), .QB (\$dummy [32]), 
        .D (L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .CLK (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_12 (.Q (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_12), .QB (\$dummy [33]), 
        .D (L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .CLK (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_13 (.Q (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_13), .QB (\$dummy [34]), 
        .D (L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .CLK (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_14 (.Q (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_14), .QB (\$dummy [35]), 
        .D (L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .CLK (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_15 (.Q (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_15), .QB (\$dummy [36]), 
        .D (L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .CLK (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_16 (.Q (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_16), .QB (\$dummy [37]), 
        .D (L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .CLK (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    inv02 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix623 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624), .A (CLK)) ;
    inv02 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix625 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626), .A (CLK)) ;
    inv02 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix627 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628), .A (CLK)) ;
    inv02 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix643 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644), .A (nx7624)) ;
    dff L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_0 (.Q (
        L1_0_L2_0_G1_MINI_ALU_BoothP_0), .QB (\$dummy [38]), .D (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .CLK (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    nor02_2x L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix567 (.Y (
             L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566), .A0 (RST), .A1 (
             L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    dff L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_1 (.Q (
        L1_0_L2_0_G1_MINI_ALU_BoothP_1), .QB (\$dummy [39]), .D (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .CLK (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_2 (.Q (
        L1_0_L2_0_G1_MINI_ALU_BoothP_2), .QB (\$dummy [40]), .D (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .CLK (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_3 (.Q (
        L1_0_L2_0_G1_MINI_ALU_BoothP_3), .QB (\$dummy [41]), .D (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .CLK (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_4 (.Q (
        L1_0_L2_0_G1_MINI_ALU_BoothP_4), .QB (\$dummy [42]), .D (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .CLK (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_5 (.Q (
        L1_0_L2_0_G1_MINI_ALU_BoothP_5), .QB (\$dummy [43]), .D (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .CLK (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_6 (.Q (
        L1_0_L2_0_G1_MINI_ALU_BoothP_6), .QB (\$dummy [44]), .D (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .CLK (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_7 (.Q (
        L1_0_L2_0_G1_MINI_ALU_BoothP_7), .QB (\$dummy [45]), .D (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .CLK (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_8 (.Q (
        L1_0_L2_0_G1_MINI_ALU_BoothP_8), .QB (\$dummy [46]), .D (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .CLK (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_9 (.Q (
        L1_0_L2_0_G1_MINI_ALU_BoothP_9), .QB (\$dummy [47]), .D (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .CLK (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_10 (.Q (
        L1_0_L2_0_G1_MINI_ALU_BoothP_10), .QB (\$dummy [48]), .D (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .CLK (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_11 (.Q (
        L1_0_L2_0_G1_MINI_ALU_BoothP_11), .QB (\$dummy [49]), .D (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .CLK (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_12 (.Q (
        L1_0_L2_0_G1_MINI_ALU_BoothP_12), .QB (\$dummy [50]), .D (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .CLK (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_13 (.Q (
        L1_0_L2_0_G1_MINI_ALU_BoothP_13), .QB (\$dummy [51]), .D (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .CLK (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_14 (.Q (
        L1_0_L2_0_G1_MINI_ALU_BoothP_14), .QB (\$dummy [52]), .D (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .CLK (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_15 (.Q (
        L1_0_L2_0_G1_MINI_ALU_BoothP_15), .QB (\$dummy [53]), .D (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .CLK (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_16 (.Q (
        L1_0_L2_0_G1_MINI_ALU_BoothP_16), .QB (\$dummy [54]), .D (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .CLK (
        L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    inv02 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix623 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624), .A (CLK)) ;
    inv02 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix625 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626), .A (CLK)) ;
    inv02 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix627 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628), .A (CLK)) ;
    inv02 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix643 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644), .A (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642)) ;
    xor2 L1_0_L2_1_G1_MINI_ALU_ix83 (.Y (L1Results_1__0), .A0 (
         L1SecondOperands_1__0), .A1 (L1FirstOperands_1__0)) ;
    xnor2 L1_0_L2_1_G1_MINI_ALU_ix380 (.Y (L1_0_L2_1_G1_MINI_ALU_nx379), .A0 (
          L1_0_L2_1_G1_MINI_ALU_nx381), .A1 (L1_0_L2_1_G1_MINI_ALU_nx383)) ;
    nand02 L1_0_L2_1_G1_MINI_ALU_ix382 (.Y (L1_0_L2_1_G1_MINI_ALU_nx381), .A0 (
           L1_0_L2_1_G1_MINI_ALU_BoothOperand_0), .A1 (nx7644)) ;
    xnor2 L1_0_L2_1_G1_MINI_ALU_ix384 (.Y (L1_0_L2_1_G1_MINI_ALU_nx383), .A0 (
          L1_0_L2_1_G1_MINI_ALU_BoothOperand_1), .A1 (
          L1_0_L2_1_G1_MINI_ALU_BoothP_1)) ;
    inv01 L1_0_L2_1_G1_MINI_ALU_ix388 (.Y (L1_0_L2_1_G1_MINI_ALU_nx387), .A (
          L1_0_L2_1_G1_MINI_ALU_BoothP_2)) ;
    xnor2 L1_0_L2_1_G1_MINI_ALU_ix390 (.Y (L1_0_L2_1_G1_MINI_ALU_nx389), .A0 (
          L1_0_L2_1_G1_MINI_ALU_nx391), .A1 (L1_0_L2_1_G1_MINI_ALU_nx395)) ;
    aoi32 L1_0_L2_1_G1_MINI_ALU_ix392 (.Y (L1_0_L2_1_G1_MINI_ALU_nx391), .A0 (
          L1_0_L2_1_G1_MINI_ALU_BoothOperand_0), .A1 (nx7644), .A2 (
          L1_0_L2_1_G1_MINI_ALU_nx154), .B0 (L1_0_L2_1_G1_MINI_ALU_BoothP_1), .B1 (
          L1_0_L2_1_G1_MINI_ALU_BoothOperand_1)) ;
    xnor2 L1_0_L2_1_G1_MINI_ALU_ix396 (.Y (L1_0_L2_1_G1_MINI_ALU_nx395), .A0 (
          L1_0_L2_1_G1_MINI_ALU_BoothOperand_2), .A1 (
          L1_0_L2_1_G1_MINI_ALU_BoothP_2)) ;
    inv01 L1_0_L2_1_G1_MINI_ALU_ix400 (.Y (L1_0_L2_1_G1_MINI_ALU_nx399), .A (
          L1_0_L2_1_G1_MINI_ALU_BoothP_3)) ;
    xnor2 L1_0_L2_1_G1_MINI_ALU_ix402 (.Y (L1_0_L2_1_G1_MINI_ALU_nx401), .A0 (
          L1_0_L2_1_G1_MINI_ALU_nx403), .A1 (L1_0_L2_1_G1_MINI_ALU_nx405)) ;
    xnor2 L1_0_L2_1_G1_MINI_ALU_ix406 (.Y (L1_0_L2_1_G1_MINI_ALU_nx405), .A0 (
          L1_0_L2_1_G1_MINI_ALU_BoothOperand_3), .A1 (
          L1_0_L2_1_G1_MINI_ALU_BoothP_3)) ;
    inv01 L1_0_L2_1_G1_MINI_ALU_ix410 (.Y (L1_0_L2_1_G1_MINI_ALU_nx409), .A (
          L1_0_L2_1_G1_MINI_ALU_BoothP_4)) ;
    xnor2 L1_0_L2_1_G1_MINI_ALU_ix412 (.Y (L1_0_L2_1_G1_MINI_ALU_nx411), .A0 (
          L1_0_L2_1_G1_MINI_ALU_nx413), .A1 (L1_0_L2_1_G1_MINI_ALU_nx415)) ;
    xnor2 L1_0_L2_1_G1_MINI_ALU_ix416 (.Y (L1_0_L2_1_G1_MINI_ALU_nx415), .A0 (
          L1_0_L2_1_G1_MINI_ALU_BoothOperand_4), .A1 (
          L1_0_L2_1_G1_MINI_ALU_BoothP_4)) ;
    inv01 L1_0_L2_1_G1_MINI_ALU_ix420 (.Y (L1_0_L2_1_G1_MINI_ALU_nx419), .A (
          L1_0_L2_1_G1_MINI_ALU_BoothP_5)) ;
    xnor2 L1_0_L2_1_G1_MINI_ALU_ix422 (.Y (L1_0_L2_1_G1_MINI_ALU_nx421), .A0 (
          L1_0_L2_1_G1_MINI_ALU_nx423), .A1 (L1_0_L2_1_G1_MINI_ALU_nx425)) ;
    xnor2 L1_0_L2_1_G1_MINI_ALU_ix426 (.Y (L1_0_L2_1_G1_MINI_ALU_nx425), .A0 (
          L1_0_L2_1_G1_MINI_ALU_BoothOperand_5), .A1 (
          L1_0_L2_1_G1_MINI_ALU_BoothP_5)) ;
    inv01 L1_0_L2_1_G1_MINI_ALU_ix430 (.Y (L1_0_L2_1_G1_MINI_ALU_nx429), .A (
          L1_0_L2_1_G1_MINI_ALU_BoothP_6)) ;
    xnor2 L1_0_L2_1_G1_MINI_ALU_ix432 (.Y (L1_0_L2_1_G1_MINI_ALU_nx431), .A0 (
          L1_0_L2_1_G1_MINI_ALU_nx433), .A1 (L1_0_L2_1_G1_MINI_ALU_nx435)) ;
    xnor2 L1_0_L2_1_G1_MINI_ALU_ix436 (.Y (L1_0_L2_1_G1_MINI_ALU_nx435), .A0 (
          L1_0_L2_1_G1_MINI_ALU_BoothOperand_6), .A1 (
          L1_0_L2_1_G1_MINI_ALU_BoothP_6)) ;
    inv01 L1_0_L2_1_G1_MINI_ALU_ix440 (.Y (L1_0_L2_1_G1_MINI_ALU_nx439), .A (
          L1_0_L2_1_G1_MINI_ALU_BoothP_7)) ;
    xnor2 L1_0_L2_1_G1_MINI_ALU_ix442 (.Y (L1_0_L2_1_G1_MINI_ALU_nx441), .A0 (
          L1_0_L2_1_G1_MINI_ALU_nx443), .A1 (L1_0_L2_1_G1_MINI_ALU_nx445)) ;
    xnor2 L1_0_L2_1_G1_MINI_ALU_ix446 (.Y (L1_0_L2_1_G1_MINI_ALU_nx445), .A0 (
          L1_0_L2_1_G1_MINI_ALU_BoothOperand_7), .A1 (
          L1_0_L2_1_G1_MINI_ALU_BoothP_7)) ;
    inv01 L1_0_L2_1_G1_MINI_ALU_ix450 (.Y (L1_0_L2_1_G1_MINI_ALU_nx449), .A (
          L1_0_L2_1_G1_MINI_ALU_BoothP_8)) ;
    xnor2 L1_0_L2_1_G1_MINI_ALU_ix452 (.Y (L1_0_L2_1_G1_MINI_ALU_nx451), .A0 (
          L1_0_L2_1_G1_MINI_ALU_nx453), .A1 (L1_0_L2_1_G1_MINI_ALU_nx455)) ;
    xnor2 L1_0_L2_1_G1_MINI_ALU_ix456 (.Y (L1_0_L2_1_G1_MINI_ALU_nx455), .A0 (
          L1_0_L2_1_G1_MINI_ALU_BoothOperand_8), .A1 (
          L1_0_L2_1_G1_MINI_ALU_BoothP_8)) ;
    xor2 L1_0_L2_1_G1_MINI_ALU_ix317 (.Y (L1_0_L2_1_G1_MINI_ALU_nx316), .A0 (
         L1_0_L2_1_G1_MINI_ALU_nx461), .A1 (L1_0_L2_1_G1_MINI_ALU_nx463)) ;
    xnor2 L1_0_L2_1_G1_MINI_ALU_ix464 (.Y (L1_0_L2_1_G1_MINI_ALU_nx463), .A0 (
          L1_0_L2_1_G1_MINI_ALU_BoothOperand_9), .A1 (
          L1_0_L2_1_G1_MINI_ALU_BoothP_9)) ;
    xor2 L1_0_L2_1_G1_MINI_ALU_ix337 (.Y (L1_0_L2_1_G1_MINI_ALU_nx336), .A0 (
         L1_0_L2_1_G1_MINI_ALU_nx467), .A1 (L1_0_L2_1_G1_MINI_ALU_nx471)) ;
    inv01 L1_0_L2_1_G1_MINI_ALU_ix470 (.Y (L1_0_L2_1_G1_MINI_ALU_nx469), .A (
          L1_0_L2_1_G1_MINI_ALU_BoothP_9)) ;
    xnor2 L1_0_L2_1_G1_MINI_ALU_ix472 (.Y (L1_0_L2_1_G1_MINI_ALU_nx471), .A0 (
          L1_0_L2_1_G1_MINI_ALU_BoothOperand_10), .A1 (
          L1_0_L2_1_G1_MINI_ALU_BoothP_10)) ;
    xor2 L1_0_L2_1_G1_MINI_ALU_ix357 (.Y (L1_0_L2_1_G1_MINI_ALU_nx356), .A0 (
         L1_0_L2_1_G1_MINI_ALU_nx475), .A1 (L1_0_L2_1_G1_MINI_ALU_nx479)) ;
    inv01 L1_0_L2_1_G1_MINI_ALU_ix478 (.Y (L1_0_L2_1_G1_MINI_ALU_nx477), .A (
          L1_0_L2_1_G1_MINI_ALU_BoothP_10)) ;
    xnor2 L1_0_L2_1_G1_MINI_ALU_ix480 (.Y (L1_0_L2_1_G1_MINI_ALU_nx479), .A0 (
          L1_0_L2_1_G1_MINI_ALU_BoothOperand_11), .A1 (
          L1_0_L2_1_G1_MINI_ALU_BoothP_11)) ;
    xor2 L1_0_L2_1_G1_MINI_ALU_ix377 (.Y (L1_0_L2_1_G1_MINI_ALU_nx376), .A0 (
         L1_0_L2_1_G1_MINI_ALU_nx483), .A1 (L1_0_L2_1_G1_MINI_ALU_nx487)) ;
    inv01 L1_0_L2_1_G1_MINI_ALU_ix486 (.Y (L1_0_L2_1_G1_MINI_ALU_nx485), .A (
          L1_0_L2_1_G1_MINI_ALU_BoothP_11)) ;
    xnor2 L1_0_L2_1_G1_MINI_ALU_ix488 (.Y (L1_0_L2_1_G1_MINI_ALU_nx487), .A0 (
          L1_0_L2_1_G1_MINI_ALU_BoothOperand_12), .A1 (
          L1_0_L2_1_G1_MINI_ALU_BoothP_12)) ;
    xor2 L1_0_L2_1_G1_MINI_ALU_ix397 (.Y (L1_0_L2_1_G1_MINI_ALU_nx396), .A0 (
         L1_0_L2_1_G1_MINI_ALU_nx491), .A1 (L1_0_L2_1_G1_MINI_ALU_nx495)) ;
    inv01 L1_0_L2_1_G1_MINI_ALU_ix494 (.Y (L1_0_L2_1_G1_MINI_ALU_nx493), .A (
          L1_0_L2_1_G1_MINI_ALU_BoothP_12)) ;
    xnor2 L1_0_L2_1_G1_MINI_ALU_ix496 (.Y (L1_0_L2_1_G1_MINI_ALU_nx495), .A0 (
          L1_0_L2_1_G1_MINI_ALU_BoothOperand_13), .A1 (
          L1_0_L2_1_G1_MINI_ALU_BoothP_13)) ;
    xor2 L1_0_L2_1_G1_MINI_ALU_ix417 (.Y (L1_0_L2_1_G1_MINI_ALU_nx416), .A0 (
         L1_0_L2_1_G1_MINI_ALU_nx499), .A1 (L1_0_L2_1_G1_MINI_ALU_nx503)) ;
    inv01 L1_0_L2_1_G1_MINI_ALU_ix502 (.Y (L1_0_L2_1_G1_MINI_ALU_nx501), .A (
          L1_0_L2_1_G1_MINI_ALU_BoothP_13)) ;
    xnor2 L1_0_L2_1_G1_MINI_ALU_ix504 (.Y (L1_0_L2_1_G1_MINI_ALU_nx503), .A0 (
          L1_0_L2_1_G1_MINI_ALU_BoothOperand_14), .A1 (
          L1_0_L2_1_G1_MINI_ALU_BoothP_14)) ;
    xor2 L1_0_L2_1_G1_MINI_ALU_ix437 (.Y (L1_0_L2_1_G1_MINI_ALU_nx436), .A0 (
         L1_0_L2_1_G1_MINI_ALU_nx507), .A1 (L1_0_L2_1_G1_MINI_ALU_nx511)) ;
    inv01 L1_0_L2_1_G1_MINI_ALU_ix510 (.Y (L1_0_L2_1_G1_MINI_ALU_nx509), .A (
          L1_0_L2_1_G1_MINI_ALU_BoothP_14)) ;
    xnor2 L1_0_L2_1_G1_MINI_ALU_ix512 (.Y (L1_0_L2_1_G1_MINI_ALU_nx511), .A0 (
          L1_0_L2_1_G1_MINI_ALU_BoothOperand_15), .A1 (
          L1_0_L2_1_G1_MINI_ALU_BoothP_15)) ;
    xnor2 L1_0_L2_1_G1_MINI_ALU_ix457 (.Y (L1_0_L2_1_G1_MINI_ALU_nx456), .A0 (
          L1_0_L2_1_G1_MINI_ALU_nx515), .A1 (L1_0_L2_1_G1_MINI_ALU_nx454)) ;
    inv01 L1_0_L2_1_G1_MINI_ALU_ix518 (.Y (L1_0_L2_1_G1_MINI_ALU_nx517), .A (
          L1_0_L2_1_G1_MINI_ALU_BoothP_15)) ;
    xor2 L1_0_L2_1_G1_MINI_ALU_ix455 (.Y (L1_0_L2_1_G1_MINI_ALU_nx454), .A0 (
         L1_0_L2_1_G1_MINI_ALU_BoothOperand_16), .A1 (
         L1_0_L2_1_G1_MINI_ALU_BoothP_16)) ;
    mux21_ni L1_0_L2_1_G1_MINI_ALU_ix91 (.Y (L1SecondOperands_1__0), .A0 (
             L1_0_L2_1_G1_MINI_ALU_BoothP_1), .A1 (WindowDin_0__1__0), .S0 (
             Instr)) ;
    mux21_ni L1_0_L2_1_G1_MINI_ALU_ix99 (.Y (L1SecondOperands_1__1), .A0 (
             L1_0_L2_1_G1_MINI_ALU_BoothP_2), .A1 (WindowDin_0__1__1), .S0 (
             Instr)) ;
    mux21_ni L1_0_L2_1_G1_MINI_ALU_ix107 (.Y (L1SecondOperands_1__2), .A0 (
             L1_0_L2_1_G1_MINI_ALU_BoothP_3), .A1 (WindowDin_0__1__2), .S0 (
             Instr)) ;
    mux21_ni L1_0_L2_1_G1_MINI_ALU_ix115 (.Y (L1SecondOperands_1__3), .A0 (
             L1_0_L2_1_G1_MINI_ALU_BoothP_4), .A1 (WindowDin_0__1__3), .S0 (
             Instr)) ;
    mux21_ni L1_0_L2_1_G1_MINI_ALU_ix123 (.Y (L1SecondOperands_1__4), .A0 (
             L1_0_L2_1_G1_MINI_ALU_BoothP_5), .A1 (WindowDin_0__1__4), .S0 (
             Instr)) ;
    mux21_ni L1_0_L2_1_G1_MINI_ALU_ix131 (.Y (L1SecondOperands_1__5), .A0 (
             L1_0_L2_1_G1_MINI_ALU_BoothP_6), .A1 (WindowDin_0__1__5), .S0 (
             Instr)) ;
    mux21_ni L1_0_L2_1_G1_MINI_ALU_ix139 (.Y (L1SecondOperands_1__6), .A0 (
             L1_0_L2_1_G1_MINI_ALU_BoothP_7), .A1 (WindowDin_0__1__6), .S0 (
             Instr)) ;
    mux21_ni L1_0_L2_1_G1_MINI_ALU_ix147 (.Y (L1SecondOperands_1__7), .A0 (
             L1_0_L2_1_G1_MINI_ALU_BoothP_8), .A1 (WindowDin_0__1__7), .S0 (
             Instr)) ;
    xor2 L1_0_L2_1_G1_MINI_ALU_ix77 (.Y (L1Results_1__1), .A0 (
         L1_0_L2_1_G1_MINI_ALU_nx529), .A1 (L1_0_L2_1_G1_MINI_ALU_nx531)) ;
    nand02 L1_0_L2_1_G1_MINI_ALU_ix530 (.Y (L1_0_L2_1_G1_MINI_ALU_nx529), .A0 (
           L1SecondOperands_1__0), .A1 (L1FirstOperands_1__0)) ;
    xnor2 L1_0_L2_1_G1_MINI_ALU_ix532 (.Y (L1_0_L2_1_G1_MINI_ALU_nx531), .A0 (
          L1SecondOperands_1__1), .A1 (L1FirstOperands_1__1)) ;
    xor2 L1_0_L2_1_G1_MINI_ALU_ix75 (.Y (L1Results_1__2), .A0 (
         L1_0_L2_1_G1_MINI_ALU_nx534), .A1 (L1_0_L2_1_G1_MINI_ALU_nx537)) ;
    aoi32 L1_0_L2_1_G1_MINI_ALU_ix535 (.Y (L1_0_L2_1_G1_MINI_ALU_nx534), .A0 (
          L1SecondOperands_1__0), .A1 (L1FirstOperands_1__0), .A2 (
          L1_0_L2_1_G1_MINI_ALU_nx30), .B0 (L1FirstOperands_1__1), .B1 (
          L1SecondOperands_1__1)) ;
    xnor2 L1_0_L2_1_G1_MINI_ALU_ix538 (.Y (L1_0_L2_1_G1_MINI_ALU_nx537), .A0 (
          L1SecondOperands_1__2), .A1 (L1FirstOperands_1__2)) ;
    xor2 L1_0_L2_1_G1_MINI_ALU_ix73 (.Y (L1Results_1__3), .A0 (
         L1_0_L2_1_G1_MINI_ALU_nx540), .A1 (L1_0_L2_1_G1_MINI_ALU_nx544)) ;
    aoi22 L1_0_L2_1_G1_MINI_ALU_ix541 (.Y (L1_0_L2_1_G1_MINI_ALU_nx540), .A0 (
          L1FirstOperands_1__2), .A1 (L1SecondOperands_1__2), .B0 (
          L1_0_L2_1_G1_MINI_ALU_nx40), .B1 (L1_0_L2_1_G1_MINI_ALU_nx24)) ;
    xnor2 L1_0_L2_1_G1_MINI_ALU_ix545 (.Y (L1_0_L2_1_G1_MINI_ALU_nx544), .A0 (
          L1SecondOperands_1__3), .A1 (L1FirstOperands_1__3)) ;
    xor2 L1_0_L2_1_G1_MINI_ALU_ix71 (.Y (L1Results_1__4), .A0 (
         L1_0_L2_1_G1_MINI_ALU_nx547), .A1 (L1_0_L2_1_G1_MINI_ALU_nx551)) ;
    aoi22 L1_0_L2_1_G1_MINI_ALU_ix548 (.Y (L1_0_L2_1_G1_MINI_ALU_nx547), .A0 (
          L1FirstOperands_1__3), .A1 (L1SecondOperands_1__3), .B0 (
          L1_0_L2_1_G1_MINI_ALU_nx44), .B1 (L1_0_L2_1_G1_MINI_ALU_nx18)) ;
    xnor2 L1_0_L2_1_G1_MINI_ALU_ix552 (.Y (L1_0_L2_1_G1_MINI_ALU_nx551), .A0 (
          L1SecondOperands_1__4), .A1 (L1FirstOperands_1__4)) ;
    xor2 L1_0_L2_1_G1_MINI_ALU_ix69 (.Y (L1Results_1__5), .A0 (
         L1_0_L2_1_G1_MINI_ALU_nx554), .A1 (L1_0_L2_1_G1_MINI_ALU_nx558)) ;
    aoi22 L1_0_L2_1_G1_MINI_ALU_ix555 (.Y (L1_0_L2_1_G1_MINI_ALU_nx554), .A0 (
          L1FirstOperands_1__4), .A1 (L1SecondOperands_1__4), .B0 (
          L1_0_L2_1_G1_MINI_ALU_nx48), .B1 (L1_0_L2_1_G1_MINI_ALU_nx12)) ;
    xnor2 L1_0_L2_1_G1_MINI_ALU_ix559 (.Y (L1_0_L2_1_G1_MINI_ALU_nx558), .A0 (
          L1SecondOperands_1__5), .A1 (L1FirstOperands_1__5)) ;
    xor2 L1_0_L2_1_G1_MINI_ALU_ix67 (.Y (L1Results_1__6), .A0 (
         L1_0_L2_1_G1_MINI_ALU_nx561), .A1 (L1_0_L2_1_G1_MINI_ALU_nx565)) ;
    aoi22 L1_0_L2_1_G1_MINI_ALU_ix562 (.Y (L1_0_L2_1_G1_MINI_ALU_nx561), .A0 (
          L1FirstOperands_1__5), .A1 (L1SecondOperands_1__5), .B0 (
          L1_0_L2_1_G1_MINI_ALU_nx52), .B1 (L1_0_L2_1_G1_MINI_ALU_nx6)) ;
    xnor2 L1_0_L2_1_G1_MINI_ALU_ix566 (.Y (L1_0_L2_1_G1_MINI_ALU_nx565), .A0 (
          L1SecondOperands_1__6), .A1 (L1FirstOperands_1__6)) ;
    xnor2 L1_0_L2_1_G1_MINI_ALU_ix65 (.Y (L1Results_1__7), .A0 (
          L1_0_L2_1_G1_MINI_ALU_nx568), .A1 (L1_0_L2_1_G1_MINI_ALU_nx62)) ;
    aoi22 L1_0_L2_1_G1_MINI_ALU_ix569 (.Y (L1_0_L2_1_G1_MINI_ALU_nx568), .A0 (
          L1FirstOperands_1__6), .A1 (L1SecondOperands_1__6), .B0 (
          L1_0_L2_1_G1_MINI_ALU_nx56), .B1 (L1_0_L2_1_G1_MINI_ALU_nx0)) ;
    xor2 L1_0_L2_1_G1_MINI_ALU_ix63 (.Y (L1_0_L2_1_G1_MINI_ALU_nx62), .A0 (
         L1SecondOperands_1__7), .A1 (L1FirstOperands_1__7)) ;
    inv01 L1_0_L2_1_G1_MINI_ALU_ix155 (.Y (L1_0_L2_1_G1_MINI_ALU_nx154), .A (
          L1_0_L2_1_G1_MINI_ALU_nx383)) ;
    inv01 L1_0_L2_1_G1_MINI_ALU_ix57 (.Y (L1_0_L2_1_G1_MINI_ALU_nx56), .A (
          L1_0_L2_1_G1_MINI_ALU_nx561)) ;
    inv01 L1_0_L2_1_G1_MINI_ALU_ix53 (.Y (L1_0_L2_1_G1_MINI_ALU_nx52), .A (
          L1_0_L2_1_G1_MINI_ALU_nx554)) ;
    inv01 L1_0_L2_1_G1_MINI_ALU_ix49 (.Y (L1_0_L2_1_G1_MINI_ALU_nx48), .A (
          L1_0_L2_1_G1_MINI_ALU_nx547)) ;
    inv01 L1_0_L2_1_G1_MINI_ALU_ix45 (.Y (L1_0_L2_1_G1_MINI_ALU_nx44), .A (
          L1_0_L2_1_G1_MINI_ALU_nx540)) ;
    inv01 L1_0_L2_1_G1_MINI_ALU_ix41 (.Y (L1_0_L2_1_G1_MINI_ALU_nx40), .A (
          L1_0_L2_1_G1_MINI_ALU_nx534)) ;
    inv01 L1_0_L2_1_G1_MINI_ALU_ix31 (.Y (L1_0_L2_1_G1_MINI_ALU_nx30), .A (
          L1_0_L2_1_G1_MINI_ALU_nx531)) ;
    inv01 L1_0_L2_1_G1_MINI_ALU_ix25 (.Y (L1_0_L2_1_G1_MINI_ALU_nx24), .A (
          L1_0_L2_1_G1_MINI_ALU_nx537)) ;
    inv01 L1_0_L2_1_G1_MINI_ALU_ix19 (.Y (L1_0_L2_1_G1_MINI_ALU_nx18), .A (
          L1_0_L2_1_G1_MINI_ALU_nx544)) ;
    inv01 L1_0_L2_1_G1_MINI_ALU_ix13 (.Y (L1_0_L2_1_G1_MINI_ALU_nx12), .A (
          L1_0_L2_1_G1_MINI_ALU_nx551)) ;
    inv01 L1_0_L2_1_G1_MINI_ALU_ix7 (.Y (L1_0_L2_1_G1_MINI_ALU_nx6), .A (
          L1_0_L2_1_G1_MINI_ALU_nx558)) ;
    inv01 L1_0_L2_1_G1_MINI_ALU_ix1 (.Y (L1_0_L2_1_G1_MINI_ALU_nx0), .A (
          L1_0_L2_1_G1_MINI_ALU_nx565)) ;
    fake_gnd L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix216 (.Y (
             L1_0_L2_1_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    nor02ii L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix81 (.Y (
            L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx80), .A0 (Instr), .A1 (Start)) ;
    aoi21 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix77 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_10), .A0 (
          FilterDin_0__1__1), .A1 (FilterDin_0__1__0), .B0 (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx4)) ;
    nor02_2x L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix5 (.Y (
             L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx4), .A0 (FilterDin_0__1__0), .A1 (
             FilterDin_0__1__1)) ;
    aoi21 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix67 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_11), .A0 (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx328), .A1 (FilterDin_0__1__2), .B0 (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx8)) ;
    nor03_2x L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix9 (.Y (
             L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx8), .A0 (FilterDin_0__1__2), .A1 (
             FilterDin_0__1__0), .A2 (FilterDin_0__1__1)) ;
    xnor2 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix59 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_12), .A0 (
          FilterDin_0__1__3), .A1 (L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx8)) ;
    xnor2 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix51 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_13), .A0 (
          FilterDin_0__1__4), .A1 (L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx12)) ;
    nor04 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix13 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx12), .A0 (FilterDin_0__1__3), .A1 (
          FilterDin_0__1__2), .A2 (FilterDin_0__1__0), .A3 (FilterDin_0__1__1)
          ) ;
    xnor2 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix43 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_14), .A0 (
          FilterDin_0__1__5), .A1 (L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx16)) ;
    nor02ii L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix17 (.Y (
            L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx16), .A0 (FilterDin_0__1__4), .A1 (
            L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx12)) ;
    xnor2 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix35 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_15), .A0 (
          FilterDin_0__1__6), .A1 (L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx20)) ;
    nor02ii L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix21 (.Y (
            L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx20), .A0 (FilterDin_0__1__5), .A1 (
            L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx16)) ;
    xnor2 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix27 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_16), .A0 (
          FilterDin_0__1__7), .A1 (L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx24)) ;
    nor02ii L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix25 (.Y (
            L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx24), .A0 (FilterDin_0__1__6), .A1 (
            L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx20)) ;
    inv01 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix329 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx328), .A (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx4)) ;
    inv02 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix383 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx384), .A (
          L1_0_L2_1_G1_MINI_ALU_BoothP_0)) ;
    dff L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_0 (.Q (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_0), .QB (\$dummy [55]), .D (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .CLK (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    nor02_2x L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix567 (.Y (
             L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566), .A0 (RST), .A1 (
             L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644)) ;
    dff L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_1 (.Q (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_1), .QB (\$dummy [56]), .D (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .CLK (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_2 (.Q (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_2), .QB (\$dummy [57]), .D (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .CLK (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_3 (.Q (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_3), .QB (\$dummy [58]), .D (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .CLK (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_4 (.Q (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_4), .QB (\$dummy [59]), .D (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .CLK (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_5 (.Q (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_5), .QB (\$dummy [60]), .D (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .CLK (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_6 (.Q (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_6), .QB (\$dummy [61]), .D (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .CLK (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_7 (.Q (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_7), .QB (\$dummy [62]), .D (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .CLK (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_8 (.Q (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_8), .QB (\$dummy [63]), .D (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .CLK (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_9 (.Q (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_9), .QB (\$dummy [64]), .D (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .CLK (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_10 (.Q (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_10), .QB (\$dummy [65]), 
        .D (L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .CLK (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_11 (.Q (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_11), .QB (\$dummy [66]), 
        .D (L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .CLK (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_12 (.Q (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_12), .QB (\$dummy [67]), 
        .D (L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .CLK (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_13 (.Q (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_13), .QB (\$dummy [68]), 
        .D (L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .CLK (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_14 (.Q (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_14), .QB (\$dummy [69]), 
        .D (L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .CLK (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_15 (.Q (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_15), .QB (\$dummy [70]), 
        .D (L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .CLK (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_16 (.Q (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_16), .QB (\$dummy [71]), 
        .D (L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .CLK (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    inv02 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix623 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624), .A (CLK)) ;
    inv02 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix625 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626), .A (CLK)) ;
    inv02 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix627 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628), .A (CLK)) ;
    inv02 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix643 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644), .A (nx7658)) ;
    dff L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_0 (.Q (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_0), .QB (\$dummy [72]), .D (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .CLK (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    nor02_2x L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix567 (.Y (
             L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566), .A0 (RST), .A1 (
             L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644)) ;
    dff L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_1 (.Q (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_1), .QB (\$dummy [73]), .D (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .CLK (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_2 (.Q (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_2), .QB (\$dummy [74]), .D (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .CLK (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_3 (.Q (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_3), .QB (\$dummy [75]), .D (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .CLK (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_4 (.Q (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_4), .QB (\$dummy [76]), .D (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .CLK (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_5 (.Q (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_5), .QB (\$dummy [77]), .D (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .CLK (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_6 (.Q (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_6), .QB (\$dummy [78]), .D (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .CLK (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_7 (.Q (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_7), .QB (\$dummy [79]), .D (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .CLK (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_8 (.Q (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_8), .QB (\$dummy [80]), .D (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .CLK (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_9 (.Q (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_9), .QB (\$dummy [81]), .D (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .CLK (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_10 (.Q (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_10), .QB (\$dummy [82]), 
        .D (L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .CLK (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_11 (.Q (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_11), .QB (\$dummy [83]), 
        .D (L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .CLK (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_12 (.Q (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_12), .QB (\$dummy [84]), 
        .D (L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .CLK (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_13 (.Q (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_13), .QB (\$dummy [85]), 
        .D (L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .CLK (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_14 (.Q (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_14), .QB (\$dummy [86]), 
        .D (L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .CLK (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_15 (.Q (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_15), .QB (\$dummy [87]), 
        .D (L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .CLK (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_16 (.Q (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_16), .QB (\$dummy [88]), 
        .D (L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .CLK (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    inv02 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix623 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624), .A (CLK)) ;
    inv02 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix625 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626), .A (CLK)) ;
    inv02 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix627 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628), .A (CLK)) ;
    inv02 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix643 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644), .A (nx7664)) ;
    dff L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_0 (.Q (
        L1_0_L2_1_G1_MINI_ALU_BoothP_0), .QB (\$dummy [89]), .D (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .CLK (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    nor02_2x L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix567 (.Y (
             L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566), .A0 (RST), .A1 (
             L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    dff L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_1 (.Q (
        L1_0_L2_1_G1_MINI_ALU_BoothP_1), .QB (\$dummy [90]), .D (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .CLK (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_2 (.Q (
        L1_0_L2_1_G1_MINI_ALU_BoothP_2), .QB (\$dummy [91]), .D (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .CLK (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_3 (.Q (
        L1_0_L2_1_G1_MINI_ALU_BoothP_3), .QB (\$dummy [92]), .D (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .CLK (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_4 (.Q (
        L1_0_L2_1_G1_MINI_ALU_BoothP_4), .QB (\$dummy [93]), .D (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .CLK (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_5 (.Q (
        L1_0_L2_1_G1_MINI_ALU_BoothP_5), .QB (\$dummy [94]), .D (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .CLK (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_6 (.Q (
        L1_0_L2_1_G1_MINI_ALU_BoothP_6), .QB (\$dummy [95]), .D (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .CLK (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_7 (.Q (
        L1_0_L2_1_G1_MINI_ALU_BoothP_7), .QB (\$dummy [96]), .D (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .CLK (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_8 (.Q (
        L1_0_L2_1_G1_MINI_ALU_BoothP_8), .QB (\$dummy [97]), .D (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .CLK (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_9 (.Q (
        L1_0_L2_1_G1_MINI_ALU_BoothP_9), .QB (\$dummy [98]), .D (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .CLK (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_10 (.Q (
        L1_0_L2_1_G1_MINI_ALU_BoothP_10), .QB (\$dummy [99]), .D (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .CLK (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_11 (.Q (
        L1_0_L2_1_G1_MINI_ALU_BoothP_11), .QB (\$dummy [100]), .D (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .CLK (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_12 (.Q (
        L1_0_L2_1_G1_MINI_ALU_BoothP_12), .QB (\$dummy [101]), .D (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .CLK (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_13 (.Q (
        L1_0_L2_1_G1_MINI_ALU_BoothP_13), .QB (\$dummy [102]), .D (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .CLK (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_14 (.Q (
        L1_0_L2_1_G1_MINI_ALU_BoothP_14), .QB (\$dummy [103]), .D (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .CLK (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_15 (.Q (
        L1_0_L2_1_G1_MINI_ALU_BoothP_15), .QB (\$dummy [104]), .D (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .CLK (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_16 (.Q (
        L1_0_L2_1_G1_MINI_ALU_BoothP_16), .QB (\$dummy [105]), .D (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .CLK (
        L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    inv02 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix623 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624), .A (CLK)) ;
    inv02 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix625 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626), .A (CLK)) ;
    inv02 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix627 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628), .A (CLK)) ;
    inv02 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix643 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644), .A (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642)) ;
    xor2 L1_0_L2_2_G1_MINI_ALU_ix83 (.Y (L1Results_2__0), .A0 (
         L1SecondOperands_2__0), .A1 (L1FirstOperands_2__0)) ;
    xnor2 L1_0_L2_2_G1_MINI_ALU_ix380 (.Y (L1_0_L2_2_G1_MINI_ALU_nx379), .A0 (
          L1_0_L2_2_G1_MINI_ALU_nx381), .A1 (L1_0_L2_2_G1_MINI_ALU_nx383)) ;
    nand02 L1_0_L2_2_G1_MINI_ALU_ix382 (.Y (L1_0_L2_2_G1_MINI_ALU_nx381), .A0 (
           L1_0_L2_2_G1_MINI_ALU_BoothOperand_0), .A1 (nx7684)) ;
    xnor2 L1_0_L2_2_G1_MINI_ALU_ix384 (.Y (L1_0_L2_2_G1_MINI_ALU_nx383), .A0 (
          L1_0_L2_2_G1_MINI_ALU_BoothOperand_1), .A1 (
          L1_0_L2_2_G1_MINI_ALU_BoothP_1)) ;
    inv01 L1_0_L2_2_G1_MINI_ALU_ix388 (.Y (L1_0_L2_2_G1_MINI_ALU_nx387), .A (
          L1_0_L2_2_G1_MINI_ALU_BoothP_2)) ;
    xnor2 L1_0_L2_2_G1_MINI_ALU_ix390 (.Y (L1_0_L2_2_G1_MINI_ALU_nx389), .A0 (
          L1_0_L2_2_G1_MINI_ALU_nx391), .A1 (L1_0_L2_2_G1_MINI_ALU_nx395)) ;
    aoi32 L1_0_L2_2_G1_MINI_ALU_ix392 (.Y (L1_0_L2_2_G1_MINI_ALU_nx391), .A0 (
          L1_0_L2_2_G1_MINI_ALU_BoothOperand_0), .A1 (nx7684), .A2 (
          L1_0_L2_2_G1_MINI_ALU_nx154), .B0 (L1_0_L2_2_G1_MINI_ALU_BoothP_1), .B1 (
          L1_0_L2_2_G1_MINI_ALU_BoothOperand_1)) ;
    xnor2 L1_0_L2_2_G1_MINI_ALU_ix396 (.Y (L1_0_L2_2_G1_MINI_ALU_nx395), .A0 (
          L1_0_L2_2_G1_MINI_ALU_BoothOperand_2), .A1 (
          L1_0_L2_2_G1_MINI_ALU_BoothP_2)) ;
    inv01 L1_0_L2_2_G1_MINI_ALU_ix400 (.Y (L1_0_L2_2_G1_MINI_ALU_nx399), .A (
          L1_0_L2_2_G1_MINI_ALU_BoothP_3)) ;
    xnor2 L1_0_L2_2_G1_MINI_ALU_ix402 (.Y (L1_0_L2_2_G1_MINI_ALU_nx401), .A0 (
          L1_0_L2_2_G1_MINI_ALU_nx403), .A1 (L1_0_L2_2_G1_MINI_ALU_nx405)) ;
    xnor2 L1_0_L2_2_G1_MINI_ALU_ix406 (.Y (L1_0_L2_2_G1_MINI_ALU_nx405), .A0 (
          L1_0_L2_2_G1_MINI_ALU_BoothOperand_3), .A1 (
          L1_0_L2_2_G1_MINI_ALU_BoothP_3)) ;
    inv01 L1_0_L2_2_G1_MINI_ALU_ix410 (.Y (L1_0_L2_2_G1_MINI_ALU_nx409), .A (
          L1_0_L2_2_G1_MINI_ALU_BoothP_4)) ;
    xnor2 L1_0_L2_2_G1_MINI_ALU_ix412 (.Y (L1_0_L2_2_G1_MINI_ALU_nx411), .A0 (
          L1_0_L2_2_G1_MINI_ALU_nx413), .A1 (L1_0_L2_2_G1_MINI_ALU_nx415)) ;
    xnor2 L1_0_L2_2_G1_MINI_ALU_ix416 (.Y (L1_0_L2_2_G1_MINI_ALU_nx415), .A0 (
          L1_0_L2_2_G1_MINI_ALU_BoothOperand_4), .A1 (
          L1_0_L2_2_G1_MINI_ALU_BoothP_4)) ;
    inv01 L1_0_L2_2_G1_MINI_ALU_ix420 (.Y (L1_0_L2_2_G1_MINI_ALU_nx419), .A (
          L1_0_L2_2_G1_MINI_ALU_BoothP_5)) ;
    xnor2 L1_0_L2_2_G1_MINI_ALU_ix422 (.Y (L1_0_L2_2_G1_MINI_ALU_nx421), .A0 (
          L1_0_L2_2_G1_MINI_ALU_nx423), .A1 (L1_0_L2_2_G1_MINI_ALU_nx425)) ;
    xnor2 L1_0_L2_2_G1_MINI_ALU_ix426 (.Y (L1_0_L2_2_G1_MINI_ALU_nx425), .A0 (
          L1_0_L2_2_G1_MINI_ALU_BoothOperand_5), .A1 (
          L1_0_L2_2_G1_MINI_ALU_BoothP_5)) ;
    inv01 L1_0_L2_2_G1_MINI_ALU_ix430 (.Y (L1_0_L2_2_G1_MINI_ALU_nx429), .A (
          L1_0_L2_2_G1_MINI_ALU_BoothP_6)) ;
    xnor2 L1_0_L2_2_G1_MINI_ALU_ix432 (.Y (L1_0_L2_2_G1_MINI_ALU_nx431), .A0 (
          L1_0_L2_2_G1_MINI_ALU_nx433), .A1 (L1_0_L2_2_G1_MINI_ALU_nx435)) ;
    xnor2 L1_0_L2_2_G1_MINI_ALU_ix436 (.Y (L1_0_L2_2_G1_MINI_ALU_nx435), .A0 (
          L1_0_L2_2_G1_MINI_ALU_BoothOperand_6), .A1 (
          L1_0_L2_2_G1_MINI_ALU_BoothP_6)) ;
    inv01 L1_0_L2_2_G1_MINI_ALU_ix440 (.Y (L1_0_L2_2_G1_MINI_ALU_nx439), .A (
          L1_0_L2_2_G1_MINI_ALU_BoothP_7)) ;
    xnor2 L1_0_L2_2_G1_MINI_ALU_ix442 (.Y (L1_0_L2_2_G1_MINI_ALU_nx441), .A0 (
          L1_0_L2_2_G1_MINI_ALU_nx443), .A1 (L1_0_L2_2_G1_MINI_ALU_nx445)) ;
    xnor2 L1_0_L2_2_G1_MINI_ALU_ix446 (.Y (L1_0_L2_2_G1_MINI_ALU_nx445), .A0 (
          L1_0_L2_2_G1_MINI_ALU_BoothOperand_7), .A1 (
          L1_0_L2_2_G1_MINI_ALU_BoothP_7)) ;
    inv01 L1_0_L2_2_G1_MINI_ALU_ix450 (.Y (L1_0_L2_2_G1_MINI_ALU_nx449), .A (
          L1_0_L2_2_G1_MINI_ALU_BoothP_8)) ;
    xnor2 L1_0_L2_2_G1_MINI_ALU_ix452 (.Y (L1_0_L2_2_G1_MINI_ALU_nx451), .A0 (
          L1_0_L2_2_G1_MINI_ALU_nx453), .A1 (L1_0_L2_2_G1_MINI_ALU_nx455)) ;
    xnor2 L1_0_L2_2_G1_MINI_ALU_ix456 (.Y (L1_0_L2_2_G1_MINI_ALU_nx455), .A0 (
          L1_0_L2_2_G1_MINI_ALU_BoothOperand_8), .A1 (
          L1_0_L2_2_G1_MINI_ALU_BoothP_8)) ;
    xor2 L1_0_L2_2_G1_MINI_ALU_ix317 (.Y (L1_0_L2_2_G1_MINI_ALU_nx316), .A0 (
         L1_0_L2_2_G1_MINI_ALU_nx461), .A1 (L1_0_L2_2_G1_MINI_ALU_nx463)) ;
    xnor2 L1_0_L2_2_G1_MINI_ALU_ix464 (.Y (L1_0_L2_2_G1_MINI_ALU_nx463), .A0 (
          L1_0_L2_2_G1_MINI_ALU_BoothOperand_9), .A1 (
          L1_0_L2_2_G1_MINI_ALU_BoothP_9)) ;
    xor2 L1_0_L2_2_G1_MINI_ALU_ix337 (.Y (L1_0_L2_2_G1_MINI_ALU_nx336), .A0 (
         L1_0_L2_2_G1_MINI_ALU_nx467), .A1 (L1_0_L2_2_G1_MINI_ALU_nx471)) ;
    inv01 L1_0_L2_2_G1_MINI_ALU_ix470 (.Y (L1_0_L2_2_G1_MINI_ALU_nx469), .A (
          L1_0_L2_2_G1_MINI_ALU_BoothP_9)) ;
    xnor2 L1_0_L2_2_G1_MINI_ALU_ix472 (.Y (L1_0_L2_2_G1_MINI_ALU_nx471), .A0 (
          L1_0_L2_2_G1_MINI_ALU_BoothOperand_10), .A1 (
          L1_0_L2_2_G1_MINI_ALU_BoothP_10)) ;
    xor2 L1_0_L2_2_G1_MINI_ALU_ix357 (.Y (L1_0_L2_2_G1_MINI_ALU_nx356), .A0 (
         L1_0_L2_2_G1_MINI_ALU_nx475), .A1 (L1_0_L2_2_G1_MINI_ALU_nx479)) ;
    inv01 L1_0_L2_2_G1_MINI_ALU_ix478 (.Y (L1_0_L2_2_G1_MINI_ALU_nx477), .A (
          L1_0_L2_2_G1_MINI_ALU_BoothP_10)) ;
    xnor2 L1_0_L2_2_G1_MINI_ALU_ix480 (.Y (L1_0_L2_2_G1_MINI_ALU_nx479), .A0 (
          L1_0_L2_2_G1_MINI_ALU_BoothOperand_11), .A1 (
          L1_0_L2_2_G1_MINI_ALU_BoothP_11)) ;
    xor2 L1_0_L2_2_G1_MINI_ALU_ix377 (.Y (L1_0_L2_2_G1_MINI_ALU_nx376), .A0 (
         L1_0_L2_2_G1_MINI_ALU_nx483), .A1 (L1_0_L2_2_G1_MINI_ALU_nx487)) ;
    inv01 L1_0_L2_2_G1_MINI_ALU_ix486 (.Y (L1_0_L2_2_G1_MINI_ALU_nx485), .A (
          L1_0_L2_2_G1_MINI_ALU_BoothP_11)) ;
    xnor2 L1_0_L2_2_G1_MINI_ALU_ix488 (.Y (L1_0_L2_2_G1_MINI_ALU_nx487), .A0 (
          L1_0_L2_2_G1_MINI_ALU_BoothOperand_12), .A1 (
          L1_0_L2_2_G1_MINI_ALU_BoothP_12)) ;
    xor2 L1_0_L2_2_G1_MINI_ALU_ix397 (.Y (L1_0_L2_2_G1_MINI_ALU_nx396), .A0 (
         L1_0_L2_2_G1_MINI_ALU_nx491), .A1 (L1_0_L2_2_G1_MINI_ALU_nx495)) ;
    inv01 L1_0_L2_2_G1_MINI_ALU_ix494 (.Y (L1_0_L2_2_G1_MINI_ALU_nx493), .A (
          L1_0_L2_2_G1_MINI_ALU_BoothP_12)) ;
    xnor2 L1_0_L2_2_G1_MINI_ALU_ix496 (.Y (L1_0_L2_2_G1_MINI_ALU_nx495), .A0 (
          L1_0_L2_2_G1_MINI_ALU_BoothOperand_13), .A1 (
          L1_0_L2_2_G1_MINI_ALU_BoothP_13)) ;
    xor2 L1_0_L2_2_G1_MINI_ALU_ix417 (.Y (L1_0_L2_2_G1_MINI_ALU_nx416), .A0 (
         L1_0_L2_2_G1_MINI_ALU_nx499), .A1 (L1_0_L2_2_G1_MINI_ALU_nx503)) ;
    inv01 L1_0_L2_2_G1_MINI_ALU_ix502 (.Y (L1_0_L2_2_G1_MINI_ALU_nx501), .A (
          L1_0_L2_2_G1_MINI_ALU_BoothP_13)) ;
    xnor2 L1_0_L2_2_G1_MINI_ALU_ix504 (.Y (L1_0_L2_2_G1_MINI_ALU_nx503), .A0 (
          L1_0_L2_2_G1_MINI_ALU_BoothOperand_14), .A1 (
          L1_0_L2_2_G1_MINI_ALU_BoothP_14)) ;
    xor2 L1_0_L2_2_G1_MINI_ALU_ix437 (.Y (L1_0_L2_2_G1_MINI_ALU_nx436), .A0 (
         L1_0_L2_2_G1_MINI_ALU_nx507), .A1 (L1_0_L2_2_G1_MINI_ALU_nx511)) ;
    inv01 L1_0_L2_2_G1_MINI_ALU_ix510 (.Y (L1_0_L2_2_G1_MINI_ALU_nx509), .A (
          L1_0_L2_2_G1_MINI_ALU_BoothP_14)) ;
    xnor2 L1_0_L2_2_G1_MINI_ALU_ix512 (.Y (L1_0_L2_2_G1_MINI_ALU_nx511), .A0 (
          L1_0_L2_2_G1_MINI_ALU_BoothOperand_15), .A1 (
          L1_0_L2_2_G1_MINI_ALU_BoothP_15)) ;
    xnor2 L1_0_L2_2_G1_MINI_ALU_ix457 (.Y (L1_0_L2_2_G1_MINI_ALU_nx456), .A0 (
          L1_0_L2_2_G1_MINI_ALU_nx515), .A1 (L1_0_L2_2_G1_MINI_ALU_nx454)) ;
    inv01 L1_0_L2_2_G1_MINI_ALU_ix518 (.Y (L1_0_L2_2_G1_MINI_ALU_nx517), .A (
          L1_0_L2_2_G1_MINI_ALU_BoothP_15)) ;
    xor2 L1_0_L2_2_G1_MINI_ALU_ix455 (.Y (L1_0_L2_2_G1_MINI_ALU_nx454), .A0 (
         L1_0_L2_2_G1_MINI_ALU_BoothOperand_16), .A1 (
         L1_0_L2_2_G1_MINI_ALU_BoothP_16)) ;
    mux21_ni L1_0_L2_2_G1_MINI_ALU_ix91 (.Y (L1SecondOperands_2__0), .A0 (
             L1_0_L2_2_G1_MINI_ALU_BoothP_1), .A1 (WindowDin_0__2__0), .S0 (
             Instr)) ;
    mux21_ni L1_0_L2_2_G1_MINI_ALU_ix99 (.Y (L1SecondOperands_2__1), .A0 (
             L1_0_L2_2_G1_MINI_ALU_BoothP_2), .A1 (WindowDin_0__2__1), .S0 (
             Instr)) ;
    mux21_ni L1_0_L2_2_G1_MINI_ALU_ix107 (.Y (L1SecondOperands_2__2), .A0 (
             L1_0_L2_2_G1_MINI_ALU_BoothP_3), .A1 (WindowDin_0__2__2), .S0 (
             Instr)) ;
    mux21_ni L1_0_L2_2_G1_MINI_ALU_ix115 (.Y (L1SecondOperands_2__3), .A0 (
             L1_0_L2_2_G1_MINI_ALU_BoothP_4), .A1 (WindowDin_0__2__3), .S0 (
             Instr)) ;
    mux21_ni L1_0_L2_2_G1_MINI_ALU_ix123 (.Y (L1SecondOperands_2__4), .A0 (
             L1_0_L2_2_G1_MINI_ALU_BoothP_5), .A1 (WindowDin_0__2__4), .S0 (
             Instr)) ;
    mux21_ni L1_0_L2_2_G1_MINI_ALU_ix131 (.Y (L1SecondOperands_2__5), .A0 (
             L1_0_L2_2_G1_MINI_ALU_BoothP_6), .A1 (WindowDin_0__2__5), .S0 (
             Instr)) ;
    mux21_ni L1_0_L2_2_G1_MINI_ALU_ix139 (.Y (L1SecondOperands_2__6), .A0 (
             L1_0_L2_2_G1_MINI_ALU_BoothP_7), .A1 (WindowDin_0__2__6), .S0 (
             Instr)) ;
    mux21_ni L1_0_L2_2_G1_MINI_ALU_ix147 (.Y (L1SecondOperands_2__7), .A0 (
             L1_0_L2_2_G1_MINI_ALU_BoothP_8), .A1 (WindowDin_0__2__7), .S0 (
             Instr)) ;
    xor2 L1_0_L2_2_G1_MINI_ALU_ix77 (.Y (L1Results_2__1), .A0 (
         L1_0_L2_2_G1_MINI_ALU_nx529), .A1 (L1_0_L2_2_G1_MINI_ALU_nx531)) ;
    nand02 L1_0_L2_2_G1_MINI_ALU_ix530 (.Y (L1_0_L2_2_G1_MINI_ALU_nx529), .A0 (
           L1SecondOperands_2__0), .A1 (L1FirstOperands_2__0)) ;
    xnor2 L1_0_L2_2_G1_MINI_ALU_ix532 (.Y (L1_0_L2_2_G1_MINI_ALU_nx531), .A0 (
          L1SecondOperands_2__1), .A1 (L1FirstOperands_2__1)) ;
    xor2 L1_0_L2_2_G1_MINI_ALU_ix75 (.Y (L1Results_2__2), .A0 (
         L1_0_L2_2_G1_MINI_ALU_nx534), .A1 (L1_0_L2_2_G1_MINI_ALU_nx537)) ;
    aoi32 L1_0_L2_2_G1_MINI_ALU_ix535 (.Y (L1_0_L2_2_G1_MINI_ALU_nx534), .A0 (
          L1SecondOperands_2__0), .A1 (L1FirstOperands_2__0), .A2 (
          L1_0_L2_2_G1_MINI_ALU_nx30), .B0 (L1FirstOperands_2__1), .B1 (
          L1SecondOperands_2__1)) ;
    xnor2 L1_0_L2_2_G1_MINI_ALU_ix538 (.Y (L1_0_L2_2_G1_MINI_ALU_nx537), .A0 (
          L1SecondOperands_2__2), .A1 (L1FirstOperands_2__2)) ;
    xor2 L1_0_L2_2_G1_MINI_ALU_ix73 (.Y (L1Results_2__3), .A0 (
         L1_0_L2_2_G1_MINI_ALU_nx540), .A1 (L1_0_L2_2_G1_MINI_ALU_nx544)) ;
    aoi22 L1_0_L2_2_G1_MINI_ALU_ix541 (.Y (L1_0_L2_2_G1_MINI_ALU_nx540), .A0 (
          L1FirstOperands_2__2), .A1 (L1SecondOperands_2__2), .B0 (
          L1_0_L2_2_G1_MINI_ALU_nx40), .B1 (L1_0_L2_2_G1_MINI_ALU_nx24)) ;
    xnor2 L1_0_L2_2_G1_MINI_ALU_ix545 (.Y (L1_0_L2_2_G1_MINI_ALU_nx544), .A0 (
          L1SecondOperands_2__3), .A1 (L1FirstOperands_2__3)) ;
    xor2 L1_0_L2_2_G1_MINI_ALU_ix71 (.Y (L1Results_2__4), .A0 (
         L1_0_L2_2_G1_MINI_ALU_nx547), .A1 (L1_0_L2_2_G1_MINI_ALU_nx551)) ;
    aoi22 L1_0_L2_2_G1_MINI_ALU_ix548 (.Y (L1_0_L2_2_G1_MINI_ALU_nx547), .A0 (
          L1FirstOperands_2__3), .A1 (L1SecondOperands_2__3), .B0 (
          L1_0_L2_2_G1_MINI_ALU_nx44), .B1 (L1_0_L2_2_G1_MINI_ALU_nx18)) ;
    xnor2 L1_0_L2_2_G1_MINI_ALU_ix552 (.Y (L1_0_L2_2_G1_MINI_ALU_nx551), .A0 (
          L1SecondOperands_2__4), .A1 (L1FirstOperands_2__4)) ;
    xor2 L1_0_L2_2_G1_MINI_ALU_ix69 (.Y (L1Results_2__5), .A0 (
         L1_0_L2_2_G1_MINI_ALU_nx554), .A1 (L1_0_L2_2_G1_MINI_ALU_nx558)) ;
    aoi22 L1_0_L2_2_G1_MINI_ALU_ix555 (.Y (L1_0_L2_2_G1_MINI_ALU_nx554), .A0 (
          L1FirstOperands_2__4), .A1 (L1SecondOperands_2__4), .B0 (
          L1_0_L2_2_G1_MINI_ALU_nx48), .B1 (L1_0_L2_2_G1_MINI_ALU_nx12)) ;
    xnor2 L1_0_L2_2_G1_MINI_ALU_ix559 (.Y (L1_0_L2_2_G1_MINI_ALU_nx558), .A0 (
          L1SecondOperands_2__5), .A1 (L1FirstOperands_2__5)) ;
    xor2 L1_0_L2_2_G1_MINI_ALU_ix67 (.Y (L1Results_2__6), .A0 (
         L1_0_L2_2_G1_MINI_ALU_nx561), .A1 (L1_0_L2_2_G1_MINI_ALU_nx565)) ;
    aoi22 L1_0_L2_2_G1_MINI_ALU_ix562 (.Y (L1_0_L2_2_G1_MINI_ALU_nx561), .A0 (
          L1FirstOperands_2__5), .A1 (L1SecondOperands_2__5), .B0 (
          L1_0_L2_2_G1_MINI_ALU_nx52), .B1 (L1_0_L2_2_G1_MINI_ALU_nx6)) ;
    xnor2 L1_0_L2_2_G1_MINI_ALU_ix566 (.Y (L1_0_L2_2_G1_MINI_ALU_nx565), .A0 (
          L1SecondOperands_2__6), .A1 (L1FirstOperands_2__6)) ;
    xnor2 L1_0_L2_2_G1_MINI_ALU_ix65 (.Y (L1Results_2__7), .A0 (
          L1_0_L2_2_G1_MINI_ALU_nx568), .A1 (L1_0_L2_2_G1_MINI_ALU_nx62)) ;
    aoi22 L1_0_L2_2_G1_MINI_ALU_ix569 (.Y (L1_0_L2_2_G1_MINI_ALU_nx568), .A0 (
          L1FirstOperands_2__6), .A1 (L1SecondOperands_2__6), .B0 (
          L1_0_L2_2_G1_MINI_ALU_nx56), .B1 (L1_0_L2_2_G1_MINI_ALU_nx0)) ;
    xor2 L1_0_L2_2_G1_MINI_ALU_ix63 (.Y (L1_0_L2_2_G1_MINI_ALU_nx62), .A0 (
         L1SecondOperands_2__7), .A1 (L1FirstOperands_2__7)) ;
    inv01 L1_0_L2_2_G1_MINI_ALU_ix155 (.Y (L1_0_L2_2_G1_MINI_ALU_nx154), .A (
          L1_0_L2_2_G1_MINI_ALU_nx383)) ;
    inv01 L1_0_L2_2_G1_MINI_ALU_ix57 (.Y (L1_0_L2_2_G1_MINI_ALU_nx56), .A (
          L1_0_L2_2_G1_MINI_ALU_nx561)) ;
    inv01 L1_0_L2_2_G1_MINI_ALU_ix53 (.Y (L1_0_L2_2_G1_MINI_ALU_nx52), .A (
          L1_0_L2_2_G1_MINI_ALU_nx554)) ;
    inv01 L1_0_L2_2_G1_MINI_ALU_ix49 (.Y (L1_0_L2_2_G1_MINI_ALU_nx48), .A (
          L1_0_L2_2_G1_MINI_ALU_nx547)) ;
    inv01 L1_0_L2_2_G1_MINI_ALU_ix45 (.Y (L1_0_L2_2_G1_MINI_ALU_nx44), .A (
          L1_0_L2_2_G1_MINI_ALU_nx540)) ;
    inv01 L1_0_L2_2_G1_MINI_ALU_ix41 (.Y (L1_0_L2_2_G1_MINI_ALU_nx40), .A (
          L1_0_L2_2_G1_MINI_ALU_nx534)) ;
    inv01 L1_0_L2_2_G1_MINI_ALU_ix31 (.Y (L1_0_L2_2_G1_MINI_ALU_nx30), .A (
          L1_0_L2_2_G1_MINI_ALU_nx531)) ;
    inv01 L1_0_L2_2_G1_MINI_ALU_ix25 (.Y (L1_0_L2_2_G1_MINI_ALU_nx24), .A (
          L1_0_L2_2_G1_MINI_ALU_nx537)) ;
    inv01 L1_0_L2_2_G1_MINI_ALU_ix19 (.Y (L1_0_L2_2_G1_MINI_ALU_nx18), .A (
          L1_0_L2_2_G1_MINI_ALU_nx544)) ;
    inv01 L1_0_L2_2_G1_MINI_ALU_ix13 (.Y (L1_0_L2_2_G1_MINI_ALU_nx12), .A (
          L1_0_L2_2_G1_MINI_ALU_nx551)) ;
    inv01 L1_0_L2_2_G1_MINI_ALU_ix7 (.Y (L1_0_L2_2_G1_MINI_ALU_nx6), .A (
          L1_0_L2_2_G1_MINI_ALU_nx558)) ;
    inv01 L1_0_L2_2_G1_MINI_ALU_ix1 (.Y (L1_0_L2_2_G1_MINI_ALU_nx0), .A (
          L1_0_L2_2_G1_MINI_ALU_nx565)) ;
    fake_gnd L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix216 (.Y (
             L1_0_L2_2_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    nor02ii L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix81 (.Y (
            L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx80), .A0 (Instr), .A1 (Start)) ;
    aoi21 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix77 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_10), .A0 (
          FilterDin_0__2__1), .A1 (FilterDin_0__2__0), .B0 (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx4)) ;
    nor02_2x L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix5 (.Y (
             L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx4), .A0 (FilterDin_0__2__0), .A1 (
             FilterDin_0__2__1)) ;
    aoi21 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix67 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_11), .A0 (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx328), .A1 (FilterDin_0__2__2), .B0 (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx8)) ;
    nor03_2x L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix9 (.Y (
             L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx8), .A0 (FilterDin_0__2__2), .A1 (
             FilterDin_0__2__0), .A2 (FilterDin_0__2__1)) ;
    xnor2 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix59 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_12), .A0 (
          FilterDin_0__2__3), .A1 (L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx8)) ;
    xnor2 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix51 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_13), .A0 (
          FilterDin_0__2__4), .A1 (L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx12)) ;
    nor04 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix13 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx12), .A0 (FilterDin_0__2__3), .A1 (
          FilterDin_0__2__2), .A2 (FilterDin_0__2__0), .A3 (FilterDin_0__2__1)
          ) ;
    xnor2 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix43 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_14), .A0 (
          FilterDin_0__2__5), .A1 (L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx16)) ;
    nor02ii L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix17 (.Y (
            L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx16), .A0 (FilterDin_0__2__4), .A1 (
            L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx12)) ;
    xnor2 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix35 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_15), .A0 (
          FilterDin_0__2__6), .A1 (L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx20)) ;
    nor02ii L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix21 (.Y (
            L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx20), .A0 (FilterDin_0__2__5), .A1 (
            L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx16)) ;
    xnor2 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix27 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_16), .A0 (
          FilterDin_0__2__7), .A1 (L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx24)) ;
    nor02ii L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix25 (.Y (
            L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx24), .A0 (FilterDin_0__2__6), .A1 (
            L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx20)) ;
    inv01 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix329 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx328), .A (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx4)) ;
    inv02 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix383 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx384), .A (
          L1_0_L2_2_G1_MINI_ALU_BoothP_0)) ;
    dff L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_0 (.Q (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_0), .QB (\$dummy [106]), 
        .D (L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .CLK (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    nor02_2x L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix567 (.Y (
             L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566), .A0 (RST), .A1 (
             L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644)) ;
    dff L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_1 (.Q (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_1), .QB (\$dummy [107]), 
        .D (L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .CLK (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_2 (.Q (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_2), .QB (\$dummy [108]), 
        .D (L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .CLK (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_3 (.Q (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_3), .QB (\$dummy [109]), 
        .D (L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .CLK (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_4 (.Q (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_4), .QB (\$dummy [110]), 
        .D (L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .CLK (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_5 (.Q (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_5), .QB (\$dummy [111]), 
        .D (L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .CLK (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_6 (.Q (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_6), .QB (\$dummy [112]), 
        .D (L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .CLK (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_7 (.Q (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_7), .QB (\$dummy [113]), 
        .D (L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .CLK (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_8 (.Q (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_8), .QB (\$dummy [114]), 
        .D (L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .CLK (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_9 (.Q (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_9), .QB (\$dummy [115]), 
        .D (L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .CLK (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_10 (.Q (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_10), .QB (\$dummy [116])
        , .D (L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .CLK (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_11 (.Q (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_11), .QB (\$dummy [117])
        , .D (L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .CLK (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_12 (.Q (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_12), .QB (\$dummy [118])
        , .D (L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .CLK (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_13 (.Q (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_13), .QB (\$dummy [119])
        , .D (L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .CLK (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_14 (.Q (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_14), .QB (\$dummy [120])
        , .D (L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .CLK (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_15 (.Q (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_15), .QB (\$dummy [121])
        , .D (L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .CLK (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_16 (.Q (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_16), .QB (\$dummy [122])
        , .D (L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .CLK (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    inv02 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix623 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624), .A (CLK)) ;
    inv02 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix625 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626), .A (CLK)) ;
    inv02 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix627 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628), .A (CLK)) ;
    inv02 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix643 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644), .A (nx7698)) ;
    dff L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_0 (.Q (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_0), .QB (\$dummy [123]), 
        .D (L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .CLK (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    nor02_2x L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix567 (.Y (
             L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566), .A0 (RST), .A1 (
             L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644)) ;
    dff L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_1 (.Q (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_1), .QB (\$dummy [124]), 
        .D (L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .CLK (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_2 (.Q (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_2), .QB (\$dummy [125]), 
        .D (L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .CLK (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_3 (.Q (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_3), .QB (\$dummy [126]), 
        .D (L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .CLK (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_4 (.Q (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_4), .QB (\$dummy [127]), 
        .D (L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .CLK (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_5 (.Q (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_5), .QB (\$dummy [128]), 
        .D (L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .CLK (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_6 (.Q (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_6), .QB (\$dummy [129]), 
        .D (L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .CLK (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_7 (.Q (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_7), .QB (\$dummy [130]), 
        .D (L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .CLK (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_8 (.Q (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_8), .QB (\$dummy [131]), 
        .D (L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .CLK (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_9 (.Q (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_9), .QB (\$dummy [132]), 
        .D (L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .CLK (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_10 (.Q (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_10), .QB (\$dummy [133])
        , .D (L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .CLK (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_11 (.Q (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_11), .QB (\$dummy [134])
        , .D (L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .CLK (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_12 (.Q (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_12), .QB (\$dummy [135])
        , .D (L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .CLK (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_13 (.Q (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_13), .QB (\$dummy [136])
        , .D (L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .CLK (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_14 (.Q (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_14), .QB (\$dummy [137])
        , .D (L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .CLK (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_15 (.Q (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_15), .QB (\$dummy [138])
        , .D (L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .CLK (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_16 (.Q (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_16), .QB (\$dummy [139])
        , .D (L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .CLK (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    inv02 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix623 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624), .A (CLK)) ;
    inv02 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix625 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626), .A (CLK)) ;
    inv02 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix627 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628), .A (CLK)) ;
    inv02 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix643 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644), .A (nx7704)) ;
    dff L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_0 (.Q (
        L1_0_L2_2_G1_MINI_ALU_BoothP_0), .QB (\$dummy [140]), .D (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .CLK (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    nor02_2x L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix567 (.Y (
             L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566), .A0 (RST), .A1 (
             L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    dff L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_1 (.Q (
        L1_0_L2_2_G1_MINI_ALU_BoothP_1), .QB (\$dummy [141]), .D (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .CLK (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_2 (.Q (
        L1_0_L2_2_G1_MINI_ALU_BoothP_2), .QB (\$dummy [142]), .D (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .CLK (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_3 (.Q (
        L1_0_L2_2_G1_MINI_ALU_BoothP_3), .QB (\$dummy [143]), .D (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .CLK (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_4 (.Q (
        L1_0_L2_2_G1_MINI_ALU_BoothP_4), .QB (\$dummy [144]), .D (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .CLK (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_5 (.Q (
        L1_0_L2_2_G1_MINI_ALU_BoothP_5), .QB (\$dummy [145]), .D (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .CLK (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_6 (.Q (
        L1_0_L2_2_G1_MINI_ALU_BoothP_6), .QB (\$dummy [146]), .D (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .CLK (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_7 (.Q (
        L1_0_L2_2_G1_MINI_ALU_BoothP_7), .QB (\$dummy [147]), .D (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .CLK (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_8 (.Q (
        L1_0_L2_2_G1_MINI_ALU_BoothP_8), .QB (\$dummy [148]), .D (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .CLK (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_9 (.Q (
        L1_0_L2_2_G1_MINI_ALU_BoothP_9), .QB (\$dummy [149]), .D (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .CLK (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_10 (.Q (
        L1_0_L2_2_G1_MINI_ALU_BoothP_10), .QB (\$dummy [150]), .D (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .CLK (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_11 (.Q (
        L1_0_L2_2_G1_MINI_ALU_BoothP_11), .QB (\$dummy [151]), .D (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .CLK (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_12 (.Q (
        L1_0_L2_2_G1_MINI_ALU_BoothP_12), .QB (\$dummy [152]), .D (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .CLK (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_13 (.Q (
        L1_0_L2_2_G1_MINI_ALU_BoothP_13), .QB (\$dummy [153]), .D (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .CLK (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_14 (.Q (
        L1_0_L2_2_G1_MINI_ALU_BoothP_14), .QB (\$dummy [154]), .D (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .CLK (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_15 (.Q (
        L1_0_L2_2_G1_MINI_ALU_BoothP_15), .QB (\$dummy [155]), .D (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .CLK (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_16 (.Q (
        L1_0_L2_2_G1_MINI_ALU_BoothP_16), .QB (\$dummy [156]), .D (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .CLK (
        L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    inv02 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix623 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624), .A (CLK)) ;
    inv02 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix625 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626), .A (CLK)) ;
    inv02 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix627 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628), .A (CLK)) ;
    inv02 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix643 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644), .A (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642)) ;
    xor2 L1_0_L2_3_G1_MINI_ALU_ix83 (.Y (L1Results_3__0), .A0 (
         L1SecondOperands_3__0), .A1 (L1FirstOperands_3__0)) ;
    xnor2 L1_0_L2_3_G1_MINI_ALU_ix380 (.Y (L1_0_L2_3_G1_MINI_ALU_nx379), .A0 (
          L1_0_L2_3_G1_MINI_ALU_nx381), .A1 (L1_0_L2_3_G1_MINI_ALU_nx383)) ;
    nand02 L1_0_L2_3_G1_MINI_ALU_ix382 (.Y (L1_0_L2_3_G1_MINI_ALU_nx381), .A0 (
           L1_0_L2_3_G1_MINI_ALU_BoothOperand_0), .A1 (nx7724)) ;
    xnor2 L1_0_L2_3_G1_MINI_ALU_ix384 (.Y (L1_0_L2_3_G1_MINI_ALU_nx383), .A0 (
          L1_0_L2_3_G1_MINI_ALU_BoothOperand_1), .A1 (
          L1_0_L2_3_G1_MINI_ALU_BoothP_1)) ;
    inv01 L1_0_L2_3_G1_MINI_ALU_ix388 (.Y (L1_0_L2_3_G1_MINI_ALU_nx387), .A (
          L1_0_L2_3_G1_MINI_ALU_BoothP_2)) ;
    xnor2 L1_0_L2_3_G1_MINI_ALU_ix390 (.Y (L1_0_L2_3_G1_MINI_ALU_nx389), .A0 (
          L1_0_L2_3_G1_MINI_ALU_nx391), .A1 (L1_0_L2_3_G1_MINI_ALU_nx395)) ;
    aoi32 L1_0_L2_3_G1_MINI_ALU_ix392 (.Y (L1_0_L2_3_G1_MINI_ALU_nx391), .A0 (
          L1_0_L2_3_G1_MINI_ALU_BoothOperand_0), .A1 (nx7724), .A2 (
          L1_0_L2_3_G1_MINI_ALU_nx154), .B0 (L1_0_L2_3_G1_MINI_ALU_BoothP_1), .B1 (
          L1_0_L2_3_G1_MINI_ALU_BoothOperand_1)) ;
    xnor2 L1_0_L2_3_G1_MINI_ALU_ix396 (.Y (L1_0_L2_3_G1_MINI_ALU_nx395), .A0 (
          L1_0_L2_3_G1_MINI_ALU_BoothOperand_2), .A1 (
          L1_0_L2_3_G1_MINI_ALU_BoothP_2)) ;
    inv01 L1_0_L2_3_G1_MINI_ALU_ix400 (.Y (L1_0_L2_3_G1_MINI_ALU_nx399), .A (
          L1_0_L2_3_G1_MINI_ALU_BoothP_3)) ;
    xnor2 L1_0_L2_3_G1_MINI_ALU_ix402 (.Y (L1_0_L2_3_G1_MINI_ALU_nx401), .A0 (
          L1_0_L2_3_G1_MINI_ALU_nx403), .A1 (L1_0_L2_3_G1_MINI_ALU_nx405)) ;
    xnor2 L1_0_L2_3_G1_MINI_ALU_ix406 (.Y (L1_0_L2_3_G1_MINI_ALU_nx405), .A0 (
          L1_0_L2_3_G1_MINI_ALU_BoothOperand_3), .A1 (
          L1_0_L2_3_G1_MINI_ALU_BoothP_3)) ;
    inv01 L1_0_L2_3_G1_MINI_ALU_ix410 (.Y (L1_0_L2_3_G1_MINI_ALU_nx409), .A (
          L1_0_L2_3_G1_MINI_ALU_BoothP_4)) ;
    xnor2 L1_0_L2_3_G1_MINI_ALU_ix412 (.Y (L1_0_L2_3_G1_MINI_ALU_nx411), .A0 (
          L1_0_L2_3_G1_MINI_ALU_nx413), .A1 (L1_0_L2_3_G1_MINI_ALU_nx415)) ;
    xnor2 L1_0_L2_3_G1_MINI_ALU_ix416 (.Y (L1_0_L2_3_G1_MINI_ALU_nx415), .A0 (
          L1_0_L2_3_G1_MINI_ALU_BoothOperand_4), .A1 (
          L1_0_L2_3_G1_MINI_ALU_BoothP_4)) ;
    inv01 L1_0_L2_3_G1_MINI_ALU_ix420 (.Y (L1_0_L2_3_G1_MINI_ALU_nx419), .A (
          L1_0_L2_3_G1_MINI_ALU_BoothP_5)) ;
    xnor2 L1_0_L2_3_G1_MINI_ALU_ix422 (.Y (L1_0_L2_3_G1_MINI_ALU_nx421), .A0 (
          L1_0_L2_3_G1_MINI_ALU_nx423), .A1 (L1_0_L2_3_G1_MINI_ALU_nx425)) ;
    xnor2 L1_0_L2_3_G1_MINI_ALU_ix426 (.Y (L1_0_L2_3_G1_MINI_ALU_nx425), .A0 (
          L1_0_L2_3_G1_MINI_ALU_BoothOperand_5), .A1 (
          L1_0_L2_3_G1_MINI_ALU_BoothP_5)) ;
    inv01 L1_0_L2_3_G1_MINI_ALU_ix430 (.Y (L1_0_L2_3_G1_MINI_ALU_nx429), .A (
          L1_0_L2_3_G1_MINI_ALU_BoothP_6)) ;
    xnor2 L1_0_L2_3_G1_MINI_ALU_ix432 (.Y (L1_0_L2_3_G1_MINI_ALU_nx431), .A0 (
          L1_0_L2_3_G1_MINI_ALU_nx433), .A1 (L1_0_L2_3_G1_MINI_ALU_nx435)) ;
    xnor2 L1_0_L2_3_G1_MINI_ALU_ix436 (.Y (L1_0_L2_3_G1_MINI_ALU_nx435), .A0 (
          L1_0_L2_3_G1_MINI_ALU_BoothOperand_6), .A1 (
          L1_0_L2_3_G1_MINI_ALU_BoothP_6)) ;
    inv01 L1_0_L2_3_G1_MINI_ALU_ix440 (.Y (L1_0_L2_3_G1_MINI_ALU_nx439), .A (
          L1_0_L2_3_G1_MINI_ALU_BoothP_7)) ;
    xnor2 L1_0_L2_3_G1_MINI_ALU_ix442 (.Y (L1_0_L2_3_G1_MINI_ALU_nx441), .A0 (
          L1_0_L2_3_G1_MINI_ALU_nx443), .A1 (L1_0_L2_3_G1_MINI_ALU_nx445)) ;
    xnor2 L1_0_L2_3_G1_MINI_ALU_ix446 (.Y (L1_0_L2_3_G1_MINI_ALU_nx445), .A0 (
          L1_0_L2_3_G1_MINI_ALU_BoothOperand_7), .A1 (
          L1_0_L2_3_G1_MINI_ALU_BoothP_7)) ;
    inv01 L1_0_L2_3_G1_MINI_ALU_ix450 (.Y (L1_0_L2_3_G1_MINI_ALU_nx449), .A (
          L1_0_L2_3_G1_MINI_ALU_BoothP_8)) ;
    xnor2 L1_0_L2_3_G1_MINI_ALU_ix452 (.Y (L1_0_L2_3_G1_MINI_ALU_nx451), .A0 (
          L1_0_L2_3_G1_MINI_ALU_nx453), .A1 (L1_0_L2_3_G1_MINI_ALU_nx455)) ;
    xnor2 L1_0_L2_3_G1_MINI_ALU_ix456 (.Y (L1_0_L2_3_G1_MINI_ALU_nx455), .A0 (
          L1_0_L2_3_G1_MINI_ALU_BoothOperand_8), .A1 (
          L1_0_L2_3_G1_MINI_ALU_BoothP_8)) ;
    xor2 L1_0_L2_3_G1_MINI_ALU_ix317 (.Y (L1_0_L2_3_G1_MINI_ALU_nx316), .A0 (
         L1_0_L2_3_G1_MINI_ALU_nx461), .A1 (L1_0_L2_3_G1_MINI_ALU_nx463)) ;
    xnor2 L1_0_L2_3_G1_MINI_ALU_ix464 (.Y (L1_0_L2_3_G1_MINI_ALU_nx463), .A0 (
          L1_0_L2_3_G1_MINI_ALU_BoothOperand_9), .A1 (
          L1_0_L2_3_G1_MINI_ALU_BoothP_9)) ;
    xor2 L1_0_L2_3_G1_MINI_ALU_ix337 (.Y (L1_0_L2_3_G1_MINI_ALU_nx336), .A0 (
         L1_0_L2_3_G1_MINI_ALU_nx467), .A1 (L1_0_L2_3_G1_MINI_ALU_nx471)) ;
    inv01 L1_0_L2_3_G1_MINI_ALU_ix470 (.Y (L1_0_L2_3_G1_MINI_ALU_nx469), .A (
          L1_0_L2_3_G1_MINI_ALU_BoothP_9)) ;
    xnor2 L1_0_L2_3_G1_MINI_ALU_ix472 (.Y (L1_0_L2_3_G1_MINI_ALU_nx471), .A0 (
          L1_0_L2_3_G1_MINI_ALU_BoothOperand_10), .A1 (
          L1_0_L2_3_G1_MINI_ALU_BoothP_10)) ;
    xor2 L1_0_L2_3_G1_MINI_ALU_ix357 (.Y (L1_0_L2_3_G1_MINI_ALU_nx356), .A0 (
         L1_0_L2_3_G1_MINI_ALU_nx475), .A1 (L1_0_L2_3_G1_MINI_ALU_nx479)) ;
    inv01 L1_0_L2_3_G1_MINI_ALU_ix478 (.Y (L1_0_L2_3_G1_MINI_ALU_nx477), .A (
          L1_0_L2_3_G1_MINI_ALU_BoothP_10)) ;
    xnor2 L1_0_L2_3_G1_MINI_ALU_ix480 (.Y (L1_0_L2_3_G1_MINI_ALU_nx479), .A0 (
          L1_0_L2_3_G1_MINI_ALU_BoothOperand_11), .A1 (
          L1_0_L2_3_G1_MINI_ALU_BoothP_11)) ;
    xor2 L1_0_L2_3_G1_MINI_ALU_ix377 (.Y (L1_0_L2_3_G1_MINI_ALU_nx376), .A0 (
         L1_0_L2_3_G1_MINI_ALU_nx483), .A1 (L1_0_L2_3_G1_MINI_ALU_nx487)) ;
    inv01 L1_0_L2_3_G1_MINI_ALU_ix486 (.Y (L1_0_L2_3_G1_MINI_ALU_nx485), .A (
          L1_0_L2_3_G1_MINI_ALU_BoothP_11)) ;
    xnor2 L1_0_L2_3_G1_MINI_ALU_ix488 (.Y (L1_0_L2_3_G1_MINI_ALU_nx487), .A0 (
          L1_0_L2_3_G1_MINI_ALU_BoothOperand_12), .A1 (
          L1_0_L2_3_G1_MINI_ALU_BoothP_12)) ;
    xor2 L1_0_L2_3_G1_MINI_ALU_ix397 (.Y (L1_0_L2_3_G1_MINI_ALU_nx396), .A0 (
         L1_0_L2_3_G1_MINI_ALU_nx491), .A1 (L1_0_L2_3_G1_MINI_ALU_nx495)) ;
    inv01 L1_0_L2_3_G1_MINI_ALU_ix494 (.Y (L1_0_L2_3_G1_MINI_ALU_nx493), .A (
          L1_0_L2_3_G1_MINI_ALU_BoothP_12)) ;
    xnor2 L1_0_L2_3_G1_MINI_ALU_ix496 (.Y (L1_0_L2_3_G1_MINI_ALU_nx495), .A0 (
          L1_0_L2_3_G1_MINI_ALU_BoothOperand_13), .A1 (
          L1_0_L2_3_G1_MINI_ALU_BoothP_13)) ;
    xor2 L1_0_L2_3_G1_MINI_ALU_ix417 (.Y (L1_0_L2_3_G1_MINI_ALU_nx416), .A0 (
         L1_0_L2_3_G1_MINI_ALU_nx499), .A1 (L1_0_L2_3_G1_MINI_ALU_nx503)) ;
    inv01 L1_0_L2_3_G1_MINI_ALU_ix502 (.Y (L1_0_L2_3_G1_MINI_ALU_nx501), .A (
          L1_0_L2_3_G1_MINI_ALU_BoothP_13)) ;
    xnor2 L1_0_L2_3_G1_MINI_ALU_ix504 (.Y (L1_0_L2_3_G1_MINI_ALU_nx503), .A0 (
          L1_0_L2_3_G1_MINI_ALU_BoothOperand_14), .A1 (
          L1_0_L2_3_G1_MINI_ALU_BoothP_14)) ;
    xor2 L1_0_L2_3_G1_MINI_ALU_ix437 (.Y (L1_0_L2_3_G1_MINI_ALU_nx436), .A0 (
         L1_0_L2_3_G1_MINI_ALU_nx507), .A1 (L1_0_L2_3_G1_MINI_ALU_nx511)) ;
    inv01 L1_0_L2_3_G1_MINI_ALU_ix510 (.Y (L1_0_L2_3_G1_MINI_ALU_nx509), .A (
          L1_0_L2_3_G1_MINI_ALU_BoothP_14)) ;
    xnor2 L1_0_L2_3_G1_MINI_ALU_ix512 (.Y (L1_0_L2_3_G1_MINI_ALU_nx511), .A0 (
          L1_0_L2_3_G1_MINI_ALU_BoothOperand_15), .A1 (
          L1_0_L2_3_G1_MINI_ALU_BoothP_15)) ;
    xnor2 L1_0_L2_3_G1_MINI_ALU_ix457 (.Y (L1_0_L2_3_G1_MINI_ALU_nx456), .A0 (
          L1_0_L2_3_G1_MINI_ALU_nx515), .A1 (L1_0_L2_3_G1_MINI_ALU_nx454)) ;
    inv01 L1_0_L2_3_G1_MINI_ALU_ix518 (.Y (L1_0_L2_3_G1_MINI_ALU_nx517), .A (
          L1_0_L2_3_G1_MINI_ALU_BoothP_15)) ;
    xor2 L1_0_L2_3_G1_MINI_ALU_ix455 (.Y (L1_0_L2_3_G1_MINI_ALU_nx454), .A0 (
         L1_0_L2_3_G1_MINI_ALU_BoothOperand_16), .A1 (
         L1_0_L2_3_G1_MINI_ALU_BoothP_16)) ;
    mux21_ni L1_0_L2_3_G1_MINI_ALU_ix91 (.Y (L1SecondOperands_3__0), .A0 (
             L1_0_L2_3_G1_MINI_ALU_BoothP_1), .A1 (WindowDin_0__3__0), .S0 (
             Instr)) ;
    mux21_ni L1_0_L2_3_G1_MINI_ALU_ix99 (.Y (L1SecondOperands_3__1), .A0 (
             L1_0_L2_3_G1_MINI_ALU_BoothP_2), .A1 (WindowDin_0__3__1), .S0 (
             Instr)) ;
    mux21_ni L1_0_L2_3_G1_MINI_ALU_ix107 (.Y (L1SecondOperands_3__2), .A0 (
             L1_0_L2_3_G1_MINI_ALU_BoothP_3), .A1 (WindowDin_0__3__2), .S0 (
             Instr)) ;
    mux21_ni L1_0_L2_3_G1_MINI_ALU_ix115 (.Y (L1SecondOperands_3__3), .A0 (
             L1_0_L2_3_G1_MINI_ALU_BoothP_4), .A1 (WindowDin_0__3__3), .S0 (
             Instr)) ;
    mux21_ni L1_0_L2_3_G1_MINI_ALU_ix123 (.Y (L1SecondOperands_3__4), .A0 (
             L1_0_L2_3_G1_MINI_ALU_BoothP_5), .A1 (WindowDin_0__3__4), .S0 (
             Instr)) ;
    mux21_ni L1_0_L2_3_G1_MINI_ALU_ix131 (.Y (L1SecondOperands_3__5), .A0 (
             L1_0_L2_3_G1_MINI_ALU_BoothP_6), .A1 (WindowDin_0__3__5), .S0 (
             Instr)) ;
    mux21_ni L1_0_L2_3_G1_MINI_ALU_ix139 (.Y (L1SecondOperands_3__6), .A0 (
             L1_0_L2_3_G1_MINI_ALU_BoothP_7), .A1 (WindowDin_0__3__6), .S0 (
             Instr)) ;
    mux21_ni L1_0_L2_3_G1_MINI_ALU_ix147 (.Y (L1SecondOperands_3__7), .A0 (
             L1_0_L2_3_G1_MINI_ALU_BoothP_8), .A1 (WindowDin_0__3__7), .S0 (
             Instr)) ;
    xor2 L1_0_L2_3_G1_MINI_ALU_ix77 (.Y (L1Results_3__1), .A0 (
         L1_0_L2_3_G1_MINI_ALU_nx529), .A1 (L1_0_L2_3_G1_MINI_ALU_nx531)) ;
    nand02 L1_0_L2_3_G1_MINI_ALU_ix530 (.Y (L1_0_L2_3_G1_MINI_ALU_nx529), .A0 (
           L1SecondOperands_3__0), .A1 (L1FirstOperands_3__0)) ;
    xnor2 L1_0_L2_3_G1_MINI_ALU_ix532 (.Y (L1_0_L2_3_G1_MINI_ALU_nx531), .A0 (
          L1SecondOperands_3__1), .A1 (L1FirstOperands_3__1)) ;
    xor2 L1_0_L2_3_G1_MINI_ALU_ix75 (.Y (L1Results_3__2), .A0 (
         L1_0_L2_3_G1_MINI_ALU_nx534), .A1 (L1_0_L2_3_G1_MINI_ALU_nx537)) ;
    aoi32 L1_0_L2_3_G1_MINI_ALU_ix535 (.Y (L1_0_L2_3_G1_MINI_ALU_nx534), .A0 (
          L1SecondOperands_3__0), .A1 (L1FirstOperands_3__0), .A2 (
          L1_0_L2_3_G1_MINI_ALU_nx30), .B0 (L1FirstOperands_3__1), .B1 (
          L1SecondOperands_3__1)) ;
    xnor2 L1_0_L2_3_G1_MINI_ALU_ix538 (.Y (L1_0_L2_3_G1_MINI_ALU_nx537), .A0 (
          L1SecondOperands_3__2), .A1 (L1FirstOperands_3__2)) ;
    xor2 L1_0_L2_3_G1_MINI_ALU_ix73 (.Y (L1Results_3__3), .A0 (
         L1_0_L2_3_G1_MINI_ALU_nx540), .A1 (L1_0_L2_3_G1_MINI_ALU_nx544)) ;
    aoi22 L1_0_L2_3_G1_MINI_ALU_ix541 (.Y (L1_0_L2_3_G1_MINI_ALU_nx540), .A0 (
          L1FirstOperands_3__2), .A1 (L1SecondOperands_3__2), .B0 (
          L1_0_L2_3_G1_MINI_ALU_nx40), .B1 (L1_0_L2_3_G1_MINI_ALU_nx24)) ;
    xnor2 L1_0_L2_3_G1_MINI_ALU_ix545 (.Y (L1_0_L2_3_G1_MINI_ALU_nx544), .A0 (
          L1SecondOperands_3__3), .A1 (L1FirstOperands_3__3)) ;
    xor2 L1_0_L2_3_G1_MINI_ALU_ix71 (.Y (L1Results_3__4), .A0 (
         L1_0_L2_3_G1_MINI_ALU_nx547), .A1 (L1_0_L2_3_G1_MINI_ALU_nx551)) ;
    aoi22 L1_0_L2_3_G1_MINI_ALU_ix548 (.Y (L1_0_L2_3_G1_MINI_ALU_nx547), .A0 (
          L1FirstOperands_3__3), .A1 (L1SecondOperands_3__3), .B0 (
          L1_0_L2_3_G1_MINI_ALU_nx44), .B1 (L1_0_L2_3_G1_MINI_ALU_nx18)) ;
    xnor2 L1_0_L2_3_G1_MINI_ALU_ix552 (.Y (L1_0_L2_3_G1_MINI_ALU_nx551), .A0 (
          L1SecondOperands_3__4), .A1 (L1FirstOperands_3__4)) ;
    xor2 L1_0_L2_3_G1_MINI_ALU_ix69 (.Y (L1Results_3__5), .A0 (
         L1_0_L2_3_G1_MINI_ALU_nx554), .A1 (L1_0_L2_3_G1_MINI_ALU_nx558)) ;
    aoi22 L1_0_L2_3_G1_MINI_ALU_ix555 (.Y (L1_0_L2_3_G1_MINI_ALU_nx554), .A0 (
          L1FirstOperands_3__4), .A1 (L1SecondOperands_3__4), .B0 (
          L1_0_L2_3_G1_MINI_ALU_nx48), .B1 (L1_0_L2_3_G1_MINI_ALU_nx12)) ;
    xnor2 L1_0_L2_3_G1_MINI_ALU_ix559 (.Y (L1_0_L2_3_G1_MINI_ALU_nx558), .A0 (
          L1SecondOperands_3__5), .A1 (L1FirstOperands_3__5)) ;
    xor2 L1_0_L2_3_G1_MINI_ALU_ix67 (.Y (L1Results_3__6), .A0 (
         L1_0_L2_3_G1_MINI_ALU_nx561), .A1 (L1_0_L2_3_G1_MINI_ALU_nx565)) ;
    aoi22 L1_0_L2_3_G1_MINI_ALU_ix562 (.Y (L1_0_L2_3_G1_MINI_ALU_nx561), .A0 (
          L1FirstOperands_3__5), .A1 (L1SecondOperands_3__5), .B0 (
          L1_0_L2_3_G1_MINI_ALU_nx52), .B1 (L1_0_L2_3_G1_MINI_ALU_nx6)) ;
    xnor2 L1_0_L2_3_G1_MINI_ALU_ix566 (.Y (L1_0_L2_3_G1_MINI_ALU_nx565), .A0 (
          L1SecondOperands_3__6), .A1 (L1FirstOperands_3__6)) ;
    xnor2 L1_0_L2_3_G1_MINI_ALU_ix65 (.Y (L1Results_3__7), .A0 (
          L1_0_L2_3_G1_MINI_ALU_nx568), .A1 (L1_0_L2_3_G1_MINI_ALU_nx62)) ;
    aoi22 L1_0_L2_3_G1_MINI_ALU_ix569 (.Y (L1_0_L2_3_G1_MINI_ALU_nx568), .A0 (
          L1FirstOperands_3__6), .A1 (L1SecondOperands_3__6), .B0 (
          L1_0_L2_3_G1_MINI_ALU_nx56), .B1 (L1_0_L2_3_G1_MINI_ALU_nx0)) ;
    xor2 L1_0_L2_3_G1_MINI_ALU_ix63 (.Y (L1_0_L2_3_G1_MINI_ALU_nx62), .A0 (
         L1SecondOperands_3__7), .A1 (L1FirstOperands_3__7)) ;
    inv01 L1_0_L2_3_G1_MINI_ALU_ix155 (.Y (L1_0_L2_3_G1_MINI_ALU_nx154), .A (
          L1_0_L2_3_G1_MINI_ALU_nx383)) ;
    inv01 L1_0_L2_3_G1_MINI_ALU_ix57 (.Y (L1_0_L2_3_G1_MINI_ALU_nx56), .A (
          L1_0_L2_3_G1_MINI_ALU_nx561)) ;
    inv01 L1_0_L2_3_G1_MINI_ALU_ix53 (.Y (L1_0_L2_3_G1_MINI_ALU_nx52), .A (
          L1_0_L2_3_G1_MINI_ALU_nx554)) ;
    inv01 L1_0_L2_3_G1_MINI_ALU_ix49 (.Y (L1_0_L2_3_G1_MINI_ALU_nx48), .A (
          L1_0_L2_3_G1_MINI_ALU_nx547)) ;
    inv01 L1_0_L2_3_G1_MINI_ALU_ix45 (.Y (L1_0_L2_3_G1_MINI_ALU_nx44), .A (
          L1_0_L2_3_G1_MINI_ALU_nx540)) ;
    inv01 L1_0_L2_3_G1_MINI_ALU_ix41 (.Y (L1_0_L2_3_G1_MINI_ALU_nx40), .A (
          L1_0_L2_3_G1_MINI_ALU_nx534)) ;
    inv01 L1_0_L2_3_G1_MINI_ALU_ix31 (.Y (L1_0_L2_3_G1_MINI_ALU_nx30), .A (
          L1_0_L2_3_G1_MINI_ALU_nx531)) ;
    inv01 L1_0_L2_3_G1_MINI_ALU_ix25 (.Y (L1_0_L2_3_G1_MINI_ALU_nx24), .A (
          L1_0_L2_3_G1_MINI_ALU_nx537)) ;
    inv01 L1_0_L2_3_G1_MINI_ALU_ix19 (.Y (L1_0_L2_3_G1_MINI_ALU_nx18), .A (
          L1_0_L2_3_G1_MINI_ALU_nx544)) ;
    inv01 L1_0_L2_3_G1_MINI_ALU_ix13 (.Y (L1_0_L2_3_G1_MINI_ALU_nx12), .A (
          L1_0_L2_3_G1_MINI_ALU_nx551)) ;
    inv01 L1_0_L2_3_G1_MINI_ALU_ix7 (.Y (L1_0_L2_3_G1_MINI_ALU_nx6), .A (
          L1_0_L2_3_G1_MINI_ALU_nx558)) ;
    inv01 L1_0_L2_3_G1_MINI_ALU_ix1 (.Y (L1_0_L2_3_G1_MINI_ALU_nx0), .A (
          L1_0_L2_3_G1_MINI_ALU_nx565)) ;
    fake_gnd L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix216 (.Y (
             L1_0_L2_3_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    nor02ii L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix81 (.Y (
            L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx80), .A0 (Instr), .A1 (Start)) ;
    aoi21 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix77 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_10), .A0 (
          FilterDin_0__3__1), .A1 (FilterDin_0__3__0), .B0 (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx4)) ;
    nor02_2x L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix5 (.Y (
             L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx4), .A0 (FilterDin_0__3__0), .A1 (
             FilterDin_0__3__1)) ;
    aoi21 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix67 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_11), .A0 (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx328), .A1 (FilterDin_0__3__2), .B0 (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx8)) ;
    nor03_2x L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix9 (.Y (
             L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx8), .A0 (FilterDin_0__3__2), .A1 (
             FilterDin_0__3__0), .A2 (FilterDin_0__3__1)) ;
    xnor2 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix59 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_12), .A0 (
          FilterDin_0__3__3), .A1 (L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx8)) ;
    xnor2 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix51 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_13), .A0 (
          FilterDin_0__3__4), .A1 (L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx12)) ;
    nor04 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix13 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx12), .A0 (FilterDin_0__3__3), .A1 (
          FilterDin_0__3__2), .A2 (FilterDin_0__3__0), .A3 (FilterDin_0__3__1)
          ) ;
    xnor2 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix43 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_14), .A0 (
          FilterDin_0__3__5), .A1 (L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx16)) ;
    nor02ii L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix17 (.Y (
            L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx16), .A0 (FilterDin_0__3__4), .A1 (
            L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx12)) ;
    xnor2 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix35 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_15), .A0 (
          FilterDin_0__3__6), .A1 (L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx20)) ;
    nor02ii L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix21 (.Y (
            L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx20), .A0 (FilterDin_0__3__5), .A1 (
            L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx16)) ;
    xnor2 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix27 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_16), .A0 (
          FilterDin_0__3__7), .A1 (L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx24)) ;
    nor02ii L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix25 (.Y (
            L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx24), .A0 (FilterDin_0__3__6), .A1 (
            L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx20)) ;
    inv01 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix329 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx328), .A (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx4)) ;
    inv02 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix383 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx384), .A (
          L1_0_L2_3_G1_MINI_ALU_BoothP_0)) ;
    dff L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_0 (.Q (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_0), .QB (\$dummy [157]), 
        .D (L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .CLK (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    nor02_2x L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix567 (.Y (
             L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566), .A0 (RST), .A1 (
             L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644)) ;
    dff L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_1 (.Q (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_1), .QB (\$dummy [158]), 
        .D (L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .CLK (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_2 (.Q (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_2), .QB (\$dummy [159]), 
        .D (L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .CLK (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_3 (.Q (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_3), .QB (\$dummy [160]), 
        .D (L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .CLK (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_4 (.Q (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_4), .QB (\$dummy [161]), 
        .D (L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .CLK (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_5 (.Q (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_5), .QB (\$dummy [162]), 
        .D (L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .CLK (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_6 (.Q (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_6), .QB (\$dummy [163]), 
        .D (L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .CLK (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_7 (.Q (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_7), .QB (\$dummy [164]), 
        .D (L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .CLK (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_8 (.Q (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_8), .QB (\$dummy [165]), 
        .D (L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .CLK (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_9 (.Q (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_9), .QB (\$dummy [166]), 
        .D (L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .CLK (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_10 (.Q (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_10), .QB (\$dummy [167])
        , .D (L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .CLK (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_11 (.Q (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_11), .QB (\$dummy [168])
        , .D (L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .CLK (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_12 (.Q (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_12), .QB (\$dummy [169])
        , .D (L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .CLK (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_13 (.Q (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_13), .QB (\$dummy [170])
        , .D (L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .CLK (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_14 (.Q (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_14), .QB (\$dummy [171])
        , .D (L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .CLK (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_15 (.Q (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_15), .QB (\$dummy [172])
        , .D (L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .CLK (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_16 (.Q (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_16), .QB (\$dummy [173])
        , .D (L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .CLK (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    inv02 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix623 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624), .A (CLK)) ;
    inv02 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix625 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626), .A (CLK)) ;
    inv02 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix627 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628), .A (CLK)) ;
    inv02 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix643 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644), .A (nx7738)) ;
    dff L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_0 (.Q (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_0), .QB (\$dummy [174]), 
        .D (L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .CLK (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    nor02_2x L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix567 (.Y (
             L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566), .A0 (RST), .A1 (
             L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644)) ;
    dff L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_1 (.Q (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_1), .QB (\$dummy [175]), 
        .D (L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .CLK (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_2 (.Q (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_2), .QB (\$dummy [176]), 
        .D (L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .CLK (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_3 (.Q (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_3), .QB (\$dummy [177]), 
        .D (L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .CLK (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_4 (.Q (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_4), .QB (\$dummy [178]), 
        .D (L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .CLK (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_5 (.Q (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_5), .QB (\$dummy [179]), 
        .D (L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .CLK (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_6 (.Q (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_6), .QB (\$dummy [180]), 
        .D (L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .CLK (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_7 (.Q (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_7), .QB (\$dummy [181]), 
        .D (L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .CLK (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_8 (.Q (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_8), .QB (\$dummy [182]), 
        .D (L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .CLK (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_9 (.Q (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_9), .QB (\$dummy [183]), 
        .D (L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .CLK (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_10 (.Q (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_10), .QB (\$dummy [184])
        , .D (L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .CLK (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_11 (.Q (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_11), .QB (\$dummy [185])
        , .D (L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .CLK (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_12 (.Q (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_12), .QB (\$dummy [186])
        , .D (L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .CLK (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_13 (.Q (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_13), .QB (\$dummy [187])
        , .D (L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .CLK (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_14 (.Q (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_14), .QB (\$dummy [188])
        , .D (L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .CLK (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_15 (.Q (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_15), .QB (\$dummy [189])
        , .D (L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .CLK (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_16 (.Q (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_16), .QB (\$dummy [190])
        , .D (L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .CLK (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    inv02 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix623 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624), .A (CLK)) ;
    inv02 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix625 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626), .A (CLK)) ;
    inv02 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix627 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628), .A (CLK)) ;
    inv02 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix643 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644), .A (nx7744)) ;
    dff L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_0 (.Q (
        L1_0_L2_3_G1_MINI_ALU_BoothP_0), .QB (\$dummy [191]), .D (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .CLK (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    nor02_2x L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix567 (.Y (
             L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566), .A0 (RST), .A1 (
             L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    dff L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_1 (.Q (
        L1_0_L2_3_G1_MINI_ALU_BoothP_1), .QB (\$dummy [192]), .D (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .CLK (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_2 (.Q (
        L1_0_L2_3_G1_MINI_ALU_BoothP_2), .QB (\$dummy [193]), .D (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .CLK (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_3 (.Q (
        L1_0_L2_3_G1_MINI_ALU_BoothP_3), .QB (\$dummy [194]), .D (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .CLK (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_4 (.Q (
        L1_0_L2_3_G1_MINI_ALU_BoothP_4), .QB (\$dummy [195]), .D (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .CLK (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_5 (.Q (
        L1_0_L2_3_G1_MINI_ALU_BoothP_5), .QB (\$dummy [196]), .D (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .CLK (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_6 (.Q (
        L1_0_L2_3_G1_MINI_ALU_BoothP_6), .QB (\$dummy [197]), .D (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .CLK (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_7 (.Q (
        L1_0_L2_3_G1_MINI_ALU_BoothP_7), .QB (\$dummy [198]), .D (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .CLK (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_8 (.Q (
        L1_0_L2_3_G1_MINI_ALU_BoothP_8), .QB (\$dummy [199]), .D (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .CLK (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_9 (.Q (
        L1_0_L2_3_G1_MINI_ALU_BoothP_9), .QB (\$dummy [200]), .D (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .CLK (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_10 (.Q (
        L1_0_L2_3_G1_MINI_ALU_BoothP_10), .QB (\$dummy [201]), .D (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .CLK (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_11 (.Q (
        L1_0_L2_3_G1_MINI_ALU_BoothP_11), .QB (\$dummy [202]), .D (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .CLK (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_12 (.Q (
        L1_0_L2_3_G1_MINI_ALU_BoothP_12), .QB (\$dummy [203]), .D (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .CLK (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_13 (.Q (
        L1_0_L2_3_G1_MINI_ALU_BoothP_13), .QB (\$dummy [204]), .D (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .CLK (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_14 (.Q (
        L1_0_L2_3_G1_MINI_ALU_BoothP_14), .QB (\$dummy [205]), .D (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .CLK (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_15 (.Q (
        L1_0_L2_3_G1_MINI_ALU_BoothP_15), .QB (\$dummy [206]), .D (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .CLK (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_16 (.Q (
        L1_0_L2_3_G1_MINI_ALU_BoothP_16), .QB (\$dummy [207]), .D (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .CLK (
        L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    inv02 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix623 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624), .A (CLK)) ;
    inv02 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix625 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626), .A (CLK)) ;
    inv02 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix627 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628), .A (CLK)) ;
    inv02 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix643 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644), .A (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642)) ;
    xor2 L1_0_L2_4_G1_MINI_ALU_ix83 (.Y (L1Results_4__0), .A0 (
         L1SecondOperands_4__0), .A1 (L1FirstOperands_4__0)) ;
    xnor2 L1_0_L2_4_G1_MINI_ALU_ix380 (.Y (L1_0_L2_4_G1_MINI_ALU_nx379), .A0 (
          L1_0_L2_4_G1_MINI_ALU_nx381), .A1 (L1_0_L2_4_G1_MINI_ALU_nx383)) ;
    nand02 L1_0_L2_4_G1_MINI_ALU_ix382 (.Y (L1_0_L2_4_G1_MINI_ALU_nx381), .A0 (
           L1_0_L2_4_G1_MINI_ALU_BoothOperand_0), .A1 (nx7764)) ;
    xnor2 L1_0_L2_4_G1_MINI_ALU_ix384 (.Y (L1_0_L2_4_G1_MINI_ALU_nx383), .A0 (
          L1_0_L2_4_G1_MINI_ALU_BoothOperand_1), .A1 (
          L1_0_L2_4_G1_MINI_ALU_BoothP_1)) ;
    inv01 L1_0_L2_4_G1_MINI_ALU_ix388 (.Y (L1_0_L2_4_G1_MINI_ALU_nx387), .A (
          L1_0_L2_4_G1_MINI_ALU_BoothP_2)) ;
    xnor2 L1_0_L2_4_G1_MINI_ALU_ix390 (.Y (L1_0_L2_4_G1_MINI_ALU_nx389), .A0 (
          L1_0_L2_4_G1_MINI_ALU_nx391), .A1 (L1_0_L2_4_G1_MINI_ALU_nx395)) ;
    aoi32 L1_0_L2_4_G1_MINI_ALU_ix392 (.Y (L1_0_L2_4_G1_MINI_ALU_nx391), .A0 (
          L1_0_L2_4_G1_MINI_ALU_BoothOperand_0), .A1 (nx7764), .A2 (
          L1_0_L2_4_G1_MINI_ALU_nx154), .B0 (L1_0_L2_4_G1_MINI_ALU_BoothP_1), .B1 (
          L1_0_L2_4_G1_MINI_ALU_BoothOperand_1)) ;
    xnor2 L1_0_L2_4_G1_MINI_ALU_ix396 (.Y (L1_0_L2_4_G1_MINI_ALU_nx395), .A0 (
          L1_0_L2_4_G1_MINI_ALU_BoothOperand_2), .A1 (
          L1_0_L2_4_G1_MINI_ALU_BoothP_2)) ;
    inv01 L1_0_L2_4_G1_MINI_ALU_ix400 (.Y (L1_0_L2_4_G1_MINI_ALU_nx399), .A (
          L1_0_L2_4_G1_MINI_ALU_BoothP_3)) ;
    xnor2 L1_0_L2_4_G1_MINI_ALU_ix402 (.Y (L1_0_L2_4_G1_MINI_ALU_nx401), .A0 (
          L1_0_L2_4_G1_MINI_ALU_nx403), .A1 (L1_0_L2_4_G1_MINI_ALU_nx405)) ;
    xnor2 L1_0_L2_4_G1_MINI_ALU_ix406 (.Y (L1_0_L2_4_G1_MINI_ALU_nx405), .A0 (
          L1_0_L2_4_G1_MINI_ALU_BoothOperand_3), .A1 (
          L1_0_L2_4_G1_MINI_ALU_BoothP_3)) ;
    inv01 L1_0_L2_4_G1_MINI_ALU_ix410 (.Y (L1_0_L2_4_G1_MINI_ALU_nx409), .A (
          L1_0_L2_4_G1_MINI_ALU_BoothP_4)) ;
    xnor2 L1_0_L2_4_G1_MINI_ALU_ix412 (.Y (L1_0_L2_4_G1_MINI_ALU_nx411), .A0 (
          L1_0_L2_4_G1_MINI_ALU_nx413), .A1 (L1_0_L2_4_G1_MINI_ALU_nx415)) ;
    xnor2 L1_0_L2_4_G1_MINI_ALU_ix416 (.Y (L1_0_L2_4_G1_MINI_ALU_nx415), .A0 (
          L1_0_L2_4_G1_MINI_ALU_BoothOperand_4), .A1 (
          L1_0_L2_4_G1_MINI_ALU_BoothP_4)) ;
    inv01 L1_0_L2_4_G1_MINI_ALU_ix420 (.Y (L1_0_L2_4_G1_MINI_ALU_nx419), .A (
          L1_0_L2_4_G1_MINI_ALU_BoothP_5)) ;
    xnor2 L1_0_L2_4_G1_MINI_ALU_ix422 (.Y (L1_0_L2_4_G1_MINI_ALU_nx421), .A0 (
          L1_0_L2_4_G1_MINI_ALU_nx423), .A1 (L1_0_L2_4_G1_MINI_ALU_nx425)) ;
    xnor2 L1_0_L2_4_G1_MINI_ALU_ix426 (.Y (L1_0_L2_4_G1_MINI_ALU_nx425), .A0 (
          L1_0_L2_4_G1_MINI_ALU_BoothOperand_5), .A1 (
          L1_0_L2_4_G1_MINI_ALU_BoothP_5)) ;
    inv01 L1_0_L2_4_G1_MINI_ALU_ix430 (.Y (L1_0_L2_4_G1_MINI_ALU_nx429), .A (
          L1_0_L2_4_G1_MINI_ALU_BoothP_6)) ;
    xnor2 L1_0_L2_4_G1_MINI_ALU_ix432 (.Y (L1_0_L2_4_G1_MINI_ALU_nx431), .A0 (
          L1_0_L2_4_G1_MINI_ALU_nx433), .A1 (L1_0_L2_4_G1_MINI_ALU_nx435)) ;
    xnor2 L1_0_L2_4_G1_MINI_ALU_ix436 (.Y (L1_0_L2_4_G1_MINI_ALU_nx435), .A0 (
          L1_0_L2_4_G1_MINI_ALU_BoothOperand_6), .A1 (
          L1_0_L2_4_G1_MINI_ALU_BoothP_6)) ;
    inv01 L1_0_L2_4_G1_MINI_ALU_ix440 (.Y (L1_0_L2_4_G1_MINI_ALU_nx439), .A (
          L1_0_L2_4_G1_MINI_ALU_BoothP_7)) ;
    xnor2 L1_0_L2_4_G1_MINI_ALU_ix442 (.Y (L1_0_L2_4_G1_MINI_ALU_nx441), .A0 (
          L1_0_L2_4_G1_MINI_ALU_nx443), .A1 (L1_0_L2_4_G1_MINI_ALU_nx445)) ;
    xnor2 L1_0_L2_4_G1_MINI_ALU_ix446 (.Y (L1_0_L2_4_G1_MINI_ALU_nx445), .A0 (
          L1_0_L2_4_G1_MINI_ALU_BoothOperand_7), .A1 (
          L1_0_L2_4_G1_MINI_ALU_BoothP_7)) ;
    inv01 L1_0_L2_4_G1_MINI_ALU_ix450 (.Y (L1_0_L2_4_G1_MINI_ALU_nx449), .A (
          L1_0_L2_4_G1_MINI_ALU_BoothP_8)) ;
    xnor2 L1_0_L2_4_G1_MINI_ALU_ix452 (.Y (L1_0_L2_4_G1_MINI_ALU_nx451), .A0 (
          L1_0_L2_4_G1_MINI_ALU_nx453), .A1 (L1_0_L2_4_G1_MINI_ALU_nx455)) ;
    xnor2 L1_0_L2_4_G1_MINI_ALU_ix456 (.Y (L1_0_L2_4_G1_MINI_ALU_nx455), .A0 (
          L1_0_L2_4_G1_MINI_ALU_BoothOperand_8), .A1 (
          L1_0_L2_4_G1_MINI_ALU_BoothP_8)) ;
    xor2 L1_0_L2_4_G1_MINI_ALU_ix317 (.Y (L1_0_L2_4_G1_MINI_ALU_nx316), .A0 (
         L1_0_L2_4_G1_MINI_ALU_nx461), .A1 (L1_0_L2_4_G1_MINI_ALU_nx463)) ;
    xnor2 L1_0_L2_4_G1_MINI_ALU_ix464 (.Y (L1_0_L2_4_G1_MINI_ALU_nx463), .A0 (
          L1_0_L2_4_G1_MINI_ALU_BoothOperand_9), .A1 (
          L1_0_L2_4_G1_MINI_ALU_BoothP_9)) ;
    xor2 L1_0_L2_4_G1_MINI_ALU_ix337 (.Y (L1_0_L2_4_G1_MINI_ALU_nx336), .A0 (
         L1_0_L2_4_G1_MINI_ALU_nx467), .A1 (L1_0_L2_4_G1_MINI_ALU_nx471)) ;
    inv01 L1_0_L2_4_G1_MINI_ALU_ix470 (.Y (L1_0_L2_4_G1_MINI_ALU_nx469), .A (
          L1_0_L2_4_G1_MINI_ALU_BoothP_9)) ;
    xnor2 L1_0_L2_4_G1_MINI_ALU_ix472 (.Y (L1_0_L2_4_G1_MINI_ALU_nx471), .A0 (
          L1_0_L2_4_G1_MINI_ALU_BoothOperand_10), .A1 (
          L1_0_L2_4_G1_MINI_ALU_BoothP_10)) ;
    xor2 L1_0_L2_4_G1_MINI_ALU_ix357 (.Y (L1_0_L2_4_G1_MINI_ALU_nx356), .A0 (
         L1_0_L2_4_G1_MINI_ALU_nx475), .A1 (L1_0_L2_4_G1_MINI_ALU_nx479)) ;
    inv01 L1_0_L2_4_G1_MINI_ALU_ix478 (.Y (L1_0_L2_4_G1_MINI_ALU_nx477), .A (
          L1_0_L2_4_G1_MINI_ALU_BoothP_10)) ;
    xnor2 L1_0_L2_4_G1_MINI_ALU_ix480 (.Y (L1_0_L2_4_G1_MINI_ALU_nx479), .A0 (
          L1_0_L2_4_G1_MINI_ALU_BoothOperand_11), .A1 (
          L1_0_L2_4_G1_MINI_ALU_BoothP_11)) ;
    xor2 L1_0_L2_4_G1_MINI_ALU_ix377 (.Y (L1_0_L2_4_G1_MINI_ALU_nx376), .A0 (
         L1_0_L2_4_G1_MINI_ALU_nx483), .A1 (L1_0_L2_4_G1_MINI_ALU_nx487)) ;
    inv01 L1_0_L2_4_G1_MINI_ALU_ix486 (.Y (L1_0_L2_4_G1_MINI_ALU_nx485), .A (
          L1_0_L2_4_G1_MINI_ALU_BoothP_11)) ;
    xnor2 L1_0_L2_4_G1_MINI_ALU_ix488 (.Y (L1_0_L2_4_G1_MINI_ALU_nx487), .A0 (
          L1_0_L2_4_G1_MINI_ALU_BoothOperand_12), .A1 (
          L1_0_L2_4_G1_MINI_ALU_BoothP_12)) ;
    xor2 L1_0_L2_4_G1_MINI_ALU_ix397 (.Y (L1_0_L2_4_G1_MINI_ALU_nx396), .A0 (
         L1_0_L2_4_G1_MINI_ALU_nx491), .A1 (L1_0_L2_4_G1_MINI_ALU_nx495)) ;
    inv01 L1_0_L2_4_G1_MINI_ALU_ix494 (.Y (L1_0_L2_4_G1_MINI_ALU_nx493), .A (
          L1_0_L2_4_G1_MINI_ALU_BoothP_12)) ;
    xnor2 L1_0_L2_4_G1_MINI_ALU_ix496 (.Y (L1_0_L2_4_G1_MINI_ALU_nx495), .A0 (
          L1_0_L2_4_G1_MINI_ALU_BoothOperand_13), .A1 (
          L1_0_L2_4_G1_MINI_ALU_BoothP_13)) ;
    xor2 L1_0_L2_4_G1_MINI_ALU_ix417 (.Y (L1_0_L2_4_G1_MINI_ALU_nx416), .A0 (
         L1_0_L2_4_G1_MINI_ALU_nx499), .A1 (L1_0_L2_4_G1_MINI_ALU_nx503)) ;
    inv01 L1_0_L2_4_G1_MINI_ALU_ix502 (.Y (L1_0_L2_4_G1_MINI_ALU_nx501), .A (
          L1_0_L2_4_G1_MINI_ALU_BoothP_13)) ;
    xnor2 L1_0_L2_4_G1_MINI_ALU_ix504 (.Y (L1_0_L2_4_G1_MINI_ALU_nx503), .A0 (
          L1_0_L2_4_G1_MINI_ALU_BoothOperand_14), .A1 (
          L1_0_L2_4_G1_MINI_ALU_BoothP_14)) ;
    xor2 L1_0_L2_4_G1_MINI_ALU_ix437 (.Y (L1_0_L2_4_G1_MINI_ALU_nx436), .A0 (
         L1_0_L2_4_G1_MINI_ALU_nx507), .A1 (L1_0_L2_4_G1_MINI_ALU_nx511)) ;
    inv01 L1_0_L2_4_G1_MINI_ALU_ix510 (.Y (L1_0_L2_4_G1_MINI_ALU_nx509), .A (
          L1_0_L2_4_G1_MINI_ALU_BoothP_14)) ;
    xnor2 L1_0_L2_4_G1_MINI_ALU_ix512 (.Y (L1_0_L2_4_G1_MINI_ALU_nx511), .A0 (
          L1_0_L2_4_G1_MINI_ALU_BoothOperand_15), .A1 (
          L1_0_L2_4_G1_MINI_ALU_BoothP_15)) ;
    xnor2 L1_0_L2_4_G1_MINI_ALU_ix457 (.Y (L1_0_L2_4_G1_MINI_ALU_nx456), .A0 (
          L1_0_L2_4_G1_MINI_ALU_nx515), .A1 (L1_0_L2_4_G1_MINI_ALU_nx454)) ;
    inv01 L1_0_L2_4_G1_MINI_ALU_ix518 (.Y (L1_0_L2_4_G1_MINI_ALU_nx517), .A (
          L1_0_L2_4_G1_MINI_ALU_BoothP_15)) ;
    xor2 L1_0_L2_4_G1_MINI_ALU_ix455 (.Y (L1_0_L2_4_G1_MINI_ALU_nx454), .A0 (
         L1_0_L2_4_G1_MINI_ALU_BoothOperand_16), .A1 (
         L1_0_L2_4_G1_MINI_ALU_BoothP_16)) ;
    mux21_ni L1_0_L2_4_G1_MINI_ALU_ix91 (.Y (L1SecondOperands_4__0), .A0 (
             L1_0_L2_4_G1_MINI_ALU_BoothP_1), .A1 (WindowDin_0__4__0), .S0 (
             Instr)) ;
    mux21_ni L1_0_L2_4_G1_MINI_ALU_ix99 (.Y (L1SecondOperands_4__1), .A0 (
             L1_0_L2_4_G1_MINI_ALU_BoothP_2), .A1 (WindowDin_0__4__1), .S0 (
             Instr)) ;
    mux21_ni L1_0_L2_4_G1_MINI_ALU_ix107 (.Y (L1SecondOperands_4__2), .A0 (
             L1_0_L2_4_G1_MINI_ALU_BoothP_3), .A1 (WindowDin_0__4__2), .S0 (
             Instr)) ;
    mux21_ni L1_0_L2_4_G1_MINI_ALU_ix115 (.Y (L1SecondOperands_4__3), .A0 (
             L1_0_L2_4_G1_MINI_ALU_BoothP_4), .A1 (WindowDin_0__4__3), .S0 (
             Instr)) ;
    mux21_ni L1_0_L2_4_G1_MINI_ALU_ix123 (.Y (L1SecondOperands_4__4), .A0 (
             L1_0_L2_4_G1_MINI_ALU_BoothP_5), .A1 (WindowDin_0__4__4), .S0 (
             Instr)) ;
    mux21_ni L1_0_L2_4_G1_MINI_ALU_ix131 (.Y (L1SecondOperands_4__5), .A0 (
             L1_0_L2_4_G1_MINI_ALU_BoothP_6), .A1 (WindowDin_0__4__5), .S0 (
             Instr)) ;
    mux21_ni L1_0_L2_4_G1_MINI_ALU_ix139 (.Y (L1SecondOperands_4__6), .A0 (
             L1_0_L2_4_G1_MINI_ALU_BoothP_7), .A1 (WindowDin_0__4__6), .S0 (
             Instr)) ;
    mux21_ni L1_0_L2_4_G1_MINI_ALU_ix147 (.Y (L1SecondOperands_4__7), .A0 (
             L1_0_L2_4_G1_MINI_ALU_BoothP_8), .A1 (WindowDin_0__4__7), .S0 (
             Instr)) ;
    xor2 L1_0_L2_4_G1_MINI_ALU_ix77 (.Y (L1Results_4__1), .A0 (
         L1_0_L2_4_G1_MINI_ALU_nx529), .A1 (L1_0_L2_4_G1_MINI_ALU_nx531)) ;
    nand02 L1_0_L2_4_G1_MINI_ALU_ix530 (.Y (L1_0_L2_4_G1_MINI_ALU_nx529), .A0 (
           L1SecondOperands_4__0), .A1 (L1FirstOperands_4__0)) ;
    xnor2 L1_0_L2_4_G1_MINI_ALU_ix532 (.Y (L1_0_L2_4_G1_MINI_ALU_nx531), .A0 (
          L1SecondOperands_4__1), .A1 (L1FirstOperands_4__1)) ;
    xor2 L1_0_L2_4_G1_MINI_ALU_ix75 (.Y (L1Results_4__2), .A0 (
         L1_0_L2_4_G1_MINI_ALU_nx534), .A1 (L1_0_L2_4_G1_MINI_ALU_nx537)) ;
    aoi32 L1_0_L2_4_G1_MINI_ALU_ix535 (.Y (L1_0_L2_4_G1_MINI_ALU_nx534), .A0 (
          L1SecondOperands_4__0), .A1 (L1FirstOperands_4__0), .A2 (
          L1_0_L2_4_G1_MINI_ALU_nx30), .B0 (L1FirstOperands_4__1), .B1 (
          L1SecondOperands_4__1)) ;
    xnor2 L1_0_L2_4_G1_MINI_ALU_ix538 (.Y (L1_0_L2_4_G1_MINI_ALU_nx537), .A0 (
          L1SecondOperands_4__2), .A1 (L1FirstOperands_4__2)) ;
    xor2 L1_0_L2_4_G1_MINI_ALU_ix73 (.Y (L1Results_4__3), .A0 (
         L1_0_L2_4_G1_MINI_ALU_nx540), .A1 (L1_0_L2_4_G1_MINI_ALU_nx544)) ;
    aoi22 L1_0_L2_4_G1_MINI_ALU_ix541 (.Y (L1_0_L2_4_G1_MINI_ALU_nx540), .A0 (
          L1FirstOperands_4__2), .A1 (L1SecondOperands_4__2), .B0 (
          L1_0_L2_4_G1_MINI_ALU_nx40), .B1 (L1_0_L2_4_G1_MINI_ALU_nx24)) ;
    xnor2 L1_0_L2_4_G1_MINI_ALU_ix545 (.Y (L1_0_L2_4_G1_MINI_ALU_nx544), .A0 (
          L1SecondOperands_4__3), .A1 (L1FirstOperands_4__3)) ;
    xor2 L1_0_L2_4_G1_MINI_ALU_ix71 (.Y (L1Results_4__4), .A0 (
         L1_0_L2_4_G1_MINI_ALU_nx547), .A1 (L1_0_L2_4_G1_MINI_ALU_nx551)) ;
    aoi22 L1_0_L2_4_G1_MINI_ALU_ix548 (.Y (L1_0_L2_4_G1_MINI_ALU_nx547), .A0 (
          L1FirstOperands_4__3), .A1 (L1SecondOperands_4__3), .B0 (
          L1_0_L2_4_G1_MINI_ALU_nx44), .B1 (L1_0_L2_4_G1_MINI_ALU_nx18)) ;
    xnor2 L1_0_L2_4_G1_MINI_ALU_ix552 (.Y (L1_0_L2_4_G1_MINI_ALU_nx551), .A0 (
          L1SecondOperands_4__4), .A1 (L1FirstOperands_4__4)) ;
    xor2 L1_0_L2_4_G1_MINI_ALU_ix69 (.Y (L1Results_4__5), .A0 (
         L1_0_L2_4_G1_MINI_ALU_nx554), .A1 (L1_0_L2_4_G1_MINI_ALU_nx558)) ;
    aoi22 L1_0_L2_4_G1_MINI_ALU_ix555 (.Y (L1_0_L2_4_G1_MINI_ALU_nx554), .A0 (
          L1FirstOperands_4__4), .A1 (L1SecondOperands_4__4), .B0 (
          L1_0_L2_4_G1_MINI_ALU_nx48), .B1 (L1_0_L2_4_G1_MINI_ALU_nx12)) ;
    xnor2 L1_0_L2_4_G1_MINI_ALU_ix559 (.Y (L1_0_L2_4_G1_MINI_ALU_nx558), .A0 (
          L1SecondOperands_4__5), .A1 (L1FirstOperands_4__5)) ;
    xor2 L1_0_L2_4_G1_MINI_ALU_ix67 (.Y (L1Results_4__6), .A0 (
         L1_0_L2_4_G1_MINI_ALU_nx561), .A1 (L1_0_L2_4_G1_MINI_ALU_nx565)) ;
    aoi22 L1_0_L2_4_G1_MINI_ALU_ix562 (.Y (L1_0_L2_4_G1_MINI_ALU_nx561), .A0 (
          L1FirstOperands_4__5), .A1 (L1SecondOperands_4__5), .B0 (
          L1_0_L2_4_G1_MINI_ALU_nx52), .B1 (L1_0_L2_4_G1_MINI_ALU_nx6)) ;
    xnor2 L1_0_L2_4_G1_MINI_ALU_ix566 (.Y (L1_0_L2_4_G1_MINI_ALU_nx565), .A0 (
          L1SecondOperands_4__6), .A1 (L1FirstOperands_4__6)) ;
    xnor2 L1_0_L2_4_G1_MINI_ALU_ix65 (.Y (L1Results_4__7), .A0 (
          L1_0_L2_4_G1_MINI_ALU_nx568), .A1 (L1_0_L2_4_G1_MINI_ALU_nx62)) ;
    aoi22 L1_0_L2_4_G1_MINI_ALU_ix569 (.Y (L1_0_L2_4_G1_MINI_ALU_nx568), .A0 (
          L1FirstOperands_4__6), .A1 (L1SecondOperands_4__6), .B0 (
          L1_0_L2_4_G1_MINI_ALU_nx56), .B1 (L1_0_L2_4_G1_MINI_ALU_nx0)) ;
    xor2 L1_0_L2_4_G1_MINI_ALU_ix63 (.Y (L1_0_L2_4_G1_MINI_ALU_nx62), .A0 (
         L1SecondOperands_4__7), .A1 (L1FirstOperands_4__7)) ;
    inv01 L1_0_L2_4_G1_MINI_ALU_ix155 (.Y (L1_0_L2_4_G1_MINI_ALU_nx154), .A (
          L1_0_L2_4_G1_MINI_ALU_nx383)) ;
    inv01 L1_0_L2_4_G1_MINI_ALU_ix57 (.Y (L1_0_L2_4_G1_MINI_ALU_nx56), .A (
          L1_0_L2_4_G1_MINI_ALU_nx561)) ;
    inv01 L1_0_L2_4_G1_MINI_ALU_ix53 (.Y (L1_0_L2_4_G1_MINI_ALU_nx52), .A (
          L1_0_L2_4_G1_MINI_ALU_nx554)) ;
    inv01 L1_0_L2_4_G1_MINI_ALU_ix49 (.Y (L1_0_L2_4_G1_MINI_ALU_nx48), .A (
          L1_0_L2_4_G1_MINI_ALU_nx547)) ;
    inv01 L1_0_L2_4_G1_MINI_ALU_ix45 (.Y (L1_0_L2_4_G1_MINI_ALU_nx44), .A (
          L1_0_L2_4_G1_MINI_ALU_nx540)) ;
    inv01 L1_0_L2_4_G1_MINI_ALU_ix41 (.Y (L1_0_L2_4_G1_MINI_ALU_nx40), .A (
          L1_0_L2_4_G1_MINI_ALU_nx534)) ;
    inv01 L1_0_L2_4_G1_MINI_ALU_ix31 (.Y (L1_0_L2_4_G1_MINI_ALU_nx30), .A (
          L1_0_L2_4_G1_MINI_ALU_nx531)) ;
    inv01 L1_0_L2_4_G1_MINI_ALU_ix25 (.Y (L1_0_L2_4_G1_MINI_ALU_nx24), .A (
          L1_0_L2_4_G1_MINI_ALU_nx537)) ;
    inv01 L1_0_L2_4_G1_MINI_ALU_ix19 (.Y (L1_0_L2_4_G1_MINI_ALU_nx18), .A (
          L1_0_L2_4_G1_MINI_ALU_nx544)) ;
    inv01 L1_0_L2_4_G1_MINI_ALU_ix13 (.Y (L1_0_L2_4_G1_MINI_ALU_nx12), .A (
          L1_0_L2_4_G1_MINI_ALU_nx551)) ;
    inv01 L1_0_L2_4_G1_MINI_ALU_ix7 (.Y (L1_0_L2_4_G1_MINI_ALU_nx6), .A (
          L1_0_L2_4_G1_MINI_ALU_nx558)) ;
    inv01 L1_0_L2_4_G1_MINI_ALU_ix1 (.Y (L1_0_L2_4_G1_MINI_ALU_nx0), .A (
          L1_0_L2_4_G1_MINI_ALU_nx565)) ;
    fake_gnd L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix216 (.Y (
             L1_0_L2_4_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    nor02ii L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix81 (.Y (
            L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx80), .A0 (Instr), .A1 (Start)) ;
    aoi21 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix77 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_10), .A0 (
          FilterDin_0__4__1), .A1 (FilterDin_0__4__0), .B0 (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx4)) ;
    nor02_2x L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix5 (.Y (
             L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx4), .A0 (FilterDin_0__4__0), .A1 (
             FilterDin_0__4__1)) ;
    aoi21 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix67 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_11), .A0 (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx328), .A1 (FilterDin_0__4__2), .B0 (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx8)) ;
    nor03_2x L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix9 (.Y (
             L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx8), .A0 (FilterDin_0__4__2), .A1 (
             FilterDin_0__4__0), .A2 (FilterDin_0__4__1)) ;
    xnor2 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix59 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_12), .A0 (
          FilterDin_0__4__3), .A1 (L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx8)) ;
    xnor2 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix51 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_13), .A0 (
          FilterDin_0__4__4), .A1 (L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx12)) ;
    nor04 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix13 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx12), .A0 (FilterDin_0__4__3), .A1 (
          FilterDin_0__4__2), .A2 (FilterDin_0__4__0), .A3 (FilterDin_0__4__1)
          ) ;
    xnor2 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix43 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_14), .A0 (
          FilterDin_0__4__5), .A1 (L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx16)) ;
    nor02ii L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix17 (.Y (
            L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx16), .A0 (FilterDin_0__4__4), .A1 (
            L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx12)) ;
    xnor2 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix35 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_15), .A0 (
          FilterDin_0__4__6), .A1 (L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx20)) ;
    nor02ii L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix21 (.Y (
            L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx20), .A0 (FilterDin_0__4__5), .A1 (
            L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx16)) ;
    xnor2 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix27 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_16), .A0 (
          FilterDin_0__4__7), .A1 (L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx24)) ;
    nor02ii L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix25 (.Y (
            L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx24), .A0 (FilterDin_0__4__6), .A1 (
            L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx20)) ;
    inv01 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix329 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx328), .A (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx4)) ;
    inv02 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix383 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx384), .A (
          L1_0_L2_4_G1_MINI_ALU_BoothP_0)) ;
    dff L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_0 (.Q (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_0), .QB (\$dummy [208]), 
        .D (L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .CLK (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    nor02_2x L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix567 (.Y (
             L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566), .A0 (RST), .A1 (
             L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644)) ;
    dff L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_1 (.Q (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_1), .QB (\$dummy [209]), 
        .D (L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .CLK (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_2 (.Q (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_2), .QB (\$dummy [210]), 
        .D (L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .CLK (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_3 (.Q (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_3), .QB (\$dummy [211]), 
        .D (L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .CLK (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_4 (.Q (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_4), .QB (\$dummy [212]), 
        .D (L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .CLK (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_5 (.Q (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_5), .QB (\$dummy [213]), 
        .D (L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .CLK (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_6 (.Q (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_6), .QB (\$dummy [214]), 
        .D (L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .CLK (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_7 (.Q (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_7), .QB (\$dummy [215]), 
        .D (L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .CLK (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_8 (.Q (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_8), .QB (\$dummy [216]), 
        .D (L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .CLK (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_9 (.Q (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_9), .QB (\$dummy [217]), 
        .D (L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .CLK (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_10 (.Q (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_10), .QB (\$dummy [218])
        , .D (L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .CLK (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_11 (.Q (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_11), .QB (\$dummy [219])
        , .D (L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .CLK (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_12 (.Q (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_12), .QB (\$dummy [220])
        , .D (L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .CLK (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_13 (.Q (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_13), .QB (\$dummy [221])
        , .D (L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .CLK (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_14 (.Q (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_14), .QB (\$dummy [222])
        , .D (L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .CLK (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_15 (.Q (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_15), .QB (\$dummy [223])
        , .D (L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .CLK (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_16 (.Q (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_16), .QB (\$dummy [224])
        , .D (L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .CLK (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    inv02 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix623 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624), .A (CLK)) ;
    inv02 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix625 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626), .A (CLK)) ;
    inv02 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix627 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628), .A (CLK)) ;
    inv02 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix643 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644), .A (nx7778)) ;
    dff L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_0 (.Q (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_0), .QB (\$dummy [225]), 
        .D (L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .CLK (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    nor02_2x L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix567 (.Y (
             L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566), .A0 (RST), .A1 (
             L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644)) ;
    dff L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_1 (.Q (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_1), .QB (\$dummy [226]), 
        .D (L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .CLK (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_2 (.Q (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_2), .QB (\$dummy [227]), 
        .D (L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .CLK (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_3 (.Q (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_3), .QB (\$dummy [228]), 
        .D (L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .CLK (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_4 (.Q (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_4), .QB (\$dummy [229]), 
        .D (L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .CLK (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_5 (.Q (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_5), .QB (\$dummy [230]), 
        .D (L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .CLK (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_6 (.Q (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_6), .QB (\$dummy [231]), 
        .D (L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .CLK (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_7 (.Q (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_7), .QB (\$dummy [232]), 
        .D (L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .CLK (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_8 (.Q (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_8), .QB (\$dummy [233]), 
        .D (L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .CLK (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_9 (.Q (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_9), .QB (\$dummy [234]), 
        .D (L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .CLK (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_10 (.Q (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_10), .QB (\$dummy [235])
        , .D (L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .CLK (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_11 (.Q (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_11), .QB (\$dummy [236])
        , .D (L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .CLK (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_12 (.Q (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_12), .QB (\$dummy [237])
        , .D (L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .CLK (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_13 (.Q (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_13), .QB (\$dummy [238])
        , .D (L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .CLK (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_14 (.Q (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_14), .QB (\$dummy [239])
        , .D (L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .CLK (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_15 (.Q (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_15), .QB (\$dummy [240])
        , .D (L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .CLK (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_16 (.Q (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_16), .QB (\$dummy [241])
        , .D (L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .CLK (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    inv02 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix623 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624), .A (CLK)) ;
    inv02 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix625 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626), .A (CLK)) ;
    inv02 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix627 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628), .A (CLK)) ;
    inv02 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix643 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644), .A (nx7784)) ;
    dff L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_0 (.Q (
        L1_0_L2_4_G1_MINI_ALU_BoothP_0), .QB (\$dummy [242]), .D (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .CLK (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    nor02_2x L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix567 (.Y (
             L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566), .A0 (RST), .A1 (
             L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    dff L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_1 (.Q (
        L1_0_L2_4_G1_MINI_ALU_BoothP_1), .QB (\$dummy [243]), .D (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .CLK (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_2 (.Q (
        L1_0_L2_4_G1_MINI_ALU_BoothP_2), .QB (\$dummy [244]), .D (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .CLK (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_3 (.Q (
        L1_0_L2_4_G1_MINI_ALU_BoothP_3), .QB (\$dummy [245]), .D (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .CLK (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_4 (.Q (
        L1_0_L2_4_G1_MINI_ALU_BoothP_4), .QB (\$dummy [246]), .D (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .CLK (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_5 (.Q (
        L1_0_L2_4_G1_MINI_ALU_BoothP_5), .QB (\$dummy [247]), .D (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .CLK (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_6 (.Q (
        L1_0_L2_4_G1_MINI_ALU_BoothP_6), .QB (\$dummy [248]), .D (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .CLK (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_7 (.Q (
        L1_0_L2_4_G1_MINI_ALU_BoothP_7), .QB (\$dummy [249]), .D (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .CLK (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_8 (.Q (
        L1_0_L2_4_G1_MINI_ALU_BoothP_8), .QB (\$dummy [250]), .D (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .CLK (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_9 (.Q (
        L1_0_L2_4_G1_MINI_ALU_BoothP_9), .QB (\$dummy [251]), .D (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .CLK (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_10 (.Q (
        L1_0_L2_4_G1_MINI_ALU_BoothP_10), .QB (\$dummy [252]), .D (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .CLK (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_11 (.Q (
        L1_0_L2_4_G1_MINI_ALU_BoothP_11), .QB (\$dummy [253]), .D (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .CLK (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_12 (.Q (
        L1_0_L2_4_G1_MINI_ALU_BoothP_12), .QB (\$dummy [254]), .D (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .CLK (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_13 (.Q (
        L1_0_L2_4_G1_MINI_ALU_BoothP_13), .QB (\$dummy [255]), .D (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .CLK (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_14 (.Q (
        L1_0_L2_4_G1_MINI_ALU_BoothP_14), .QB (\$dummy [256]), .D (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .CLK (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_15 (.Q (
        L1_0_L2_4_G1_MINI_ALU_BoothP_15), .QB (\$dummy [257]), .D (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .CLK (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_16 (.Q (
        L1_0_L2_4_G1_MINI_ALU_BoothP_16), .QB (\$dummy [258]), .D (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .CLK (
        L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    inv02 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix623 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624), .A (CLK)) ;
    inv02 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix625 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626), .A (CLK)) ;
    inv02 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix627 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628), .A (CLK)) ;
    inv02 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix643 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644), .A (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642)) ;
    xor2 L1_1_L2_0_G1_MINI_ALU_ix83 (.Y (L1Results_5__0), .A0 (
         L1SecondOperands_5__0), .A1 (L1FirstOperands_5__0)) ;
    xnor2 L1_1_L2_0_G1_MINI_ALU_ix380 (.Y (L1_1_L2_0_G1_MINI_ALU_nx379), .A0 (
          L1_1_L2_0_G1_MINI_ALU_nx381), .A1 (L1_1_L2_0_G1_MINI_ALU_nx383)) ;
    nand02 L1_1_L2_0_G1_MINI_ALU_ix382 (.Y (L1_1_L2_0_G1_MINI_ALU_nx381), .A0 (
           L1_1_L2_0_G1_MINI_ALU_BoothOperand_0), .A1 (nx7804)) ;
    xnor2 L1_1_L2_0_G1_MINI_ALU_ix384 (.Y (L1_1_L2_0_G1_MINI_ALU_nx383), .A0 (
          L1_1_L2_0_G1_MINI_ALU_BoothOperand_1), .A1 (
          L1_1_L2_0_G1_MINI_ALU_BoothP_1)) ;
    inv01 L1_1_L2_0_G1_MINI_ALU_ix388 (.Y (L1_1_L2_0_G1_MINI_ALU_nx387), .A (
          L1_1_L2_0_G1_MINI_ALU_BoothP_2)) ;
    xnor2 L1_1_L2_0_G1_MINI_ALU_ix390 (.Y (L1_1_L2_0_G1_MINI_ALU_nx389), .A0 (
          L1_1_L2_0_G1_MINI_ALU_nx391), .A1 (L1_1_L2_0_G1_MINI_ALU_nx395)) ;
    aoi32 L1_1_L2_0_G1_MINI_ALU_ix392 (.Y (L1_1_L2_0_G1_MINI_ALU_nx391), .A0 (
          L1_1_L2_0_G1_MINI_ALU_BoothOperand_0), .A1 (nx7804), .A2 (
          L1_1_L2_0_G1_MINI_ALU_nx154), .B0 (L1_1_L2_0_G1_MINI_ALU_BoothP_1), .B1 (
          L1_1_L2_0_G1_MINI_ALU_BoothOperand_1)) ;
    xnor2 L1_1_L2_0_G1_MINI_ALU_ix396 (.Y (L1_1_L2_0_G1_MINI_ALU_nx395), .A0 (
          L1_1_L2_0_G1_MINI_ALU_BoothOperand_2), .A1 (
          L1_1_L2_0_G1_MINI_ALU_BoothP_2)) ;
    inv01 L1_1_L2_0_G1_MINI_ALU_ix400 (.Y (L1_1_L2_0_G1_MINI_ALU_nx399), .A (
          L1_1_L2_0_G1_MINI_ALU_BoothP_3)) ;
    xnor2 L1_1_L2_0_G1_MINI_ALU_ix402 (.Y (L1_1_L2_0_G1_MINI_ALU_nx401), .A0 (
          L1_1_L2_0_G1_MINI_ALU_nx403), .A1 (L1_1_L2_0_G1_MINI_ALU_nx405)) ;
    xnor2 L1_1_L2_0_G1_MINI_ALU_ix406 (.Y (L1_1_L2_0_G1_MINI_ALU_nx405), .A0 (
          L1_1_L2_0_G1_MINI_ALU_BoothOperand_3), .A1 (
          L1_1_L2_0_G1_MINI_ALU_BoothP_3)) ;
    inv01 L1_1_L2_0_G1_MINI_ALU_ix410 (.Y (L1_1_L2_0_G1_MINI_ALU_nx409), .A (
          L1_1_L2_0_G1_MINI_ALU_BoothP_4)) ;
    xnor2 L1_1_L2_0_G1_MINI_ALU_ix412 (.Y (L1_1_L2_0_G1_MINI_ALU_nx411), .A0 (
          L1_1_L2_0_G1_MINI_ALU_nx413), .A1 (L1_1_L2_0_G1_MINI_ALU_nx415)) ;
    xnor2 L1_1_L2_0_G1_MINI_ALU_ix416 (.Y (L1_1_L2_0_G1_MINI_ALU_nx415), .A0 (
          L1_1_L2_0_G1_MINI_ALU_BoothOperand_4), .A1 (
          L1_1_L2_0_G1_MINI_ALU_BoothP_4)) ;
    inv01 L1_1_L2_0_G1_MINI_ALU_ix420 (.Y (L1_1_L2_0_G1_MINI_ALU_nx419), .A (
          L1_1_L2_0_G1_MINI_ALU_BoothP_5)) ;
    xnor2 L1_1_L2_0_G1_MINI_ALU_ix422 (.Y (L1_1_L2_0_G1_MINI_ALU_nx421), .A0 (
          L1_1_L2_0_G1_MINI_ALU_nx423), .A1 (L1_1_L2_0_G1_MINI_ALU_nx425)) ;
    xnor2 L1_1_L2_0_G1_MINI_ALU_ix426 (.Y (L1_1_L2_0_G1_MINI_ALU_nx425), .A0 (
          L1_1_L2_0_G1_MINI_ALU_BoothOperand_5), .A1 (
          L1_1_L2_0_G1_MINI_ALU_BoothP_5)) ;
    inv01 L1_1_L2_0_G1_MINI_ALU_ix430 (.Y (L1_1_L2_0_G1_MINI_ALU_nx429), .A (
          L1_1_L2_0_G1_MINI_ALU_BoothP_6)) ;
    xnor2 L1_1_L2_0_G1_MINI_ALU_ix432 (.Y (L1_1_L2_0_G1_MINI_ALU_nx431), .A0 (
          L1_1_L2_0_G1_MINI_ALU_nx433), .A1 (L1_1_L2_0_G1_MINI_ALU_nx435)) ;
    xnor2 L1_1_L2_0_G1_MINI_ALU_ix436 (.Y (L1_1_L2_0_G1_MINI_ALU_nx435), .A0 (
          L1_1_L2_0_G1_MINI_ALU_BoothOperand_6), .A1 (
          L1_1_L2_0_G1_MINI_ALU_BoothP_6)) ;
    inv01 L1_1_L2_0_G1_MINI_ALU_ix440 (.Y (L1_1_L2_0_G1_MINI_ALU_nx439), .A (
          L1_1_L2_0_G1_MINI_ALU_BoothP_7)) ;
    xnor2 L1_1_L2_0_G1_MINI_ALU_ix442 (.Y (L1_1_L2_0_G1_MINI_ALU_nx441), .A0 (
          L1_1_L2_0_G1_MINI_ALU_nx443), .A1 (L1_1_L2_0_G1_MINI_ALU_nx445)) ;
    xnor2 L1_1_L2_0_G1_MINI_ALU_ix446 (.Y (L1_1_L2_0_G1_MINI_ALU_nx445), .A0 (
          L1_1_L2_0_G1_MINI_ALU_BoothOperand_7), .A1 (
          L1_1_L2_0_G1_MINI_ALU_BoothP_7)) ;
    inv01 L1_1_L2_0_G1_MINI_ALU_ix450 (.Y (L1_1_L2_0_G1_MINI_ALU_nx449), .A (
          L1_1_L2_0_G1_MINI_ALU_BoothP_8)) ;
    xnor2 L1_1_L2_0_G1_MINI_ALU_ix452 (.Y (L1_1_L2_0_G1_MINI_ALU_nx451), .A0 (
          L1_1_L2_0_G1_MINI_ALU_nx453), .A1 (L1_1_L2_0_G1_MINI_ALU_nx455)) ;
    xnor2 L1_1_L2_0_G1_MINI_ALU_ix456 (.Y (L1_1_L2_0_G1_MINI_ALU_nx455), .A0 (
          L1_1_L2_0_G1_MINI_ALU_BoothOperand_8), .A1 (
          L1_1_L2_0_G1_MINI_ALU_BoothP_8)) ;
    xor2 L1_1_L2_0_G1_MINI_ALU_ix317 (.Y (L1_1_L2_0_G1_MINI_ALU_nx316), .A0 (
         L1_1_L2_0_G1_MINI_ALU_nx461), .A1 (L1_1_L2_0_G1_MINI_ALU_nx463)) ;
    xnor2 L1_1_L2_0_G1_MINI_ALU_ix464 (.Y (L1_1_L2_0_G1_MINI_ALU_nx463), .A0 (
          L1_1_L2_0_G1_MINI_ALU_BoothOperand_9), .A1 (
          L1_1_L2_0_G1_MINI_ALU_BoothP_9)) ;
    xor2 L1_1_L2_0_G1_MINI_ALU_ix337 (.Y (L1_1_L2_0_G1_MINI_ALU_nx336), .A0 (
         L1_1_L2_0_G1_MINI_ALU_nx467), .A1 (L1_1_L2_0_G1_MINI_ALU_nx471)) ;
    inv01 L1_1_L2_0_G1_MINI_ALU_ix470 (.Y (L1_1_L2_0_G1_MINI_ALU_nx469), .A (
          L1_1_L2_0_G1_MINI_ALU_BoothP_9)) ;
    xnor2 L1_1_L2_0_G1_MINI_ALU_ix472 (.Y (L1_1_L2_0_G1_MINI_ALU_nx471), .A0 (
          L1_1_L2_0_G1_MINI_ALU_BoothOperand_10), .A1 (
          L1_1_L2_0_G1_MINI_ALU_BoothP_10)) ;
    xor2 L1_1_L2_0_G1_MINI_ALU_ix357 (.Y (L1_1_L2_0_G1_MINI_ALU_nx356), .A0 (
         L1_1_L2_0_G1_MINI_ALU_nx475), .A1 (L1_1_L2_0_G1_MINI_ALU_nx479)) ;
    inv01 L1_1_L2_0_G1_MINI_ALU_ix478 (.Y (L1_1_L2_0_G1_MINI_ALU_nx477), .A (
          L1_1_L2_0_G1_MINI_ALU_BoothP_10)) ;
    xnor2 L1_1_L2_0_G1_MINI_ALU_ix480 (.Y (L1_1_L2_0_G1_MINI_ALU_nx479), .A0 (
          L1_1_L2_0_G1_MINI_ALU_BoothOperand_11), .A1 (
          L1_1_L2_0_G1_MINI_ALU_BoothP_11)) ;
    xor2 L1_1_L2_0_G1_MINI_ALU_ix377 (.Y (L1_1_L2_0_G1_MINI_ALU_nx376), .A0 (
         L1_1_L2_0_G1_MINI_ALU_nx483), .A1 (L1_1_L2_0_G1_MINI_ALU_nx487)) ;
    inv01 L1_1_L2_0_G1_MINI_ALU_ix486 (.Y (L1_1_L2_0_G1_MINI_ALU_nx485), .A (
          L1_1_L2_0_G1_MINI_ALU_BoothP_11)) ;
    xnor2 L1_1_L2_0_G1_MINI_ALU_ix488 (.Y (L1_1_L2_0_G1_MINI_ALU_nx487), .A0 (
          L1_1_L2_0_G1_MINI_ALU_BoothOperand_12), .A1 (
          L1_1_L2_0_G1_MINI_ALU_BoothP_12)) ;
    xor2 L1_1_L2_0_G1_MINI_ALU_ix397 (.Y (L1_1_L2_0_G1_MINI_ALU_nx396), .A0 (
         L1_1_L2_0_G1_MINI_ALU_nx491), .A1 (L1_1_L2_0_G1_MINI_ALU_nx495)) ;
    inv01 L1_1_L2_0_G1_MINI_ALU_ix494 (.Y (L1_1_L2_0_G1_MINI_ALU_nx493), .A (
          L1_1_L2_0_G1_MINI_ALU_BoothP_12)) ;
    xnor2 L1_1_L2_0_G1_MINI_ALU_ix496 (.Y (L1_1_L2_0_G1_MINI_ALU_nx495), .A0 (
          L1_1_L2_0_G1_MINI_ALU_BoothOperand_13), .A1 (
          L1_1_L2_0_G1_MINI_ALU_BoothP_13)) ;
    xor2 L1_1_L2_0_G1_MINI_ALU_ix417 (.Y (L1_1_L2_0_G1_MINI_ALU_nx416), .A0 (
         L1_1_L2_0_G1_MINI_ALU_nx499), .A1 (L1_1_L2_0_G1_MINI_ALU_nx503)) ;
    inv01 L1_1_L2_0_G1_MINI_ALU_ix502 (.Y (L1_1_L2_0_G1_MINI_ALU_nx501), .A (
          L1_1_L2_0_G1_MINI_ALU_BoothP_13)) ;
    xnor2 L1_1_L2_0_G1_MINI_ALU_ix504 (.Y (L1_1_L2_0_G1_MINI_ALU_nx503), .A0 (
          L1_1_L2_0_G1_MINI_ALU_BoothOperand_14), .A1 (
          L1_1_L2_0_G1_MINI_ALU_BoothP_14)) ;
    xor2 L1_1_L2_0_G1_MINI_ALU_ix437 (.Y (L1_1_L2_0_G1_MINI_ALU_nx436), .A0 (
         L1_1_L2_0_G1_MINI_ALU_nx507), .A1 (L1_1_L2_0_G1_MINI_ALU_nx511)) ;
    inv01 L1_1_L2_0_G1_MINI_ALU_ix510 (.Y (L1_1_L2_0_G1_MINI_ALU_nx509), .A (
          L1_1_L2_0_G1_MINI_ALU_BoothP_14)) ;
    xnor2 L1_1_L2_0_G1_MINI_ALU_ix512 (.Y (L1_1_L2_0_G1_MINI_ALU_nx511), .A0 (
          L1_1_L2_0_G1_MINI_ALU_BoothOperand_15), .A1 (
          L1_1_L2_0_G1_MINI_ALU_BoothP_15)) ;
    xnor2 L1_1_L2_0_G1_MINI_ALU_ix457 (.Y (L1_1_L2_0_G1_MINI_ALU_nx456), .A0 (
          L1_1_L2_0_G1_MINI_ALU_nx515), .A1 (L1_1_L2_0_G1_MINI_ALU_nx454)) ;
    inv01 L1_1_L2_0_G1_MINI_ALU_ix518 (.Y (L1_1_L2_0_G1_MINI_ALU_nx517), .A (
          L1_1_L2_0_G1_MINI_ALU_BoothP_15)) ;
    xor2 L1_1_L2_0_G1_MINI_ALU_ix455 (.Y (L1_1_L2_0_G1_MINI_ALU_nx454), .A0 (
         L1_1_L2_0_G1_MINI_ALU_BoothOperand_16), .A1 (
         L1_1_L2_0_G1_MINI_ALU_BoothP_16)) ;
    mux21_ni L1_1_L2_0_G1_MINI_ALU_ix91 (.Y (L1SecondOperands_5__0), .A0 (
             L1_1_L2_0_G1_MINI_ALU_BoothP_1), .A1 (WindowDin_1__0__0), .S0 (
             Instr)) ;
    mux21_ni L1_1_L2_0_G1_MINI_ALU_ix99 (.Y (L1SecondOperands_5__1), .A0 (
             L1_1_L2_0_G1_MINI_ALU_BoothP_2), .A1 (WindowDin_1__0__1), .S0 (
             Instr)) ;
    mux21_ni L1_1_L2_0_G1_MINI_ALU_ix107 (.Y (L1SecondOperands_5__2), .A0 (
             L1_1_L2_0_G1_MINI_ALU_BoothP_3), .A1 (WindowDin_1__0__2), .S0 (
             Instr)) ;
    mux21_ni L1_1_L2_0_G1_MINI_ALU_ix115 (.Y (L1SecondOperands_5__3), .A0 (
             L1_1_L2_0_G1_MINI_ALU_BoothP_4), .A1 (WindowDin_1__0__3), .S0 (
             Instr)) ;
    mux21_ni L1_1_L2_0_G1_MINI_ALU_ix123 (.Y (L1SecondOperands_5__4), .A0 (
             L1_1_L2_0_G1_MINI_ALU_BoothP_5), .A1 (WindowDin_1__0__4), .S0 (
             Instr)) ;
    mux21_ni L1_1_L2_0_G1_MINI_ALU_ix131 (.Y (L1SecondOperands_5__5), .A0 (
             L1_1_L2_0_G1_MINI_ALU_BoothP_6), .A1 (WindowDin_1__0__5), .S0 (
             Instr)) ;
    mux21_ni L1_1_L2_0_G1_MINI_ALU_ix139 (.Y (L1SecondOperands_5__6), .A0 (
             L1_1_L2_0_G1_MINI_ALU_BoothP_7), .A1 (WindowDin_1__0__6), .S0 (
             Instr)) ;
    mux21_ni L1_1_L2_0_G1_MINI_ALU_ix147 (.Y (L1SecondOperands_5__7), .A0 (
             L1_1_L2_0_G1_MINI_ALU_BoothP_8), .A1 (WindowDin_1__0__7), .S0 (
             Instr)) ;
    xor2 L1_1_L2_0_G1_MINI_ALU_ix77 (.Y (L1Results_5__1), .A0 (
         L1_1_L2_0_G1_MINI_ALU_nx529), .A1 (L1_1_L2_0_G1_MINI_ALU_nx531)) ;
    nand02 L1_1_L2_0_G1_MINI_ALU_ix530 (.Y (L1_1_L2_0_G1_MINI_ALU_nx529), .A0 (
           L1SecondOperands_5__0), .A1 (L1FirstOperands_5__0)) ;
    xnor2 L1_1_L2_0_G1_MINI_ALU_ix532 (.Y (L1_1_L2_0_G1_MINI_ALU_nx531), .A0 (
          L1SecondOperands_5__1), .A1 (L1FirstOperands_5__1)) ;
    xor2 L1_1_L2_0_G1_MINI_ALU_ix75 (.Y (L1Results_5__2), .A0 (
         L1_1_L2_0_G1_MINI_ALU_nx534), .A1 (L1_1_L2_0_G1_MINI_ALU_nx537)) ;
    aoi32 L1_1_L2_0_G1_MINI_ALU_ix535 (.Y (L1_1_L2_0_G1_MINI_ALU_nx534), .A0 (
          L1SecondOperands_5__0), .A1 (L1FirstOperands_5__0), .A2 (
          L1_1_L2_0_G1_MINI_ALU_nx30), .B0 (L1FirstOperands_5__1), .B1 (
          L1SecondOperands_5__1)) ;
    xnor2 L1_1_L2_0_G1_MINI_ALU_ix538 (.Y (L1_1_L2_0_G1_MINI_ALU_nx537), .A0 (
          L1SecondOperands_5__2), .A1 (L1FirstOperands_5__2)) ;
    xor2 L1_1_L2_0_G1_MINI_ALU_ix73 (.Y (L1Results_5__3), .A0 (
         L1_1_L2_0_G1_MINI_ALU_nx540), .A1 (L1_1_L2_0_G1_MINI_ALU_nx544)) ;
    aoi22 L1_1_L2_0_G1_MINI_ALU_ix541 (.Y (L1_1_L2_0_G1_MINI_ALU_nx540), .A0 (
          L1FirstOperands_5__2), .A1 (L1SecondOperands_5__2), .B0 (
          L1_1_L2_0_G1_MINI_ALU_nx40), .B1 (L1_1_L2_0_G1_MINI_ALU_nx24)) ;
    xnor2 L1_1_L2_0_G1_MINI_ALU_ix545 (.Y (L1_1_L2_0_G1_MINI_ALU_nx544), .A0 (
          L1SecondOperands_5__3), .A1 (L1FirstOperands_5__3)) ;
    xor2 L1_1_L2_0_G1_MINI_ALU_ix71 (.Y (L1Results_5__4), .A0 (
         L1_1_L2_0_G1_MINI_ALU_nx547), .A1 (L1_1_L2_0_G1_MINI_ALU_nx551)) ;
    aoi22 L1_1_L2_0_G1_MINI_ALU_ix548 (.Y (L1_1_L2_0_G1_MINI_ALU_nx547), .A0 (
          L1FirstOperands_5__3), .A1 (L1SecondOperands_5__3), .B0 (
          L1_1_L2_0_G1_MINI_ALU_nx44), .B1 (L1_1_L2_0_G1_MINI_ALU_nx18)) ;
    xnor2 L1_1_L2_0_G1_MINI_ALU_ix552 (.Y (L1_1_L2_0_G1_MINI_ALU_nx551), .A0 (
          L1SecondOperands_5__4), .A1 (L1FirstOperands_5__4)) ;
    xor2 L1_1_L2_0_G1_MINI_ALU_ix69 (.Y (L1Results_5__5), .A0 (
         L1_1_L2_0_G1_MINI_ALU_nx554), .A1 (L1_1_L2_0_G1_MINI_ALU_nx558)) ;
    aoi22 L1_1_L2_0_G1_MINI_ALU_ix555 (.Y (L1_1_L2_0_G1_MINI_ALU_nx554), .A0 (
          L1FirstOperands_5__4), .A1 (L1SecondOperands_5__4), .B0 (
          L1_1_L2_0_G1_MINI_ALU_nx48), .B1 (L1_1_L2_0_G1_MINI_ALU_nx12)) ;
    xnor2 L1_1_L2_0_G1_MINI_ALU_ix559 (.Y (L1_1_L2_0_G1_MINI_ALU_nx558), .A0 (
          L1SecondOperands_5__5), .A1 (L1FirstOperands_5__5)) ;
    xor2 L1_1_L2_0_G1_MINI_ALU_ix67 (.Y (L1Results_5__6), .A0 (
         L1_1_L2_0_G1_MINI_ALU_nx561), .A1 (L1_1_L2_0_G1_MINI_ALU_nx565)) ;
    aoi22 L1_1_L2_0_G1_MINI_ALU_ix562 (.Y (L1_1_L2_0_G1_MINI_ALU_nx561), .A0 (
          L1FirstOperands_5__5), .A1 (L1SecondOperands_5__5), .B0 (
          L1_1_L2_0_G1_MINI_ALU_nx52), .B1 (L1_1_L2_0_G1_MINI_ALU_nx6)) ;
    xnor2 L1_1_L2_0_G1_MINI_ALU_ix566 (.Y (L1_1_L2_0_G1_MINI_ALU_nx565), .A0 (
          L1SecondOperands_5__6), .A1 (L1FirstOperands_5__6)) ;
    xnor2 L1_1_L2_0_G1_MINI_ALU_ix65 (.Y (L1Results_5__7), .A0 (
          L1_1_L2_0_G1_MINI_ALU_nx568), .A1 (L1_1_L2_0_G1_MINI_ALU_nx62)) ;
    aoi22 L1_1_L2_0_G1_MINI_ALU_ix569 (.Y (L1_1_L2_0_G1_MINI_ALU_nx568), .A0 (
          L1FirstOperands_5__6), .A1 (L1SecondOperands_5__6), .B0 (
          L1_1_L2_0_G1_MINI_ALU_nx56), .B1 (L1_1_L2_0_G1_MINI_ALU_nx0)) ;
    xor2 L1_1_L2_0_G1_MINI_ALU_ix63 (.Y (L1_1_L2_0_G1_MINI_ALU_nx62), .A0 (
         L1SecondOperands_5__7), .A1 (L1FirstOperands_5__7)) ;
    inv01 L1_1_L2_0_G1_MINI_ALU_ix155 (.Y (L1_1_L2_0_G1_MINI_ALU_nx154), .A (
          L1_1_L2_0_G1_MINI_ALU_nx383)) ;
    inv01 L1_1_L2_0_G1_MINI_ALU_ix57 (.Y (L1_1_L2_0_G1_MINI_ALU_nx56), .A (
          L1_1_L2_0_G1_MINI_ALU_nx561)) ;
    inv01 L1_1_L2_0_G1_MINI_ALU_ix53 (.Y (L1_1_L2_0_G1_MINI_ALU_nx52), .A (
          L1_1_L2_0_G1_MINI_ALU_nx554)) ;
    inv01 L1_1_L2_0_G1_MINI_ALU_ix49 (.Y (L1_1_L2_0_G1_MINI_ALU_nx48), .A (
          L1_1_L2_0_G1_MINI_ALU_nx547)) ;
    inv01 L1_1_L2_0_G1_MINI_ALU_ix45 (.Y (L1_1_L2_0_G1_MINI_ALU_nx44), .A (
          L1_1_L2_0_G1_MINI_ALU_nx540)) ;
    inv01 L1_1_L2_0_G1_MINI_ALU_ix41 (.Y (L1_1_L2_0_G1_MINI_ALU_nx40), .A (
          L1_1_L2_0_G1_MINI_ALU_nx534)) ;
    inv01 L1_1_L2_0_G1_MINI_ALU_ix31 (.Y (L1_1_L2_0_G1_MINI_ALU_nx30), .A (
          L1_1_L2_0_G1_MINI_ALU_nx531)) ;
    inv01 L1_1_L2_0_G1_MINI_ALU_ix25 (.Y (L1_1_L2_0_G1_MINI_ALU_nx24), .A (
          L1_1_L2_0_G1_MINI_ALU_nx537)) ;
    inv01 L1_1_L2_0_G1_MINI_ALU_ix19 (.Y (L1_1_L2_0_G1_MINI_ALU_nx18), .A (
          L1_1_L2_0_G1_MINI_ALU_nx544)) ;
    inv01 L1_1_L2_0_G1_MINI_ALU_ix13 (.Y (L1_1_L2_0_G1_MINI_ALU_nx12), .A (
          L1_1_L2_0_G1_MINI_ALU_nx551)) ;
    inv01 L1_1_L2_0_G1_MINI_ALU_ix7 (.Y (L1_1_L2_0_G1_MINI_ALU_nx6), .A (
          L1_1_L2_0_G1_MINI_ALU_nx558)) ;
    inv01 L1_1_L2_0_G1_MINI_ALU_ix1 (.Y (L1_1_L2_0_G1_MINI_ALU_nx0), .A (
          L1_1_L2_0_G1_MINI_ALU_nx565)) ;
    fake_gnd L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix216 (.Y (
             L1_1_L2_0_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    nor02ii L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix81 (.Y (
            L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx80), .A0 (Instr), .A1 (Start)) ;
    aoi21 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix77 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_10), .A0 (
          FilterDin_1__0__1), .A1 (FilterDin_1__0__0), .B0 (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx4)) ;
    nor02_2x L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix5 (.Y (
             L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx4), .A0 (FilterDin_1__0__0), .A1 (
             FilterDin_1__0__1)) ;
    aoi21 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix67 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_11), .A0 (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx328), .A1 (FilterDin_1__0__2), .B0 (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx8)) ;
    nor03_2x L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix9 (.Y (
             L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx8), .A0 (FilterDin_1__0__2), .A1 (
             FilterDin_1__0__0), .A2 (FilterDin_1__0__1)) ;
    xnor2 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix59 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_12), .A0 (
          FilterDin_1__0__3), .A1 (L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx8)) ;
    xnor2 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix51 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_13), .A0 (
          FilterDin_1__0__4), .A1 (L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx12)) ;
    nor04 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix13 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx12), .A0 (FilterDin_1__0__3), .A1 (
          FilterDin_1__0__2), .A2 (FilterDin_1__0__0), .A3 (FilterDin_1__0__1)
          ) ;
    xnor2 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix43 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_14), .A0 (
          FilterDin_1__0__5), .A1 (L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx16)) ;
    nor02ii L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix17 (.Y (
            L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx16), .A0 (FilterDin_1__0__4), .A1 (
            L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx12)) ;
    xnor2 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix35 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_15), .A0 (
          FilterDin_1__0__6), .A1 (L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx20)) ;
    nor02ii L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix21 (.Y (
            L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx20), .A0 (FilterDin_1__0__5), .A1 (
            L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx16)) ;
    xnor2 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix27 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_16), .A0 (
          FilterDin_1__0__7), .A1 (L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx24)) ;
    nor02ii L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix25 (.Y (
            L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx24), .A0 (FilterDin_1__0__6), .A1 (
            L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx20)) ;
    inv01 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix329 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx328), .A (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx4)) ;
    inv02 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix383 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx384), .A (
          L1_1_L2_0_G1_MINI_ALU_BoothP_0)) ;
    dff L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_0 (.Q (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_0), .QB (\$dummy [259]), 
        .D (L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .CLK (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    nor02_2x L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix567 (.Y (
             L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566), .A0 (RST), .A1 (
             L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644)) ;
    dff L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_1 (.Q (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_1), .QB (\$dummy [260]), 
        .D (L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .CLK (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_2 (.Q (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_2), .QB (\$dummy [261]), 
        .D (L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .CLK (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_3 (.Q (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_3), .QB (\$dummy [262]), 
        .D (L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .CLK (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_4 (.Q (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_4), .QB (\$dummy [263]), 
        .D (L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .CLK (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_5 (.Q (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_5), .QB (\$dummy [264]), 
        .D (L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .CLK (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_6 (.Q (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_6), .QB (\$dummy [265]), 
        .D (L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .CLK (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_7 (.Q (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_7), .QB (\$dummy [266]), 
        .D (L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .CLK (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_8 (.Q (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_8), .QB (\$dummy [267]), 
        .D (L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .CLK (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_9 (.Q (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_9), .QB (\$dummy [268]), 
        .D (L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .CLK (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_10 (.Q (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_10), .QB (\$dummy [269])
        , .D (L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .CLK (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_11 (.Q (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_11), .QB (\$dummy [270])
        , .D (L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .CLK (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_12 (.Q (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_12), .QB (\$dummy [271])
        , .D (L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .CLK (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_13 (.Q (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_13), .QB (\$dummy [272])
        , .D (L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .CLK (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_14 (.Q (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_14), .QB (\$dummy [273])
        , .D (L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .CLK (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_15 (.Q (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_15), .QB (\$dummy [274])
        , .D (L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .CLK (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_16 (.Q (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_16), .QB (\$dummy [275])
        , .D (L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .CLK (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    inv02 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix623 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624), .A (CLK)) ;
    inv02 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix625 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626), .A (CLK)) ;
    inv02 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix627 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628), .A (CLK)) ;
    inv02 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix643 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644), .A (nx7818)) ;
    dff L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_0 (.Q (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_0), .QB (\$dummy [276]), 
        .D (L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .CLK (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    nor02_2x L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix567 (.Y (
             L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566), .A0 (RST), .A1 (
             L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644)) ;
    dff L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_1 (.Q (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_1), .QB (\$dummy [277]), 
        .D (L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .CLK (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_2 (.Q (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_2), .QB (\$dummy [278]), 
        .D (L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .CLK (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_3 (.Q (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_3), .QB (\$dummy [279]), 
        .D (L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .CLK (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_4 (.Q (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_4), .QB (\$dummy [280]), 
        .D (L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .CLK (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_5 (.Q (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_5), .QB (\$dummy [281]), 
        .D (L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .CLK (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_6 (.Q (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_6), .QB (\$dummy [282]), 
        .D (L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .CLK (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_7 (.Q (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_7), .QB (\$dummy [283]), 
        .D (L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .CLK (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_8 (.Q (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_8), .QB (\$dummy [284]), 
        .D (L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .CLK (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_9 (.Q (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_9), .QB (\$dummy [285]), 
        .D (L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .CLK (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_10 (.Q (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_10), .QB (\$dummy [286])
        , .D (L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .CLK (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_11 (.Q (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_11), .QB (\$dummy [287])
        , .D (L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .CLK (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_12 (.Q (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_12), .QB (\$dummy [288])
        , .D (L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .CLK (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_13 (.Q (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_13), .QB (\$dummy [289])
        , .D (L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .CLK (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_14 (.Q (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_14), .QB (\$dummy [290])
        , .D (L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .CLK (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_15 (.Q (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_15), .QB (\$dummy [291])
        , .D (L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .CLK (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_16 (.Q (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_16), .QB (\$dummy [292])
        , .D (L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .CLK (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    inv02 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix623 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624), .A (CLK)) ;
    inv02 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix625 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626), .A (CLK)) ;
    inv02 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix627 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628), .A (CLK)) ;
    inv02 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix643 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644), .A (nx7824)) ;
    dff L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_0 (.Q (
        L1_1_L2_0_G1_MINI_ALU_BoothP_0), .QB (\$dummy [293]), .D (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .CLK (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    nor02_2x L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix567 (.Y (
             L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566), .A0 (RST), .A1 (
             L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    dff L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_1 (.Q (
        L1_1_L2_0_G1_MINI_ALU_BoothP_1), .QB (\$dummy [294]), .D (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .CLK (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_2 (.Q (
        L1_1_L2_0_G1_MINI_ALU_BoothP_2), .QB (\$dummy [295]), .D (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .CLK (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_3 (.Q (
        L1_1_L2_0_G1_MINI_ALU_BoothP_3), .QB (\$dummy [296]), .D (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .CLK (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_4 (.Q (
        L1_1_L2_0_G1_MINI_ALU_BoothP_4), .QB (\$dummy [297]), .D (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .CLK (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_5 (.Q (
        L1_1_L2_0_G1_MINI_ALU_BoothP_5), .QB (\$dummy [298]), .D (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .CLK (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_6 (.Q (
        L1_1_L2_0_G1_MINI_ALU_BoothP_6), .QB (\$dummy [299]), .D (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .CLK (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_7 (.Q (
        L1_1_L2_0_G1_MINI_ALU_BoothP_7), .QB (\$dummy [300]), .D (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .CLK (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_8 (.Q (
        L1_1_L2_0_G1_MINI_ALU_BoothP_8), .QB (\$dummy [301]), .D (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .CLK (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_9 (.Q (
        L1_1_L2_0_G1_MINI_ALU_BoothP_9), .QB (\$dummy [302]), .D (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .CLK (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_10 (.Q (
        L1_1_L2_0_G1_MINI_ALU_BoothP_10), .QB (\$dummy [303]), .D (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .CLK (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_11 (.Q (
        L1_1_L2_0_G1_MINI_ALU_BoothP_11), .QB (\$dummy [304]), .D (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .CLK (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_12 (.Q (
        L1_1_L2_0_G1_MINI_ALU_BoothP_12), .QB (\$dummy [305]), .D (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .CLK (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_13 (.Q (
        L1_1_L2_0_G1_MINI_ALU_BoothP_13), .QB (\$dummy [306]), .D (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .CLK (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_14 (.Q (
        L1_1_L2_0_G1_MINI_ALU_BoothP_14), .QB (\$dummy [307]), .D (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .CLK (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_15 (.Q (
        L1_1_L2_0_G1_MINI_ALU_BoothP_15), .QB (\$dummy [308]), .D (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .CLK (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_16 (.Q (
        L1_1_L2_0_G1_MINI_ALU_BoothP_16), .QB (\$dummy [309]), .D (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .CLK (
        L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    inv02 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix623 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624), .A (CLK)) ;
    inv02 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix625 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626), .A (CLK)) ;
    inv02 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix627 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628), .A (CLK)) ;
    inv02 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix643 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644), .A (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642)) ;
    xor2 L1_1_L2_1_G1_MINI_ALU_ix83 (.Y (L1Results_6__0), .A0 (
         L1SecondOperands_6__0), .A1 (L1FirstOperands_6__0)) ;
    xnor2 L1_1_L2_1_G1_MINI_ALU_ix380 (.Y (L1_1_L2_1_G1_MINI_ALU_nx379), .A0 (
          L1_1_L2_1_G1_MINI_ALU_nx381), .A1 (L1_1_L2_1_G1_MINI_ALU_nx383)) ;
    nand02 L1_1_L2_1_G1_MINI_ALU_ix382 (.Y (L1_1_L2_1_G1_MINI_ALU_nx381), .A0 (
           L1_1_L2_1_G1_MINI_ALU_BoothOperand_0), .A1 (nx7844)) ;
    xnor2 L1_1_L2_1_G1_MINI_ALU_ix384 (.Y (L1_1_L2_1_G1_MINI_ALU_nx383), .A0 (
          L1_1_L2_1_G1_MINI_ALU_BoothOperand_1), .A1 (
          L1_1_L2_1_G1_MINI_ALU_BoothP_1)) ;
    inv01 L1_1_L2_1_G1_MINI_ALU_ix388 (.Y (L1_1_L2_1_G1_MINI_ALU_nx387), .A (
          L1_1_L2_1_G1_MINI_ALU_BoothP_2)) ;
    xnor2 L1_1_L2_1_G1_MINI_ALU_ix390 (.Y (L1_1_L2_1_G1_MINI_ALU_nx389), .A0 (
          L1_1_L2_1_G1_MINI_ALU_nx391), .A1 (L1_1_L2_1_G1_MINI_ALU_nx395)) ;
    aoi32 L1_1_L2_1_G1_MINI_ALU_ix392 (.Y (L1_1_L2_1_G1_MINI_ALU_nx391), .A0 (
          L1_1_L2_1_G1_MINI_ALU_BoothOperand_0), .A1 (nx7844), .A2 (
          L1_1_L2_1_G1_MINI_ALU_nx154), .B0 (L1_1_L2_1_G1_MINI_ALU_BoothP_1), .B1 (
          L1_1_L2_1_G1_MINI_ALU_BoothOperand_1)) ;
    xnor2 L1_1_L2_1_G1_MINI_ALU_ix396 (.Y (L1_1_L2_1_G1_MINI_ALU_nx395), .A0 (
          L1_1_L2_1_G1_MINI_ALU_BoothOperand_2), .A1 (
          L1_1_L2_1_G1_MINI_ALU_BoothP_2)) ;
    inv01 L1_1_L2_1_G1_MINI_ALU_ix400 (.Y (L1_1_L2_1_G1_MINI_ALU_nx399), .A (
          L1_1_L2_1_G1_MINI_ALU_BoothP_3)) ;
    xnor2 L1_1_L2_1_G1_MINI_ALU_ix402 (.Y (L1_1_L2_1_G1_MINI_ALU_nx401), .A0 (
          L1_1_L2_1_G1_MINI_ALU_nx403), .A1 (L1_1_L2_1_G1_MINI_ALU_nx405)) ;
    xnor2 L1_1_L2_1_G1_MINI_ALU_ix406 (.Y (L1_1_L2_1_G1_MINI_ALU_nx405), .A0 (
          L1_1_L2_1_G1_MINI_ALU_BoothOperand_3), .A1 (
          L1_1_L2_1_G1_MINI_ALU_BoothP_3)) ;
    inv01 L1_1_L2_1_G1_MINI_ALU_ix410 (.Y (L1_1_L2_1_G1_MINI_ALU_nx409), .A (
          L1_1_L2_1_G1_MINI_ALU_BoothP_4)) ;
    xnor2 L1_1_L2_1_G1_MINI_ALU_ix412 (.Y (L1_1_L2_1_G1_MINI_ALU_nx411), .A0 (
          L1_1_L2_1_G1_MINI_ALU_nx413), .A1 (L1_1_L2_1_G1_MINI_ALU_nx415)) ;
    xnor2 L1_1_L2_1_G1_MINI_ALU_ix416 (.Y (L1_1_L2_1_G1_MINI_ALU_nx415), .A0 (
          L1_1_L2_1_G1_MINI_ALU_BoothOperand_4), .A1 (
          L1_1_L2_1_G1_MINI_ALU_BoothP_4)) ;
    inv01 L1_1_L2_1_G1_MINI_ALU_ix420 (.Y (L1_1_L2_1_G1_MINI_ALU_nx419), .A (
          L1_1_L2_1_G1_MINI_ALU_BoothP_5)) ;
    xnor2 L1_1_L2_1_G1_MINI_ALU_ix422 (.Y (L1_1_L2_1_G1_MINI_ALU_nx421), .A0 (
          L1_1_L2_1_G1_MINI_ALU_nx423), .A1 (L1_1_L2_1_G1_MINI_ALU_nx425)) ;
    xnor2 L1_1_L2_1_G1_MINI_ALU_ix426 (.Y (L1_1_L2_1_G1_MINI_ALU_nx425), .A0 (
          L1_1_L2_1_G1_MINI_ALU_BoothOperand_5), .A1 (
          L1_1_L2_1_G1_MINI_ALU_BoothP_5)) ;
    inv01 L1_1_L2_1_G1_MINI_ALU_ix430 (.Y (L1_1_L2_1_G1_MINI_ALU_nx429), .A (
          L1_1_L2_1_G1_MINI_ALU_BoothP_6)) ;
    xnor2 L1_1_L2_1_G1_MINI_ALU_ix432 (.Y (L1_1_L2_1_G1_MINI_ALU_nx431), .A0 (
          L1_1_L2_1_G1_MINI_ALU_nx433), .A1 (L1_1_L2_1_G1_MINI_ALU_nx435)) ;
    xnor2 L1_1_L2_1_G1_MINI_ALU_ix436 (.Y (L1_1_L2_1_G1_MINI_ALU_nx435), .A0 (
          L1_1_L2_1_G1_MINI_ALU_BoothOperand_6), .A1 (
          L1_1_L2_1_G1_MINI_ALU_BoothP_6)) ;
    inv01 L1_1_L2_1_G1_MINI_ALU_ix440 (.Y (L1_1_L2_1_G1_MINI_ALU_nx439), .A (
          L1_1_L2_1_G1_MINI_ALU_BoothP_7)) ;
    xnor2 L1_1_L2_1_G1_MINI_ALU_ix442 (.Y (L1_1_L2_1_G1_MINI_ALU_nx441), .A0 (
          L1_1_L2_1_G1_MINI_ALU_nx443), .A1 (L1_1_L2_1_G1_MINI_ALU_nx445)) ;
    xnor2 L1_1_L2_1_G1_MINI_ALU_ix446 (.Y (L1_1_L2_1_G1_MINI_ALU_nx445), .A0 (
          L1_1_L2_1_G1_MINI_ALU_BoothOperand_7), .A1 (
          L1_1_L2_1_G1_MINI_ALU_BoothP_7)) ;
    inv01 L1_1_L2_1_G1_MINI_ALU_ix450 (.Y (L1_1_L2_1_G1_MINI_ALU_nx449), .A (
          L1_1_L2_1_G1_MINI_ALU_BoothP_8)) ;
    xnor2 L1_1_L2_1_G1_MINI_ALU_ix452 (.Y (L1_1_L2_1_G1_MINI_ALU_nx451), .A0 (
          L1_1_L2_1_G1_MINI_ALU_nx453), .A1 (L1_1_L2_1_G1_MINI_ALU_nx455)) ;
    xnor2 L1_1_L2_1_G1_MINI_ALU_ix456 (.Y (L1_1_L2_1_G1_MINI_ALU_nx455), .A0 (
          L1_1_L2_1_G1_MINI_ALU_BoothOperand_8), .A1 (
          L1_1_L2_1_G1_MINI_ALU_BoothP_8)) ;
    xor2 L1_1_L2_1_G1_MINI_ALU_ix317 (.Y (L1_1_L2_1_G1_MINI_ALU_nx316), .A0 (
         L1_1_L2_1_G1_MINI_ALU_nx461), .A1 (L1_1_L2_1_G1_MINI_ALU_nx463)) ;
    xnor2 L1_1_L2_1_G1_MINI_ALU_ix464 (.Y (L1_1_L2_1_G1_MINI_ALU_nx463), .A0 (
          L1_1_L2_1_G1_MINI_ALU_BoothOperand_9), .A1 (
          L1_1_L2_1_G1_MINI_ALU_BoothP_9)) ;
    xor2 L1_1_L2_1_G1_MINI_ALU_ix337 (.Y (L1_1_L2_1_G1_MINI_ALU_nx336), .A0 (
         L1_1_L2_1_G1_MINI_ALU_nx467), .A1 (L1_1_L2_1_G1_MINI_ALU_nx471)) ;
    inv01 L1_1_L2_1_G1_MINI_ALU_ix470 (.Y (L1_1_L2_1_G1_MINI_ALU_nx469), .A (
          L1_1_L2_1_G1_MINI_ALU_BoothP_9)) ;
    xnor2 L1_1_L2_1_G1_MINI_ALU_ix472 (.Y (L1_1_L2_1_G1_MINI_ALU_nx471), .A0 (
          L1_1_L2_1_G1_MINI_ALU_BoothOperand_10), .A1 (
          L1_1_L2_1_G1_MINI_ALU_BoothP_10)) ;
    xor2 L1_1_L2_1_G1_MINI_ALU_ix357 (.Y (L1_1_L2_1_G1_MINI_ALU_nx356), .A0 (
         L1_1_L2_1_G1_MINI_ALU_nx475), .A1 (L1_1_L2_1_G1_MINI_ALU_nx479)) ;
    inv01 L1_1_L2_1_G1_MINI_ALU_ix478 (.Y (L1_1_L2_1_G1_MINI_ALU_nx477), .A (
          L1_1_L2_1_G1_MINI_ALU_BoothP_10)) ;
    xnor2 L1_1_L2_1_G1_MINI_ALU_ix480 (.Y (L1_1_L2_1_G1_MINI_ALU_nx479), .A0 (
          L1_1_L2_1_G1_MINI_ALU_BoothOperand_11), .A1 (
          L1_1_L2_1_G1_MINI_ALU_BoothP_11)) ;
    xor2 L1_1_L2_1_G1_MINI_ALU_ix377 (.Y (L1_1_L2_1_G1_MINI_ALU_nx376), .A0 (
         L1_1_L2_1_G1_MINI_ALU_nx483), .A1 (L1_1_L2_1_G1_MINI_ALU_nx487)) ;
    inv01 L1_1_L2_1_G1_MINI_ALU_ix486 (.Y (L1_1_L2_1_G1_MINI_ALU_nx485), .A (
          L1_1_L2_1_G1_MINI_ALU_BoothP_11)) ;
    xnor2 L1_1_L2_1_G1_MINI_ALU_ix488 (.Y (L1_1_L2_1_G1_MINI_ALU_nx487), .A0 (
          L1_1_L2_1_G1_MINI_ALU_BoothOperand_12), .A1 (
          L1_1_L2_1_G1_MINI_ALU_BoothP_12)) ;
    xor2 L1_1_L2_1_G1_MINI_ALU_ix397 (.Y (L1_1_L2_1_G1_MINI_ALU_nx396), .A0 (
         L1_1_L2_1_G1_MINI_ALU_nx491), .A1 (L1_1_L2_1_G1_MINI_ALU_nx495)) ;
    inv01 L1_1_L2_1_G1_MINI_ALU_ix494 (.Y (L1_1_L2_1_G1_MINI_ALU_nx493), .A (
          L1_1_L2_1_G1_MINI_ALU_BoothP_12)) ;
    xnor2 L1_1_L2_1_G1_MINI_ALU_ix496 (.Y (L1_1_L2_1_G1_MINI_ALU_nx495), .A0 (
          L1_1_L2_1_G1_MINI_ALU_BoothOperand_13), .A1 (
          L1_1_L2_1_G1_MINI_ALU_BoothP_13)) ;
    xor2 L1_1_L2_1_G1_MINI_ALU_ix417 (.Y (L1_1_L2_1_G1_MINI_ALU_nx416), .A0 (
         L1_1_L2_1_G1_MINI_ALU_nx499), .A1 (L1_1_L2_1_G1_MINI_ALU_nx503)) ;
    inv01 L1_1_L2_1_G1_MINI_ALU_ix502 (.Y (L1_1_L2_1_G1_MINI_ALU_nx501), .A (
          L1_1_L2_1_G1_MINI_ALU_BoothP_13)) ;
    xnor2 L1_1_L2_1_G1_MINI_ALU_ix504 (.Y (L1_1_L2_1_G1_MINI_ALU_nx503), .A0 (
          L1_1_L2_1_G1_MINI_ALU_BoothOperand_14), .A1 (
          L1_1_L2_1_G1_MINI_ALU_BoothP_14)) ;
    xor2 L1_1_L2_1_G1_MINI_ALU_ix437 (.Y (L1_1_L2_1_G1_MINI_ALU_nx436), .A0 (
         L1_1_L2_1_G1_MINI_ALU_nx507), .A1 (L1_1_L2_1_G1_MINI_ALU_nx511)) ;
    inv01 L1_1_L2_1_G1_MINI_ALU_ix510 (.Y (L1_1_L2_1_G1_MINI_ALU_nx509), .A (
          L1_1_L2_1_G1_MINI_ALU_BoothP_14)) ;
    xnor2 L1_1_L2_1_G1_MINI_ALU_ix512 (.Y (L1_1_L2_1_G1_MINI_ALU_nx511), .A0 (
          L1_1_L2_1_G1_MINI_ALU_BoothOperand_15), .A1 (
          L1_1_L2_1_G1_MINI_ALU_BoothP_15)) ;
    xnor2 L1_1_L2_1_G1_MINI_ALU_ix457 (.Y (L1_1_L2_1_G1_MINI_ALU_nx456), .A0 (
          L1_1_L2_1_G1_MINI_ALU_nx515), .A1 (L1_1_L2_1_G1_MINI_ALU_nx454)) ;
    inv01 L1_1_L2_1_G1_MINI_ALU_ix518 (.Y (L1_1_L2_1_G1_MINI_ALU_nx517), .A (
          L1_1_L2_1_G1_MINI_ALU_BoothP_15)) ;
    xor2 L1_1_L2_1_G1_MINI_ALU_ix455 (.Y (L1_1_L2_1_G1_MINI_ALU_nx454), .A0 (
         L1_1_L2_1_G1_MINI_ALU_BoothOperand_16), .A1 (
         L1_1_L2_1_G1_MINI_ALU_BoothP_16)) ;
    mux21_ni L1_1_L2_1_G1_MINI_ALU_ix91 (.Y (L1SecondOperands_6__0), .A0 (
             L1_1_L2_1_G1_MINI_ALU_BoothP_1), .A1 (WindowDin_1__1__0), .S0 (
             Instr)) ;
    mux21_ni L1_1_L2_1_G1_MINI_ALU_ix99 (.Y (L1SecondOperands_6__1), .A0 (
             L1_1_L2_1_G1_MINI_ALU_BoothP_2), .A1 (WindowDin_1__1__1), .S0 (
             Instr)) ;
    mux21_ni L1_1_L2_1_G1_MINI_ALU_ix107 (.Y (L1SecondOperands_6__2), .A0 (
             L1_1_L2_1_G1_MINI_ALU_BoothP_3), .A1 (WindowDin_1__1__2), .S0 (
             Instr)) ;
    mux21_ni L1_1_L2_1_G1_MINI_ALU_ix115 (.Y (L1SecondOperands_6__3), .A0 (
             L1_1_L2_1_G1_MINI_ALU_BoothP_4), .A1 (WindowDin_1__1__3), .S0 (
             Instr)) ;
    mux21_ni L1_1_L2_1_G1_MINI_ALU_ix123 (.Y (L1SecondOperands_6__4), .A0 (
             L1_1_L2_1_G1_MINI_ALU_BoothP_5), .A1 (WindowDin_1__1__4), .S0 (
             Instr)) ;
    mux21_ni L1_1_L2_1_G1_MINI_ALU_ix131 (.Y (L1SecondOperands_6__5), .A0 (
             L1_1_L2_1_G1_MINI_ALU_BoothP_6), .A1 (WindowDin_1__1__5), .S0 (
             Instr)) ;
    mux21_ni L1_1_L2_1_G1_MINI_ALU_ix139 (.Y (L1SecondOperands_6__6), .A0 (
             L1_1_L2_1_G1_MINI_ALU_BoothP_7), .A1 (WindowDin_1__1__6), .S0 (
             Instr)) ;
    mux21_ni L1_1_L2_1_G1_MINI_ALU_ix147 (.Y (L1SecondOperands_6__7), .A0 (
             L1_1_L2_1_G1_MINI_ALU_BoothP_8), .A1 (WindowDin_1__1__7), .S0 (
             Instr)) ;
    xor2 L1_1_L2_1_G1_MINI_ALU_ix77 (.Y (L1Results_6__1), .A0 (
         L1_1_L2_1_G1_MINI_ALU_nx529), .A1 (L1_1_L2_1_G1_MINI_ALU_nx531)) ;
    nand02 L1_1_L2_1_G1_MINI_ALU_ix530 (.Y (L1_1_L2_1_G1_MINI_ALU_nx529), .A0 (
           L1SecondOperands_6__0), .A1 (L1FirstOperands_6__0)) ;
    xnor2 L1_1_L2_1_G1_MINI_ALU_ix532 (.Y (L1_1_L2_1_G1_MINI_ALU_nx531), .A0 (
          L1SecondOperands_6__1), .A1 (L1FirstOperands_6__1)) ;
    xor2 L1_1_L2_1_G1_MINI_ALU_ix75 (.Y (L1Results_6__2), .A0 (
         L1_1_L2_1_G1_MINI_ALU_nx534), .A1 (L1_1_L2_1_G1_MINI_ALU_nx537)) ;
    aoi32 L1_1_L2_1_G1_MINI_ALU_ix535 (.Y (L1_1_L2_1_G1_MINI_ALU_nx534), .A0 (
          L1SecondOperands_6__0), .A1 (L1FirstOperands_6__0), .A2 (
          L1_1_L2_1_G1_MINI_ALU_nx30), .B0 (L1FirstOperands_6__1), .B1 (
          L1SecondOperands_6__1)) ;
    xnor2 L1_1_L2_1_G1_MINI_ALU_ix538 (.Y (L1_1_L2_1_G1_MINI_ALU_nx537), .A0 (
          L1SecondOperands_6__2), .A1 (L1FirstOperands_6__2)) ;
    xor2 L1_1_L2_1_G1_MINI_ALU_ix73 (.Y (L1Results_6__3), .A0 (
         L1_1_L2_1_G1_MINI_ALU_nx540), .A1 (L1_1_L2_1_G1_MINI_ALU_nx544)) ;
    aoi22 L1_1_L2_1_G1_MINI_ALU_ix541 (.Y (L1_1_L2_1_G1_MINI_ALU_nx540), .A0 (
          L1FirstOperands_6__2), .A1 (L1SecondOperands_6__2), .B0 (
          L1_1_L2_1_G1_MINI_ALU_nx40), .B1 (L1_1_L2_1_G1_MINI_ALU_nx24)) ;
    xnor2 L1_1_L2_1_G1_MINI_ALU_ix545 (.Y (L1_1_L2_1_G1_MINI_ALU_nx544), .A0 (
          L1SecondOperands_6__3), .A1 (L1FirstOperands_6__3)) ;
    xor2 L1_1_L2_1_G1_MINI_ALU_ix71 (.Y (L1Results_6__4), .A0 (
         L1_1_L2_1_G1_MINI_ALU_nx547), .A1 (L1_1_L2_1_G1_MINI_ALU_nx551)) ;
    aoi22 L1_1_L2_1_G1_MINI_ALU_ix548 (.Y (L1_1_L2_1_G1_MINI_ALU_nx547), .A0 (
          L1FirstOperands_6__3), .A1 (L1SecondOperands_6__3), .B0 (
          L1_1_L2_1_G1_MINI_ALU_nx44), .B1 (L1_1_L2_1_G1_MINI_ALU_nx18)) ;
    xnor2 L1_1_L2_1_G1_MINI_ALU_ix552 (.Y (L1_1_L2_1_G1_MINI_ALU_nx551), .A0 (
          L1SecondOperands_6__4), .A1 (L1FirstOperands_6__4)) ;
    xor2 L1_1_L2_1_G1_MINI_ALU_ix69 (.Y (L1Results_6__5), .A0 (
         L1_1_L2_1_G1_MINI_ALU_nx554), .A1 (L1_1_L2_1_G1_MINI_ALU_nx558)) ;
    aoi22 L1_1_L2_1_G1_MINI_ALU_ix555 (.Y (L1_1_L2_1_G1_MINI_ALU_nx554), .A0 (
          L1FirstOperands_6__4), .A1 (L1SecondOperands_6__4), .B0 (
          L1_1_L2_1_G1_MINI_ALU_nx48), .B1 (L1_1_L2_1_G1_MINI_ALU_nx12)) ;
    xnor2 L1_1_L2_1_G1_MINI_ALU_ix559 (.Y (L1_1_L2_1_G1_MINI_ALU_nx558), .A0 (
          L1SecondOperands_6__5), .A1 (L1FirstOperands_6__5)) ;
    xor2 L1_1_L2_1_G1_MINI_ALU_ix67 (.Y (L1Results_6__6), .A0 (
         L1_1_L2_1_G1_MINI_ALU_nx561), .A1 (L1_1_L2_1_G1_MINI_ALU_nx565)) ;
    aoi22 L1_1_L2_1_G1_MINI_ALU_ix562 (.Y (L1_1_L2_1_G1_MINI_ALU_nx561), .A0 (
          L1FirstOperands_6__5), .A1 (L1SecondOperands_6__5), .B0 (
          L1_1_L2_1_G1_MINI_ALU_nx52), .B1 (L1_1_L2_1_G1_MINI_ALU_nx6)) ;
    xnor2 L1_1_L2_1_G1_MINI_ALU_ix566 (.Y (L1_1_L2_1_G1_MINI_ALU_nx565), .A0 (
          L1SecondOperands_6__6), .A1 (L1FirstOperands_6__6)) ;
    xnor2 L1_1_L2_1_G1_MINI_ALU_ix65 (.Y (L1Results_6__7), .A0 (
          L1_1_L2_1_G1_MINI_ALU_nx568), .A1 (L1_1_L2_1_G1_MINI_ALU_nx62)) ;
    aoi22 L1_1_L2_1_G1_MINI_ALU_ix569 (.Y (L1_1_L2_1_G1_MINI_ALU_nx568), .A0 (
          L1FirstOperands_6__6), .A1 (L1SecondOperands_6__6), .B0 (
          L1_1_L2_1_G1_MINI_ALU_nx56), .B1 (L1_1_L2_1_G1_MINI_ALU_nx0)) ;
    xor2 L1_1_L2_1_G1_MINI_ALU_ix63 (.Y (L1_1_L2_1_G1_MINI_ALU_nx62), .A0 (
         L1SecondOperands_6__7), .A1 (L1FirstOperands_6__7)) ;
    inv01 L1_1_L2_1_G1_MINI_ALU_ix155 (.Y (L1_1_L2_1_G1_MINI_ALU_nx154), .A (
          L1_1_L2_1_G1_MINI_ALU_nx383)) ;
    inv01 L1_1_L2_1_G1_MINI_ALU_ix57 (.Y (L1_1_L2_1_G1_MINI_ALU_nx56), .A (
          L1_1_L2_1_G1_MINI_ALU_nx561)) ;
    inv01 L1_1_L2_1_G1_MINI_ALU_ix53 (.Y (L1_1_L2_1_G1_MINI_ALU_nx52), .A (
          L1_1_L2_1_G1_MINI_ALU_nx554)) ;
    inv01 L1_1_L2_1_G1_MINI_ALU_ix49 (.Y (L1_1_L2_1_G1_MINI_ALU_nx48), .A (
          L1_1_L2_1_G1_MINI_ALU_nx547)) ;
    inv01 L1_1_L2_1_G1_MINI_ALU_ix45 (.Y (L1_1_L2_1_G1_MINI_ALU_nx44), .A (
          L1_1_L2_1_G1_MINI_ALU_nx540)) ;
    inv01 L1_1_L2_1_G1_MINI_ALU_ix41 (.Y (L1_1_L2_1_G1_MINI_ALU_nx40), .A (
          L1_1_L2_1_G1_MINI_ALU_nx534)) ;
    inv01 L1_1_L2_1_G1_MINI_ALU_ix31 (.Y (L1_1_L2_1_G1_MINI_ALU_nx30), .A (
          L1_1_L2_1_G1_MINI_ALU_nx531)) ;
    inv01 L1_1_L2_1_G1_MINI_ALU_ix25 (.Y (L1_1_L2_1_G1_MINI_ALU_nx24), .A (
          L1_1_L2_1_G1_MINI_ALU_nx537)) ;
    inv01 L1_1_L2_1_G1_MINI_ALU_ix19 (.Y (L1_1_L2_1_G1_MINI_ALU_nx18), .A (
          L1_1_L2_1_G1_MINI_ALU_nx544)) ;
    inv01 L1_1_L2_1_G1_MINI_ALU_ix13 (.Y (L1_1_L2_1_G1_MINI_ALU_nx12), .A (
          L1_1_L2_1_G1_MINI_ALU_nx551)) ;
    inv01 L1_1_L2_1_G1_MINI_ALU_ix7 (.Y (L1_1_L2_1_G1_MINI_ALU_nx6), .A (
          L1_1_L2_1_G1_MINI_ALU_nx558)) ;
    inv01 L1_1_L2_1_G1_MINI_ALU_ix1 (.Y (L1_1_L2_1_G1_MINI_ALU_nx0), .A (
          L1_1_L2_1_G1_MINI_ALU_nx565)) ;
    fake_gnd L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix216 (.Y (
             L1_1_L2_1_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    nor02ii L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix81 (.Y (
            L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx80), .A0 (Instr), .A1 (Start)) ;
    aoi21 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix77 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_10), .A0 (
          FilterDin_1__1__1), .A1 (FilterDin_1__1__0), .B0 (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx4)) ;
    nor02_2x L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix5 (.Y (
             L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx4), .A0 (FilterDin_1__1__0), .A1 (
             FilterDin_1__1__1)) ;
    aoi21 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix67 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_11), .A0 (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx328), .A1 (FilterDin_1__1__2), .B0 (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx8)) ;
    nor03_2x L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix9 (.Y (
             L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx8), .A0 (FilterDin_1__1__2), .A1 (
             FilterDin_1__1__0), .A2 (FilterDin_1__1__1)) ;
    xnor2 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix59 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_12), .A0 (
          FilterDin_1__1__3), .A1 (L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx8)) ;
    xnor2 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix51 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_13), .A0 (
          FilterDin_1__1__4), .A1 (L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx12)) ;
    nor04 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix13 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx12), .A0 (FilterDin_1__1__3), .A1 (
          FilterDin_1__1__2), .A2 (FilterDin_1__1__0), .A3 (FilterDin_1__1__1)
          ) ;
    xnor2 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix43 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_14), .A0 (
          FilterDin_1__1__5), .A1 (L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx16)) ;
    nor02ii L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix17 (.Y (
            L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx16), .A0 (FilterDin_1__1__4), .A1 (
            L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx12)) ;
    xnor2 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix35 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_15), .A0 (
          FilterDin_1__1__6), .A1 (L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx20)) ;
    nor02ii L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix21 (.Y (
            L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx20), .A0 (FilterDin_1__1__5), .A1 (
            L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx16)) ;
    xnor2 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix27 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_16), .A0 (
          FilterDin_1__1__7), .A1 (L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx24)) ;
    nor02ii L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix25 (.Y (
            L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx24), .A0 (FilterDin_1__1__6), .A1 (
            L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx20)) ;
    inv01 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix329 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx328), .A (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx4)) ;
    inv02 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix383 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx384), .A (
          L1_1_L2_1_G1_MINI_ALU_BoothP_0)) ;
    dff L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_0 (.Q (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_0), .QB (\$dummy [310]), 
        .D (L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .CLK (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    nor02_2x L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix567 (.Y (
             L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566), .A0 (RST), .A1 (
             L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644)) ;
    dff L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_1 (.Q (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_1), .QB (\$dummy [311]), 
        .D (L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .CLK (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_2 (.Q (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_2), .QB (\$dummy [312]), 
        .D (L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .CLK (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_3 (.Q (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_3), .QB (\$dummy [313]), 
        .D (L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .CLK (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_4 (.Q (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_4), .QB (\$dummy [314]), 
        .D (L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .CLK (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_5 (.Q (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_5), .QB (\$dummy [315]), 
        .D (L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .CLK (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_6 (.Q (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_6), .QB (\$dummy [316]), 
        .D (L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .CLK (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_7 (.Q (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_7), .QB (\$dummy [317]), 
        .D (L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .CLK (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_8 (.Q (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_8), .QB (\$dummy [318]), 
        .D (L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .CLK (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_9 (.Q (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_9), .QB (\$dummy [319]), 
        .D (L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .CLK (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_10 (.Q (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_10), .QB (\$dummy [320])
        , .D (L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .CLK (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_11 (.Q (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_11), .QB (\$dummy [321])
        , .D (L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .CLK (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_12 (.Q (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_12), .QB (\$dummy [322])
        , .D (L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .CLK (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_13 (.Q (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_13), .QB (\$dummy [323])
        , .D (L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .CLK (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_14 (.Q (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_14), .QB (\$dummy [324])
        , .D (L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .CLK (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_15 (.Q (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_15), .QB (\$dummy [325])
        , .D (L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .CLK (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_16 (.Q (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_16), .QB (\$dummy [326])
        , .D (L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .CLK (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    inv02 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix623 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624), .A (CLK)) ;
    inv02 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix625 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626), .A (CLK)) ;
    inv02 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix627 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628), .A (CLK)) ;
    inv02 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix643 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644), .A (nx7858)) ;
    dff L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_0 (.Q (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_0), .QB (\$dummy [327]), 
        .D (L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .CLK (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    nor02_2x L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix567 (.Y (
             L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566), .A0 (RST), .A1 (
             L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644)) ;
    dff L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_1 (.Q (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_1), .QB (\$dummy [328]), 
        .D (L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .CLK (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_2 (.Q (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_2), .QB (\$dummy [329]), 
        .D (L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .CLK (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_3 (.Q (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_3), .QB (\$dummy [330]), 
        .D (L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .CLK (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_4 (.Q (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_4), .QB (\$dummy [331]), 
        .D (L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .CLK (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_5 (.Q (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_5), .QB (\$dummy [332]), 
        .D (L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .CLK (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_6 (.Q (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_6), .QB (\$dummy [333]), 
        .D (L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .CLK (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_7 (.Q (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_7), .QB (\$dummy [334]), 
        .D (L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .CLK (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_8 (.Q (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_8), .QB (\$dummy [335]), 
        .D (L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .CLK (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_9 (.Q (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_9), .QB (\$dummy [336]), 
        .D (L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .CLK (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_10 (.Q (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_10), .QB (\$dummy [337])
        , .D (L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .CLK (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_11 (.Q (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_11), .QB (\$dummy [338])
        , .D (L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .CLK (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_12 (.Q (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_12), .QB (\$dummy [339])
        , .D (L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .CLK (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_13 (.Q (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_13), .QB (\$dummy [340])
        , .D (L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .CLK (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_14 (.Q (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_14), .QB (\$dummy [341])
        , .D (L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .CLK (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_15 (.Q (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_15), .QB (\$dummy [342])
        , .D (L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .CLK (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_16 (.Q (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_16), .QB (\$dummy [343])
        , .D (L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .CLK (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    inv02 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix623 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624), .A (CLK)) ;
    inv02 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix625 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626), .A (CLK)) ;
    inv02 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix627 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628), .A (CLK)) ;
    inv02 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix643 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644), .A (nx7864)) ;
    dff L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_0 (.Q (
        L1_1_L2_1_G1_MINI_ALU_BoothP_0), .QB (\$dummy [344]), .D (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .CLK (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    nor02_2x L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix567 (.Y (
             L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566), .A0 (RST), .A1 (
             L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    dff L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_1 (.Q (
        L1_1_L2_1_G1_MINI_ALU_BoothP_1), .QB (\$dummy [345]), .D (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .CLK (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_2 (.Q (
        L1_1_L2_1_G1_MINI_ALU_BoothP_2), .QB (\$dummy [346]), .D (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .CLK (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_3 (.Q (
        L1_1_L2_1_G1_MINI_ALU_BoothP_3), .QB (\$dummy [347]), .D (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .CLK (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_4 (.Q (
        L1_1_L2_1_G1_MINI_ALU_BoothP_4), .QB (\$dummy [348]), .D (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .CLK (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_5 (.Q (
        L1_1_L2_1_G1_MINI_ALU_BoothP_5), .QB (\$dummy [349]), .D (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .CLK (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_6 (.Q (
        L1_1_L2_1_G1_MINI_ALU_BoothP_6), .QB (\$dummy [350]), .D (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .CLK (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_7 (.Q (
        L1_1_L2_1_G1_MINI_ALU_BoothP_7), .QB (\$dummy [351]), .D (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .CLK (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_8 (.Q (
        L1_1_L2_1_G1_MINI_ALU_BoothP_8), .QB (\$dummy [352]), .D (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .CLK (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_9 (.Q (
        L1_1_L2_1_G1_MINI_ALU_BoothP_9), .QB (\$dummy [353]), .D (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .CLK (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_10 (.Q (
        L1_1_L2_1_G1_MINI_ALU_BoothP_10), .QB (\$dummy [354]), .D (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .CLK (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_11 (.Q (
        L1_1_L2_1_G1_MINI_ALU_BoothP_11), .QB (\$dummy [355]), .D (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .CLK (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_12 (.Q (
        L1_1_L2_1_G1_MINI_ALU_BoothP_12), .QB (\$dummy [356]), .D (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .CLK (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_13 (.Q (
        L1_1_L2_1_G1_MINI_ALU_BoothP_13), .QB (\$dummy [357]), .D (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .CLK (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_14 (.Q (
        L1_1_L2_1_G1_MINI_ALU_BoothP_14), .QB (\$dummy [358]), .D (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .CLK (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_15 (.Q (
        L1_1_L2_1_G1_MINI_ALU_BoothP_15), .QB (\$dummy [359]), .D (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .CLK (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_16 (.Q (
        L1_1_L2_1_G1_MINI_ALU_BoothP_16), .QB (\$dummy [360]), .D (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .CLK (
        L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    inv02 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix623 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624), .A (CLK)) ;
    inv02 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix625 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626), .A (CLK)) ;
    inv02 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix627 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628), .A (CLK)) ;
    inv02 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix643 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644), .A (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642)) ;
    xor2 L1_1_L2_2_G1_MINI_ALU_ix83 (.Y (L1Results_7__0), .A0 (
         L1SecondOperands_7__0), .A1 (L1FirstOperands_7__0)) ;
    xnor2 L1_1_L2_2_G1_MINI_ALU_ix380 (.Y (L1_1_L2_2_G1_MINI_ALU_nx379), .A0 (
          L1_1_L2_2_G1_MINI_ALU_nx381), .A1 (L1_1_L2_2_G1_MINI_ALU_nx383)) ;
    nand02 L1_1_L2_2_G1_MINI_ALU_ix382 (.Y (L1_1_L2_2_G1_MINI_ALU_nx381), .A0 (
           L1_1_L2_2_G1_MINI_ALU_BoothOperand_0), .A1 (nx7884)) ;
    xnor2 L1_1_L2_2_G1_MINI_ALU_ix384 (.Y (L1_1_L2_2_G1_MINI_ALU_nx383), .A0 (
          L1_1_L2_2_G1_MINI_ALU_BoothOperand_1), .A1 (
          L1_1_L2_2_G1_MINI_ALU_BoothP_1)) ;
    inv01 L1_1_L2_2_G1_MINI_ALU_ix388 (.Y (L1_1_L2_2_G1_MINI_ALU_nx387), .A (
          L1_1_L2_2_G1_MINI_ALU_BoothP_2)) ;
    xnor2 L1_1_L2_2_G1_MINI_ALU_ix390 (.Y (L1_1_L2_2_G1_MINI_ALU_nx389), .A0 (
          L1_1_L2_2_G1_MINI_ALU_nx391), .A1 (L1_1_L2_2_G1_MINI_ALU_nx395)) ;
    aoi32 L1_1_L2_2_G1_MINI_ALU_ix392 (.Y (L1_1_L2_2_G1_MINI_ALU_nx391), .A0 (
          L1_1_L2_2_G1_MINI_ALU_BoothOperand_0), .A1 (nx7884), .A2 (
          L1_1_L2_2_G1_MINI_ALU_nx154), .B0 (L1_1_L2_2_G1_MINI_ALU_BoothP_1), .B1 (
          L1_1_L2_2_G1_MINI_ALU_BoothOperand_1)) ;
    xnor2 L1_1_L2_2_G1_MINI_ALU_ix396 (.Y (L1_1_L2_2_G1_MINI_ALU_nx395), .A0 (
          L1_1_L2_2_G1_MINI_ALU_BoothOperand_2), .A1 (
          L1_1_L2_2_G1_MINI_ALU_BoothP_2)) ;
    inv01 L1_1_L2_2_G1_MINI_ALU_ix400 (.Y (L1_1_L2_2_G1_MINI_ALU_nx399), .A (
          L1_1_L2_2_G1_MINI_ALU_BoothP_3)) ;
    xnor2 L1_1_L2_2_G1_MINI_ALU_ix402 (.Y (L1_1_L2_2_G1_MINI_ALU_nx401), .A0 (
          L1_1_L2_2_G1_MINI_ALU_nx403), .A1 (L1_1_L2_2_G1_MINI_ALU_nx405)) ;
    xnor2 L1_1_L2_2_G1_MINI_ALU_ix406 (.Y (L1_1_L2_2_G1_MINI_ALU_nx405), .A0 (
          L1_1_L2_2_G1_MINI_ALU_BoothOperand_3), .A1 (
          L1_1_L2_2_G1_MINI_ALU_BoothP_3)) ;
    inv01 L1_1_L2_2_G1_MINI_ALU_ix410 (.Y (L1_1_L2_2_G1_MINI_ALU_nx409), .A (
          L1_1_L2_2_G1_MINI_ALU_BoothP_4)) ;
    xnor2 L1_1_L2_2_G1_MINI_ALU_ix412 (.Y (L1_1_L2_2_G1_MINI_ALU_nx411), .A0 (
          L1_1_L2_2_G1_MINI_ALU_nx413), .A1 (L1_1_L2_2_G1_MINI_ALU_nx415)) ;
    xnor2 L1_1_L2_2_G1_MINI_ALU_ix416 (.Y (L1_1_L2_2_G1_MINI_ALU_nx415), .A0 (
          L1_1_L2_2_G1_MINI_ALU_BoothOperand_4), .A1 (
          L1_1_L2_2_G1_MINI_ALU_BoothP_4)) ;
    inv01 L1_1_L2_2_G1_MINI_ALU_ix420 (.Y (L1_1_L2_2_G1_MINI_ALU_nx419), .A (
          L1_1_L2_2_G1_MINI_ALU_BoothP_5)) ;
    xnor2 L1_1_L2_2_G1_MINI_ALU_ix422 (.Y (L1_1_L2_2_G1_MINI_ALU_nx421), .A0 (
          L1_1_L2_2_G1_MINI_ALU_nx423), .A1 (L1_1_L2_2_G1_MINI_ALU_nx425)) ;
    xnor2 L1_1_L2_2_G1_MINI_ALU_ix426 (.Y (L1_1_L2_2_G1_MINI_ALU_nx425), .A0 (
          L1_1_L2_2_G1_MINI_ALU_BoothOperand_5), .A1 (
          L1_1_L2_2_G1_MINI_ALU_BoothP_5)) ;
    inv01 L1_1_L2_2_G1_MINI_ALU_ix430 (.Y (L1_1_L2_2_G1_MINI_ALU_nx429), .A (
          L1_1_L2_2_G1_MINI_ALU_BoothP_6)) ;
    xnor2 L1_1_L2_2_G1_MINI_ALU_ix432 (.Y (L1_1_L2_2_G1_MINI_ALU_nx431), .A0 (
          L1_1_L2_2_G1_MINI_ALU_nx433), .A1 (L1_1_L2_2_G1_MINI_ALU_nx435)) ;
    xnor2 L1_1_L2_2_G1_MINI_ALU_ix436 (.Y (L1_1_L2_2_G1_MINI_ALU_nx435), .A0 (
          L1_1_L2_2_G1_MINI_ALU_BoothOperand_6), .A1 (
          L1_1_L2_2_G1_MINI_ALU_BoothP_6)) ;
    inv01 L1_1_L2_2_G1_MINI_ALU_ix440 (.Y (L1_1_L2_2_G1_MINI_ALU_nx439), .A (
          L1_1_L2_2_G1_MINI_ALU_BoothP_7)) ;
    xnor2 L1_1_L2_2_G1_MINI_ALU_ix442 (.Y (L1_1_L2_2_G1_MINI_ALU_nx441), .A0 (
          L1_1_L2_2_G1_MINI_ALU_nx443), .A1 (L1_1_L2_2_G1_MINI_ALU_nx445)) ;
    xnor2 L1_1_L2_2_G1_MINI_ALU_ix446 (.Y (L1_1_L2_2_G1_MINI_ALU_nx445), .A0 (
          L1_1_L2_2_G1_MINI_ALU_BoothOperand_7), .A1 (
          L1_1_L2_2_G1_MINI_ALU_BoothP_7)) ;
    inv01 L1_1_L2_2_G1_MINI_ALU_ix450 (.Y (L1_1_L2_2_G1_MINI_ALU_nx449), .A (
          L1_1_L2_2_G1_MINI_ALU_BoothP_8)) ;
    xnor2 L1_1_L2_2_G1_MINI_ALU_ix452 (.Y (L1_1_L2_2_G1_MINI_ALU_nx451), .A0 (
          L1_1_L2_2_G1_MINI_ALU_nx453), .A1 (L1_1_L2_2_G1_MINI_ALU_nx455)) ;
    xnor2 L1_1_L2_2_G1_MINI_ALU_ix456 (.Y (L1_1_L2_2_G1_MINI_ALU_nx455), .A0 (
          L1_1_L2_2_G1_MINI_ALU_BoothOperand_8), .A1 (
          L1_1_L2_2_G1_MINI_ALU_BoothP_8)) ;
    xor2 L1_1_L2_2_G1_MINI_ALU_ix317 (.Y (L1_1_L2_2_G1_MINI_ALU_nx316), .A0 (
         L1_1_L2_2_G1_MINI_ALU_nx461), .A1 (L1_1_L2_2_G1_MINI_ALU_nx463)) ;
    xnor2 L1_1_L2_2_G1_MINI_ALU_ix464 (.Y (L1_1_L2_2_G1_MINI_ALU_nx463), .A0 (
          L1_1_L2_2_G1_MINI_ALU_BoothOperand_9), .A1 (
          L1_1_L2_2_G1_MINI_ALU_BoothP_9)) ;
    xor2 L1_1_L2_2_G1_MINI_ALU_ix337 (.Y (L1_1_L2_2_G1_MINI_ALU_nx336), .A0 (
         L1_1_L2_2_G1_MINI_ALU_nx467), .A1 (L1_1_L2_2_G1_MINI_ALU_nx471)) ;
    inv01 L1_1_L2_2_G1_MINI_ALU_ix470 (.Y (L1_1_L2_2_G1_MINI_ALU_nx469), .A (
          L1_1_L2_2_G1_MINI_ALU_BoothP_9)) ;
    xnor2 L1_1_L2_2_G1_MINI_ALU_ix472 (.Y (L1_1_L2_2_G1_MINI_ALU_nx471), .A0 (
          L1_1_L2_2_G1_MINI_ALU_BoothOperand_10), .A1 (
          L1_1_L2_2_G1_MINI_ALU_BoothP_10)) ;
    xor2 L1_1_L2_2_G1_MINI_ALU_ix357 (.Y (L1_1_L2_2_G1_MINI_ALU_nx356), .A0 (
         L1_1_L2_2_G1_MINI_ALU_nx475), .A1 (L1_1_L2_2_G1_MINI_ALU_nx479)) ;
    inv01 L1_1_L2_2_G1_MINI_ALU_ix478 (.Y (L1_1_L2_2_G1_MINI_ALU_nx477), .A (
          L1_1_L2_2_G1_MINI_ALU_BoothP_10)) ;
    xnor2 L1_1_L2_2_G1_MINI_ALU_ix480 (.Y (L1_1_L2_2_G1_MINI_ALU_nx479), .A0 (
          L1_1_L2_2_G1_MINI_ALU_BoothOperand_11), .A1 (
          L1_1_L2_2_G1_MINI_ALU_BoothP_11)) ;
    xor2 L1_1_L2_2_G1_MINI_ALU_ix377 (.Y (L1_1_L2_2_G1_MINI_ALU_nx376), .A0 (
         L1_1_L2_2_G1_MINI_ALU_nx483), .A1 (L1_1_L2_2_G1_MINI_ALU_nx487)) ;
    inv01 L1_1_L2_2_G1_MINI_ALU_ix486 (.Y (L1_1_L2_2_G1_MINI_ALU_nx485), .A (
          L1_1_L2_2_G1_MINI_ALU_BoothP_11)) ;
    xnor2 L1_1_L2_2_G1_MINI_ALU_ix488 (.Y (L1_1_L2_2_G1_MINI_ALU_nx487), .A0 (
          L1_1_L2_2_G1_MINI_ALU_BoothOperand_12), .A1 (
          L1_1_L2_2_G1_MINI_ALU_BoothP_12)) ;
    xor2 L1_1_L2_2_G1_MINI_ALU_ix397 (.Y (L1_1_L2_2_G1_MINI_ALU_nx396), .A0 (
         L1_1_L2_2_G1_MINI_ALU_nx491), .A1 (L1_1_L2_2_G1_MINI_ALU_nx495)) ;
    inv01 L1_1_L2_2_G1_MINI_ALU_ix494 (.Y (L1_1_L2_2_G1_MINI_ALU_nx493), .A (
          L1_1_L2_2_G1_MINI_ALU_BoothP_12)) ;
    xnor2 L1_1_L2_2_G1_MINI_ALU_ix496 (.Y (L1_1_L2_2_G1_MINI_ALU_nx495), .A0 (
          L1_1_L2_2_G1_MINI_ALU_BoothOperand_13), .A1 (
          L1_1_L2_2_G1_MINI_ALU_BoothP_13)) ;
    xor2 L1_1_L2_2_G1_MINI_ALU_ix417 (.Y (L1_1_L2_2_G1_MINI_ALU_nx416), .A0 (
         L1_1_L2_2_G1_MINI_ALU_nx499), .A1 (L1_1_L2_2_G1_MINI_ALU_nx503)) ;
    inv01 L1_1_L2_2_G1_MINI_ALU_ix502 (.Y (L1_1_L2_2_G1_MINI_ALU_nx501), .A (
          L1_1_L2_2_G1_MINI_ALU_BoothP_13)) ;
    xnor2 L1_1_L2_2_G1_MINI_ALU_ix504 (.Y (L1_1_L2_2_G1_MINI_ALU_nx503), .A0 (
          L1_1_L2_2_G1_MINI_ALU_BoothOperand_14), .A1 (
          L1_1_L2_2_G1_MINI_ALU_BoothP_14)) ;
    xor2 L1_1_L2_2_G1_MINI_ALU_ix437 (.Y (L1_1_L2_2_G1_MINI_ALU_nx436), .A0 (
         L1_1_L2_2_G1_MINI_ALU_nx507), .A1 (L1_1_L2_2_G1_MINI_ALU_nx511)) ;
    inv01 L1_1_L2_2_G1_MINI_ALU_ix510 (.Y (L1_1_L2_2_G1_MINI_ALU_nx509), .A (
          L1_1_L2_2_G1_MINI_ALU_BoothP_14)) ;
    xnor2 L1_1_L2_2_G1_MINI_ALU_ix512 (.Y (L1_1_L2_2_G1_MINI_ALU_nx511), .A0 (
          L1_1_L2_2_G1_MINI_ALU_BoothOperand_15), .A1 (
          L1_1_L2_2_G1_MINI_ALU_BoothP_15)) ;
    xnor2 L1_1_L2_2_G1_MINI_ALU_ix457 (.Y (L1_1_L2_2_G1_MINI_ALU_nx456), .A0 (
          L1_1_L2_2_G1_MINI_ALU_nx515), .A1 (L1_1_L2_2_G1_MINI_ALU_nx454)) ;
    inv01 L1_1_L2_2_G1_MINI_ALU_ix518 (.Y (L1_1_L2_2_G1_MINI_ALU_nx517), .A (
          L1_1_L2_2_G1_MINI_ALU_BoothP_15)) ;
    xor2 L1_1_L2_2_G1_MINI_ALU_ix455 (.Y (L1_1_L2_2_G1_MINI_ALU_nx454), .A0 (
         L1_1_L2_2_G1_MINI_ALU_BoothOperand_16), .A1 (
         L1_1_L2_2_G1_MINI_ALU_BoothP_16)) ;
    mux21_ni L1_1_L2_2_G1_MINI_ALU_ix91 (.Y (L1SecondOperands_7__0), .A0 (
             L1_1_L2_2_G1_MINI_ALU_BoothP_1), .A1 (WindowDin_1__2__0), .S0 (
             Instr)) ;
    mux21_ni L1_1_L2_2_G1_MINI_ALU_ix99 (.Y (L1SecondOperands_7__1), .A0 (
             L1_1_L2_2_G1_MINI_ALU_BoothP_2), .A1 (WindowDin_1__2__1), .S0 (
             Instr)) ;
    mux21_ni L1_1_L2_2_G1_MINI_ALU_ix107 (.Y (L1SecondOperands_7__2), .A0 (
             L1_1_L2_2_G1_MINI_ALU_BoothP_3), .A1 (WindowDin_1__2__2), .S0 (
             Instr)) ;
    mux21_ni L1_1_L2_2_G1_MINI_ALU_ix115 (.Y (L1SecondOperands_7__3), .A0 (
             L1_1_L2_2_G1_MINI_ALU_BoothP_4), .A1 (WindowDin_1__2__3), .S0 (
             Instr)) ;
    mux21_ni L1_1_L2_2_G1_MINI_ALU_ix123 (.Y (L1SecondOperands_7__4), .A0 (
             L1_1_L2_2_G1_MINI_ALU_BoothP_5), .A1 (WindowDin_1__2__4), .S0 (
             Instr)) ;
    mux21_ni L1_1_L2_2_G1_MINI_ALU_ix131 (.Y (L1SecondOperands_7__5), .A0 (
             L1_1_L2_2_G1_MINI_ALU_BoothP_6), .A1 (WindowDin_1__2__5), .S0 (
             Instr)) ;
    mux21_ni L1_1_L2_2_G1_MINI_ALU_ix139 (.Y (L1SecondOperands_7__6), .A0 (
             L1_1_L2_2_G1_MINI_ALU_BoothP_7), .A1 (WindowDin_1__2__6), .S0 (
             Instr)) ;
    mux21_ni L1_1_L2_2_G1_MINI_ALU_ix147 (.Y (L1SecondOperands_7__7), .A0 (
             L1_1_L2_2_G1_MINI_ALU_BoothP_8), .A1 (WindowDin_1__2__7), .S0 (
             Instr)) ;
    xor2 L1_1_L2_2_G1_MINI_ALU_ix77 (.Y (L1Results_7__1), .A0 (
         L1_1_L2_2_G1_MINI_ALU_nx529), .A1 (L1_1_L2_2_G1_MINI_ALU_nx531)) ;
    nand02 L1_1_L2_2_G1_MINI_ALU_ix530 (.Y (L1_1_L2_2_G1_MINI_ALU_nx529), .A0 (
           L1SecondOperands_7__0), .A1 (L1FirstOperands_7__0)) ;
    xnor2 L1_1_L2_2_G1_MINI_ALU_ix532 (.Y (L1_1_L2_2_G1_MINI_ALU_nx531), .A0 (
          L1SecondOperands_7__1), .A1 (L1FirstOperands_7__1)) ;
    xor2 L1_1_L2_2_G1_MINI_ALU_ix75 (.Y (L1Results_7__2), .A0 (
         L1_1_L2_2_G1_MINI_ALU_nx534), .A1 (L1_1_L2_2_G1_MINI_ALU_nx537)) ;
    aoi32 L1_1_L2_2_G1_MINI_ALU_ix535 (.Y (L1_1_L2_2_G1_MINI_ALU_nx534), .A0 (
          L1SecondOperands_7__0), .A1 (L1FirstOperands_7__0), .A2 (
          L1_1_L2_2_G1_MINI_ALU_nx30), .B0 (L1FirstOperands_7__1), .B1 (
          L1SecondOperands_7__1)) ;
    xnor2 L1_1_L2_2_G1_MINI_ALU_ix538 (.Y (L1_1_L2_2_G1_MINI_ALU_nx537), .A0 (
          L1SecondOperands_7__2), .A1 (L1FirstOperands_7__2)) ;
    xor2 L1_1_L2_2_G1_MINI_ALU_ix73 (.Y (L1Results_7__3), .A0 (
         L1_1_L2_2_G1_MINI_ALU_nx540), .A1 (L1_1_L2_2_G1_MINI_ALU_nx544)) ;
    aoi22 L1_1_L2_2_G1_MINI_ALU_ix541 (.Y (L1_1_L2_2_G1_MINI_ALU_nx540), .A0 (
          L1FirstOperands_7__2), .A1 (L1SecondOperands_7__2), .B0 (
          L1_1_L2_2_G1_MINI_ALU_nx40), .B1 (L1_1_L2_2_G1_MINI_ALU_nx24)) ;
    xnor2 L1_1_L2_2_G1_MINI_ALU_ix545 (.Y (L1_1_L2_2_G1_MINI_ALU_nx544), .A0 (
          L1SecondOperands_7__3), .A1 (L1FirstOperands_7__3)) ;
    xor2 L1_1_L2_2_G1_MINI_ALU_ix71 (.Y (L1Results_7__4), .A0 (
         L1_1_L2_2_G1_MINI_ALU_nx547), .A1 (L1_1_L2_2_G1_MINI_ALU_nx551)) ;
    aoi22 L1_1_L2_2_G1_MINI_ALU_ix548 (.Y (L1_1_L2_2_G1_MINI_ALU_nx547), .A0 (
          L1FirstOperands_7__3), .A1 (L1SecondOperands_7__3), .B0 (
          L1_1_L2_2_G1_MINI_ALU_nx44), .B1 (L1_1_L2_2_G1_MINI_ALU_nx18)) ;
    xnor2 L1_1_L2_2_G1_MINI_ALU_ix552 (.Y (L1_1_L2_2_G1_MINI_ALU_nx551), .A0 (
          L1SecondOperands_7__4), .A1 (L1FirstOperands_7__4)) ;
    xor2 L1_1_L2_2_G1_MINI_ALU_ix69 (.Y (L1Results_7__5), .A0 (
         L1_1_L2_2_G1_MINI_ALU_nx554), .A1 (L1_1_L2_2_G1_MINI_ALU_nx558)) ;
    aoi22 L1_1_L2_2_G1_MINI_ALU_ix555 (.Y (L1_1_L2_2_G1_MINI_ALU_nx554), .A0 (
          L1FirstOperands_7__4), .A1 (L1SecondOperands_7__4), .B0 (
          L1_1_L2_2_G1_MINI_ALU_nx48), .B1 (L1_1_L2_2_G1_MINI_ALU_nx12)) ;
    xnor2 L1_1_L2_2_G1_MINI_ALU_ix559 (.Y (L1_1_L2_2_G1_MINI_ALU_nx558), .A0 (
          L1SecondOperands_7__5), .A1 (L1FirstOperands_7__5)) ;
    xor2 L1_1_L2_2_G1_MINI_ALU_ix67 (.Y (L1Results_7__6), .A0 (
         L1_1_L2_2_G1_MINI_ALU_nx561), .A1 (L1_1_L2_2_G1_MINI_ALU_nx565)) ;
    aoi22 L1_1_L2_2_G1_MINI_ALU_ix562 (.Y (L1_1_L2_2_G1_MINI_ALU_nx561), .A0 (
          L1FirstOperands_7__5), .A1 (L1SecondOperands_7__5), .B0 (
          L1_1_L2_2_G1_MINI_ALU_nx52), .B1 (L1_1_L2_2_G1_MINI_ALU_nx6)) ;
    xnor2 L1_1_L2_2_G1_MINI_ALU_ix566 (.Y (L1_1_L2_2_G1_MINI_ALU_nx565), .A0 (
          L1SecondOperands_7__6), .A1 (L1FirstOperands_7__6)) ;
    xnor2 L1_1_L2_2_G1_MINI_ALU_ix65 (.Y (L1Results_7__7), .A0 (
          L1_1_L2_2_G1_MINI_ALU_nx568), .A1 (L1_1_L2_2_G1_MINI_ALU_nx62)) ;
    aoi22 L1_1_L2_2_G1_MINI_ALU_ix569 (.Y (L1_1_L2_2_G1_MINI_ALU_nx568), .A0 (
          L1FirstOperands_7__6), .A1 (L1SecondOperands_7__6), .B0 (
          L1_1_L2_2_G1_MINI_ALU_nx56), .B1 (L1_1_L2_2_G1_MINI_ALU_nx0)) ;
    xor2 L1_1_L2_2_G1_MINI_ALU_ix63 (.Y (L1_1_L2_2_G1_MINI_ALU_nx62), .A0 (
         L1SecondOperands_7__7), .A1 (L1FirstOperands_7__7)) ;
    inv01 L1_1_L2_2_G1_MINI_ALU_ix155 (.Y (L1_1_L2_2_G1_MINI_ALU_nx154), .A (
          L1_1_L2_2_G1_MINI_ALU_nx383)) ;
    inv01 L1_1_L2_2_G1_MINI_ALU_ix57 (.Y (L1_1_L2_2_G1_MINI_ALU_nx56), .A (
          L1_1_L2_2_G1_MINI_ALU_nx561)) ;
    inv01 L1_1_L2_2_G1_MINI_ALU_ix53 (.Y (L1_1_L2_2_G1_MINI_ALU_nx52), .A (
          L1_1_L2_2_G1_MINI_ALU_nx554)) ;
    inv01 L1_1_L2_2_G1_MINI_ALU_ix49 (.Y (L1_1_L2_2_G1_MINI_ALU_nx48), .A (
          L1_1_L2_2_G1_MINI_ALU_nx547)) ;
    inv01 L1_1_L2_2_G1_MINI_ALU_ix45 (.Y (L1_1_L2_2_G1_MINI_ALU_nx44), .A (
          L1_1_L2_2_G1_MINI_ALU_nx540)) ;
    inv01 L1_1_L2_2_G1_MINI_ALU_ix41 (.Y (L1_1_L2_2_G1_MINI_ALU_nx40), .A (
          L1_1_L2_2_G1_MINI_ALU_nx534)) ;
    inv01 L1_1_L2_2_G1_MINI_ALU_ix31 (.Y (L1_1_L2_2_G1_MINI_ALU_nx30), .A (
          L1_1_L2_2_G1_MINI_ALU_nx531)) ;
    inv01 L1_1_L2_2_G1_MINI_ALU_ix25 (.Y (L1_1_L2_2_G1_MINI_ALU_nx24), .A (
          L1_1_L2_2_G1_MINI_ALU_nx537)) ;
    inv01 L1_1_L2_2_G1_MINI_ALU_ix19 (.Y (L1_1_L2_2_G1_MINI_ALU_nx18), .A (
          L1_1_L2_2_G1_MINI_ALU_nx544)) ;
    inv01 L1_1_L2_2_G1_MINI_ALU_ix13 (.Y (L1_1_L2_2_G1_MINI_ALU_nx12), .A (
          L1_1_L2_2_G1_MINI_ALU_nx551)) ;
    inv01 L1_1_L2_2_G1_MINI_ALU_ix7 (.Y (L1_1_L2_2_G1_MINI_ALU_nx6), .A (
          L1_1_L2_2_G1_MINI_ALU_nx558)) ;
    inv01 L1_1_L2_2_G1_MINI_ALU_ix1 (.Y (L1_1_L2_2_G1_MINI_ALU_nx0), .A (
          L1_1_L2_2_G1_MINI_ALU_nx565)) ;
    fake_gnd L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix216 (.Y (
             L1_1_L2_2_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    nor02ii L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix81 (.Y (
            L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx80), .A0 (Instr), .A1 (Start)) ;
    aoi21 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix77 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_10), .A0 (
          FilterDin_1__2__1), .A1 (FilterDin_1__2__0), .B0 (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx4)) ;
    nor02_2x L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix5 (.Y (
             L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx4), .A0 (FilterDin_1__2__0), .A1 (
             FilterDin_1__2__1)) ;
    aoi21 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix67 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_11), .A0 (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx328), .A1 (FilterDin_1__2__2), .B0 (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx8)) ;
    nor03_2x L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix9 (.Y (
             L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx8), .A0 (FilterDin_1__2__2), .A1 (
             FilterDin_1__2__0), .A2 (FilterDin_1__2__1)) ;
    xnor2 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix59 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_12), .A0 (
          FilterDin_1__2__3), .A1 (L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx8)) ;
    xnor2 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix51 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_13), .A0 (
          FilterDin_1__2__4), .A1 (L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx12)) ;
    nor04 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix13 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx12), .A0 (FilterDin_1__2__3), .A1 (
          FilterDin_1__2__2), .A2 (FilterDin_1__2__0), .A3 (FilterDin_1__2__1)
          ) ;
    xnor2 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix43 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_14), .A0 (
          FilterDin_1__2__5), .A1 (L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx16)) ;
    nor02ii L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix17 (.Y (
            L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx16), .A0 (FilterDin_1__2__4), .A1 (
            L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx12)) ;
    xnor2 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix35 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_15), .A0 (
          FilterDin_1__2__6), .A1 (L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx20)) ;
    nor02ii L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix21 (.Y (
            L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx20), .A0 (FilterDin_1__2__5), .A1 (
            L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx16)) ;
    xnor2 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix27 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_16), .A0 (
          FilterDin_1__2__7), .A1 (L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx24)) ;
    nor02ii L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix25 (.Y (
            L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx24), .A0 (FilterDin_1__2__6), .A1 (
            L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx20)) ;
    inv01 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix329 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx328), .A (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx4)) ;
    inv02 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix383 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx384), .A (
          L1_1_L2_2_G1_MINI_ALU_BoothP_0)) ;
    dff L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_0 (.Q (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_0), .QB (\$dummy [361]), 
        .D (L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .CLK (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    nor02_2x L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix567 (.Y (
             L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566), .A0 (RST), .A1 (
             L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644)) ;
    dff L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_1 (.Q (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_1), .QB (\$dummy [362]), 
        .D (L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .CLK (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_2 (.Q (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_2), .QB (\$dummy [363]), 
        .D (L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .CLK (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_3 (.Q (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_3), .QB (\$dummy [364]), 
        .D (L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .CLK (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_4 (.Q (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_4), .QB (\$dummy [365]), 
        .D (L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .CLK (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_5 (.Q (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_5), .QB (\$dummy [366]), 
        .D (L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .CLK (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_6 (.Q (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_6), .QB (\$dummy [367]), 
        .D (L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .CLK (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_7 (.Q (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_7), .QB (\$dummy [368]), 
        .D (L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .CLK (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_8 (.Q (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_8), .QB (\$dummy [369]), 
        .D (L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .CLK (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_9 (.Q (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_9), .QB (\$dummy [370]), 
        .D (L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .CLK (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_10 (.Q (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_10), .QB (\$dummy [371])
        , .D (L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .CLK (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_11 (.Q (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_11), .QB (\$dummy [372])
        , .D (L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .CLK (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_12 (.Q (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_12), .QB (\$dummy [373])
        , .D (L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .CLK (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_13 (.Q (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_13), .QB (\$dummy [374])
        , .D (L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .CLK (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_14 (.Q (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_14), .QB (\$dummy [375])
        , .D (L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .CLK (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_15 (.Q (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_15), .QB (\$dummy [376])
        , .D (L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .CLK (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_16 (.Q (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_16), .QB (\$dummy [377])
        , .D (L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .CLK (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    inv02 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix623 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624), .A (CLK)) ;
    inv02 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix625 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626), .A (CLK)) ;
    inv02 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix627 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628), .A (CLK)) ;
    inv02 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix643 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644), .A (nx7898)) ;
    dff L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_0 (.Q (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_0), .QB (\$dummy [378]), 
        .D (L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .CLK (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    nor02_2x L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix567 (.Y (
             L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566), .A0 (RST), .A1 (
             L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644)) ;
    dff L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_1 (.Q (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_1), .QB (\$dummy [379]), 
        .D (L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .CLK (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_2 (.Q (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_2), .QB (\$dummy [380]), 
        .D (L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .CLK (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_3 (.Q (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_3), .QB (\$dummy [381]), 
        .D (L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .CLK (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_4 (.Q (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_4), .QB (\$dummy [382]), 
        .D (L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .CLK (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_5 (.Q (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_5), .QB (\$dummy [383]), 
        .D (L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .CLK (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_6 (.Q (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_6), .QB (\$dummy [384]), 
        .D (L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .CLK (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_7 (.Q (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_7), .QB (\$dummy [385]), 
        .D (L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .CLK (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_8 (.Q (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_8), .QB (\$dummy [386]), 
        .D (L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .CLK (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_9 (.Q (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_9), .QB (\$dummy [387]), 
        .D (L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .CLK (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_10 (.Q (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_10), .QB (\$dummy [388])
        , .D (L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .CLK (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_11 (.Q (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_11), .QB (\$dummy [389])
        , .D (L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .CLK (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_12 (.Q (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_12), .QB (\$dummy [390])
        , .D (L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .CLK (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_13 (.Q (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_13), .QB (\$dummy [391])
        , .D (L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .CLK (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_14 (.Q (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_14), .QB (\$dummy [392])
        , .D (L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .CLK (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_15 (.Q (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_15), .QB (\$dummy [393])
        , .D (L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .CLK (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_16 (.Q (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_16), .QB (\$dummy [394])
        , .D (L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .CLK (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    inv02 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix623 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624), .A (CLK)) ;
    inv02 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix625 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626), .A (CLK)) ;
    inv02 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix627 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628), .A (CLK)) ;
    inv02 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix643 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644), .A (nx7904)) ;
    dff L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_0 (.Q (
        L1_1_L2_2_G1_MINI_ALU_BoothP_0), .QB (\$dummy [395]), .D (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .CLK (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    nor02_2x L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix567 (.Y (
             L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566), .A0 (RST), .A1 (
             L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    dff L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_1 (.Q (
        L1_1_L2_2_G1_MINI_ALU_BoothP_1), .QB (\$dummy [396]), .D (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .CLK (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_2 (.Q (
        L1_1_L2_2_G1_MINI_ALU_BoothP_2), .QB (\$dummy [397]), .D (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .CLK (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_3 (.Q (
        L1_1_L2_2_G1_MINI_ALU_BoothP_3), .QB (\$dummy [398]), .D (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .CLK (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_4 (.Q (
        L1_1_L2_2_G1_MINI_ALU_BoothP_4), .QB (\$dummy [399]), .D (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .CLK (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_5 (.Q (
        L1_1_L2_2_G1_MINI_ALU_BoothP_5), .QB (\$dummy [400]), .D (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .CLK (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_6 (.Q (
        L1_1_L2_2_G1_MINI_ALU_BoothP_6), .QB (\$dummy [401]), .D (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .CLK (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_7 (.Q (
        L1_1_L2_2_G1_MINI_ALU_BoothP_7), .QB (\$dummy [402]), .D (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .CLK (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_8 (.Q (
        L1_1_L2_2_G1_MINI_ALU_BoothP_8), .QB (\$dummy [403]), .D (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .CLK (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_9 (.Q (
        L1_1_L2_2_G1_MINI_ALU_BoothP_9), .QB (\$dummy [404]), .D (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .CLK (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_10 (.Q (
        L1_1_L2_2_G1_MINI_ALU_BoothP_10), .QB (\$dummy [405]), .D (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .CLK (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_11 (.Q (
        L1_1_L2_2_G1_MINI_ALU_BoothP_11), .QB (\$dummy [406]), .D (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .CLK (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_12 (.Q (
        L1_1_L2_2_G1_MINI_ALU_BoothP_12), .QB (\$dummy [407]), .D (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .CLK (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_13 (.Q (
        L1_1_L2_2_G1_MINI_ALU_BoothP_13), .QB (\$dummy [408]), .D (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .CLK (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_14 (.Q (
        L1_1_L2_2_G1_MINI_ALU_BoothP_14), .QB (\$dummy [409]), .D (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .CLK (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_15 (.Q (
        L1_1_L2_2_G1_MINI_ALU_BoothP_15), .QB (\$dummy [410]), .D (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .CLK (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_16 (.Q (
        L1_1_L2_2_G1_MINI_ALU_BoothP_16), .QB (\$dummy [411]), .D (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .CLK (
        L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    inv02 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix623 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624), .A (CLK)) ;
    inv02 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix625 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626), .A (CLK)) ;
    inv02 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix627 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628), .A (CLK)) ;
    inv02 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix643 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644), .A (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642)) ;
    xor2 L1_1_L2_3_G1_MINI_ALU_ix83 (.Y (L1Results_8__0), .A0 (
         L1SecondOperands_8__0), .A1 (L1FirstOperands_8__0)) ;
    xnor2 L1_1_L2_3_G1_MINI_ALU_ix380 (.Y (L1_1_L2_3_G1_MINI_ALU_nx379), .A0 (
          L1_1_L2_3_G1_MINI_ALU_nx381), .A1 (L1_1_L2_3_G1_MINI_ALU_nx383)) ;
    nand02 L1_1_L2_3_G1_MINI_ALU_ix382 (.Y (L1_1_L2_3_G1_MINI_ALU_nx381), .A0 (
           L1_1_L2_3_G1_MINI_ALU_BoothOperand_0), .A1 (nx7924)) ;
    xnor2 L1_1_L2_3_G1_MINI_ALU_ix384 (.Y (L1_1_L2_3_G1_MINI_ALU_nx383), .A0 (
          L1_1_L2_3_G1_MINI_ALU_BoothOperand_1), .A1 (
          L1_1_L2_3_G1_MINI_ALU_BoothP_1)) ;
    inv01 L1_1_L2_3_G1_MINI_ALU_ix388 (.Y (L1_1_L2_3_G1_MINI_ALU_nx387), .A (
          L1_1_L2_3_G1_MINI_ALU_BoothP_2)) ;
    xnor2 L1_1_L2_3_G1_MINI_ALU_ix390 (.Y (L1_1_L2_3_G1_MINI_ALU_nx389), .A0 (
          L1_1_L2_3_G1_MINI_ALU_nx391), .A1 (L1_1_L2_3_G1_MINI_ALU_nx395)) ;
    aoi32 L1_1_L2_3_G1_MINI_ALU_ix392 (.Y (L1_1_L2_3_G1_MINI_ALU_nx391), .A0 (
          L1_1_L2_3_G1_MINI_ALU_BoothOperand_0), .A1 (nx7924), .A2 (
          L1_1_L2_3_G1_MINI_ALU_nx154), .B0 (L1_1_L2_3_G1_MINI_ALU_BoothP_1), .B1 (
          L1_1_L2_3_G1_MINI_ALU_BoothOperand_1)) ;
    xnor2 L1_1_L2_3_G1_MINI_ALU_ix396 (.Y (L1_1_L2_3_G1_MINI_ALU_nx395), .A0 (
          L1_1_L2_3_G1_MINI_ALU_BoothOperand_2), .A1 (
          L1_1_L2_3_G1_MINI_ALU_BoothP_2)) ;
    inv01 L1_1_L2_3_G1_MINI_ALU_ix400 (.Y (L1_1_L2_3_G1_MINI_ALU_nx399), .A (
          L1_1_L2_3_G1_MINI_ALU_BoothP_3)) ;
    xnor2 L1_1_L2_3_G1_MINI_ALU_ix402 (.Y (L1_1_L2_3_G1_MINI_ALU_nx401), .A0 (
          L1_1_L2_3_G1_MINI_ALU_nx403), .A1 (L1_1_L2_3_G1_MINI_ALU_nx405)) ;
    xnor2 L1_1_L2_3_G1_MINI_ALU_ix406 (.Y (L1_1_L2_3_G1_MINI_ALU_nx405), .A0 (
          L1_1_L2_3_G1_MINI_ALU_BoothOperand_3), .A1 (
          L1_1_L2_3_G1_MINI_ALU_BoothP_3)) ;
    inv01 L1_1_L2_3_G1_MINI_ALU_ix410 (.Y (L1_1_L2_3_G1_MINI_ALU_nx409), .A (
          L1_1_L2_3_G1_MINI_ALU_BoothP_4)) ;
    xnor2 L1_1_L2_3_G1_MINI_ALU_ix412 (.Y (L1_1_L2_3_G1_MINI_ALU_nx411), .A0 (
          L1_1_L2_3_G1_MINI_ALU_nx413), .A1 (L1_1_L2_3_G1_MINI_ALU_nx415)) ;
    xnor2 L1_1_L2_3_G1_MINI_ALU_ix416 (.Y (L1_1_L2_3_G1_MINI_ALU_nx415), .A0 (
          L1_1_L2_3_G1_MINI_ALU_BoothOperand_4), .A1 (
          L1_1_L2_3_G1_MINI_ALU_BoothP_4)) ;
    inv01 L1_1_L2_3_G1_MINI_ALU_ix420 (.Y (L1_1_L2_3_G1_MINI_ALU_nx419), .A (
          L1_1_L2_3_G1_MINI_ALU_BoothP_5)) ;
    xnor2 L1_1_L2_3_G1_MINI_ALU_ix422 (.Y (L1_1_L2_3_G1_MINI_ALU_nx421), .A0 (
          L1_1_L2_3_G1_MINI_ALU_nx423), .A1 (L1_1_L2_3_G1_MINI_ALU_nx425)) ;
    xnor2 L1_1_L2_3_G1_MINI_ALU_ix426 (.Y (L1_1_L2_3_G1_MINI_ALU_nx425), .A0 (
          L1_1_L2_3_G1_MINI_ALU_BoothOperand_5), .A1 (
          L1_1_L2_3_G1_MINI_ALU_BoothP_5)) ;
    inv01 L1_1_L2_3_G1_MINI_ALU_ix430 (.Y (L1_1_L2_3_G1_MINI_ALU_nx429), .A (
          L1_1_L2_3_G1_MINI_ALU_BoothP_6)) ;
    xnor2 L1_1_L2_3_G1_MINI_ALU_ix432 (.Y (L1_1_L2_3_G1_MINI_ALU_nx431), .A0 (
          L1_1_L2_3_G1_MINI_ALU_nx433), .A1 (L1_1_L2_3_G1_MINI_ALU_nx435)) ;
    xnor2 L1_1_L2_3_G1_MINI_ALU_ix436 (.Y (L1_1_L2_3_G1_MINI_ALU_nx435), .A0 (
          L1_1_L2_3_G1_MINI_ALU_BoothOperand_6), .A1 (
          L1_1_L2_3_G1_MINI_ALU_BoothP_6)) ;
    inv01 L1_1_L2_3_G1_MINI_ALU_ix440 (.Y (L1_1_L2_3_G1_MINI_ALU_nx439), .A (
          L1_1_L2_3_G1_MINI_ALU_BoothP_7)) ;
    xnor2 L1_1_L2_3_G1_MINI_ALU_ix442 (.Y (L1_1_L2_3_G1_MINI_ALU_nx441), .A0 (
          L1_1_L2_3_G1_MINI_ALU_nx443), .A1 (L1_1_L2_3_G1_MINI_ALU_nx445)) ;
    xnor2 L1_1_L2_3_G1_MINI_ALU_ix446 (.Y (L1_1_L2_3_G1_MINI_ALU_nx445), .A0 (
          L1_1_L2_3_G1_MINI_ALU_BoothOperand_7), .A1 (
          L1_1_L2_3_G1_MINI_ALU_BoothP_7)) ;
    inv01 L1_1_L2_3_G1_MINI_ALU_ix450 (.Y (L1_1_L2_3_G1_MINI_ALU_nx449), .A (
          L1_1_L2_3_G1_MINI_ALU_BoothP_8)) ;
    xnor2 L1_1_L2_3_G1_MINI_ALU_ix452 (.Y (L1_1_L2_3_G1_MINI_ALU_nx451), .A0 (
          L1_1_L2_3_G1_MINI_ALU_nx453), .A1 (L1_1_L2_3_G1_MINI_ALU_nx455)) ;
    xnor2 L1_1_L2_3_G1_MINI_ALU_ix456 (.Y (L1_1_L2_3_G1_MINI_ALU_nx455), .A0 (
          L1_1_L2_3_G1_MINI_ALU_BoothOperand_8), .A1 (
          L1_1_L2_3_G1_MINI_ALU_BoothP_8)) ;
    xor2 L1_1_L2_3_G1_MINI_ALU_ix317 (.Y (L1_1_L2_3_G1_MINI_ALU_nx316), .A0 (
         L1_1_L2_3_G1_MINI_ALU_nx461), .A1 (L1_1_L2_3_G1_MINI_ALU_nx463)) ;
    xnor2 L1_1_L2_3_G1_MINI_ALU_ix464 (.Y (L1_1_L2_3_G1_MINI_ALU_nx463), .A0 (
          L1_1_L2_3_G1_MINI_ALU_BoothOperand_9), .A1 (
          L1_1_L2_3_G1_MINI_ALU_BoothP_9)) ;
    xor2 L1_1_L2_3_G1_MINI_ALU_ix337 (.Y (L1_1_L2_3_G1_MINI_ALU_nx336), .A0 (
         L1_1_L2_3_G1_MINI_ALU_nx467), .A1 (L1_1_L2_3_G1_MINI_ALU_nx471)) ;
    inv01 L1_1_L2_3_G1_MINI_ALU_ix470 (.Y (L1_1_L2_3_G1_MINI_ALU_nx469), .A (
          L1_1_L2_3_G1_MINI_ALU_BoothP_9)) ;
    xnor2 L1_1_L2_3_G1_MINI_ALU_ix472 (.Y (L1_1_L2_3_G1_MINI_ALU_nx471), .A0 (
          L1_1_L2_3_G1_MINI_ALU_BoothOperand_10), .A1 (
          L1_1_L2_3_G1_MINI_ALU_BoothP_10)) ;
    xor2 L1_1_L2_3_G1_MINI_ALU_ix357 (.Y (L1_1_L2_3_G1_MINI_ALU_nx356), .A0 (
         L1_1_L2_3_G1_MINI_ALU_nx475), .A1 (L1_1_L2_3_G1_MINI_ALU_nx479)) ;
    inv01 L1_1_L2_3_G1_MINI_ALU_ix478 (.Y (L1_1_L2_3_G1_MINI_ALU_nx477), .A (
          L1_1_L2_3_G1_MINI_ALU_BoothP_10)) ;
    xnor2 L1_1_L2_3_G1_MINI_ALU_ix480 (.Y (L1_1_L2_3_G1_MINI_ALU_nx479), .A0 (
          L1_1_L2_3_G1_MINI_ALU_BoothOperand_11), .A1 (
          L1_1_L2_3_G1_MINI_ALU_BoothP_11)) ;
    xor2 L1_1_L2_3_G1_MINI_ALU_ix377 (.Y (L1_1_L2_3_G1_MINI_ALU_nx376), .A0 (
         L1_1_L2_3_G1_MINI_ALU_nx483), .A1 (L1_1_L2_3_G1_MINI_ALU_nx487)) ;
    inv01 L1_1_L2_3_G1_MINI_ALU_ix486 (.Y (L1_1_L2_3_G1_MINI_ALU_nx485), .A (
          L1_1_L2_3_G1_MINI_ALU_BoothP_11)) ;
    xnor2 L1_1_L2_3_G1_MINI_ALU_ix488 (.Y (L1_1_L2_3_G1_MINI_ALU_nx487), .A0 (
          L1_1_L2_3_G1_MINI_ALU_BoothOperand_12), .A1 (
          L1_1_L2_3_G1_MINI_ALU_BoothP_12)) ;
    xor2 L1_1_L2_3_G1_MINI_ALU_ix397 (.Y (L1_1_L2_3_G1_MINI_ALU_nx396), .A0 (
         L1_1_L2_3_G1_MINI_ALU_nx491), .A1 (L1_1_L2_3_G1_MINI_ALU_nx495)) ;
    inv01 L1_1_L2_3_G1_MINI_ALU_ix494 (.Y (L1_1_L2_3_G1_MINI_ALU_nx493), .A (
          L1_1_L2_3_G1_MINI_ALU_BoothP_12)) ;
    xnor2 L1_1_L2_3_G1_MINI_ALU_ix496 (.Y (L1_1_L2_3_G1_MINI_ALU_nx495), .A0 (
          L1_1_L2_3_G1_MINI_ALU_BoothOperand_13), .A1 (
          L1_1_L2_3_G1_MINI_ALU_BoothP_13)) ;
    xor2 L1_1_L2_3_G1_MINI_ALU_ix417 (.Y (L1_1_L2_3_G1_MINI_ALU_nx416), .A0 (
         L1_1_L2_3_G1_MINI_ALU_nx499), .A1 (L1_1_L2_3_G1_MINI_ALU_nx503)) ;
    inv01 L1_1_L2_3_G1_MINI_ALU_ix502 (.Y (L1_1_L2_3_G1_MINI_ALU_nx501), .A (
          L1_1_L2_3_G1_MINI_ALU_BoothP_13)) ;
    xnor2 L1_1_L2_3_G1_MINI_ALU_ix504 (.Y (L1_1_L2_3_G1_MINI_ALU_nx503), .A0 (
          L1_1_L2_3_G1_MINI_ALU_BoothOperand_14), .A1 (
          L1_1_L2_3_G1_MINI_ALU_BoothP_14)) ;
    xor2 L1_1_L2_3_G1_MINI_ALU_ix437 (.Y (L1_1_L2_3_G1_MINI_ALU_nx436), .A0 (
         L1_1_L2_3_G1_MINI_ALU_nx507), .A1 (L1_1_L2_3_G1_MINI_ALU_nx511)) ;
    inv01 L1_1_L2_3_G1_MINI_ALU_ix510 (.Y (L1_1_L2_3_G1_MINI_ALU_nx509), .A (
          L1_1_L2_3_G1_MINI_ALU_BoothP_14)) ;
    xnor2 L1_1_L2_3_G1_MINI_ALU_ix512 (.Y (L1_1_L2_3_G1_MINI_ALU_nx511), .A0 (
          L1_1_L2_3_G1_MINI_ALU_BoothOperand_15), .A1 (
          L1_1_L2_3_G1_MINI_ALU_BoothP_15)) ;
    xnor2 L1_1_L2_3_G1_MINI_ALU_ix457 (.Y (L1_1_L2_3_G1_MINI_ALU_nx456), .A0 (
          L1_1_L2_3_G1_MINI_ALU_nx515), .A1 (L1_1_L2_3_G1_MINI_ALU_nx454)) ;
    inv01 L1_1_L2_3_G1_MINI_ALU_ix518 (.Y (L1_1_L2_3_G1_MINI_ALU_nx517), .A (
          L1_1_L2_3_G1_MINI_ALU_BoothP_15)) ;
    xor2 L1_1_L2_3_G1_MINI_ALU_ix455 (.Y (L1_1_L2_3_G1_MINI_ALU_nx454), .A0 (
         L1_1_L2_3_G1_MINI_ALU_BoothOperand_16), .A1 (
         L1_1_L2_3_G1_MINI_ALU_BoothP_16)) ;
    mux21_ni L1_1_L2_3_G1_MINI_ALU_ix91 (.Y (L1SecondOperands_8__0), .A0 (
             L1_1_L2_3_G1_MINI_ALU_BoothP_1), .A1 (WindowDin_1__3__0), .S0 (
             Instr)) ;
    mux21_ni L1_1_L2_3_G1_MINI_ALU_ix99 (.Y (L1SecondOperands_8__1), .A0 (
             L1_1_L2_3_G1_MINI_ALU_BoothP_2), .A1 (WindowDin_1__3__1), .S0 (
             Instr)) ;
    mux21_ni L1_1_L2_3_G1_MINI_ALU_ix107 (.Y (L1SecondOperands_8__2), .A0 (
             L1_1_L2_3_G1_MINI_ALU_BoothP_3), .A1 (WindowDin_1__3__2), .S0 (
             Instr)) ;
    mux21_ni L1_1_L2_3_G1_MINI_ALU_ix115 (.Y (L1SecondOperands_8__3), .A0 (
             L1_1_L2_3_G1_MINI_ALU_BoothP_4), .A1 (WindowDin_1__3__3), .S0 (
             Instr)) ;
    mux21_ni L1_1_L2_3_G1_MINI_ALU_ix123 (.Y (L1SecondOperands_8__4), .A0 (
             L1_1_L2_3_G1_MINI_ALU_BoothP_5), .A1 (WindowDin_1__3__4), .S0 (
             Instr)) ;
    mux21_ni L1_1_L2_3_G1_MINI_ALU_ix131 (.Y (L1SecondOperands_8__5), .A0 (
             L1_1_L2_3_G1_MINI_ALU_BoothP_6), .A1 (WindowDin_1__3__5), .S0 (
             Instr)) ;
    mux21_ni L1_1_L2_3_G1_MINI_ALU_ix139 (.Y (L1SecondOperands_8__6), .A0 (
             L1_1_L2_3_G1_MINI_ALU_BoothP_7), .A1 (WindowDin_1__3__6), .S0 (
             Instr)) ;
    mux21_ni L1_1_L2_3_G1_MINI_ALU_ix147 (.Y (L1SecondOperands_8__7), .A0 (
             L1_1_L2_3_G1_MINI_ALU_BoothP_8), .A1 (WindowDin_1__3__7), .S0 (
             Instr)) ;
    xor2 L1_1_L2_3_G1_MINI_ALU_ix77 (.Y (L1Results_8__1), .A0 (
         L1_1_L2_3_G1_MINI_ALU_nx529), .A1 (L1_1_L2_3_G1_MINI_ALU_nx531)) ;
    nand02 L1_1_L2_3_G1_MINI_ALU_ix530 (.Y (L1_1_L2_3_G1_MINI_ALU_nx529), .A0 (
           L1SecondOperands_8__0), .A1 (L1FirstOperands_8__0)) ;
    xnor2 L1_1_L2_3_G1_MINI_ALU_ix532 (.Y (L1_1_L2_3_G1_MINI_ALU_nx531), .A0 (
          L1SecondOperands_8__1), .A1 (L1FirstOperands_8__1)) ;
    xor2 L1_1_L2_3_G1_MINI_ALU_ix75 (.Y (L1Results_8__2), .A0 (
         L1_1_L2_3_G1_MINI_ALU_nx534), .A1 (L1_1_L2_3_G1_MINI_ALU_nx537)) ;
    aoi32 L1_1_L2_3_G1_MINI_ALU_ix535 (.Y (L1_1_L2_3_G1_MINI_ALU_nx534), .A0 (
          L1SecondOperands_8__0), .A1 (L1FirstOperands_8__0), .A2 (
          L1_1_L2_3_G1_MINI_ALU_nx30), .B0 (L1FirstOperands_8__1), .B1 (
          L1SecondOperands_8__1)) ;
    xnor2 L1_1_L2_3_G1_MINI_ALU_ix538 (.Y (L1_1_L2_3_G1_MINI_ALU_nx537), .A0 (
          L1SecondOperands_8__2), .A1 (L1FirstOperands_8__2)) ;
    xor2 L1_1_L2_3_G1_MINI_ALU_ix73 (.Y (L1Results_8__3), .A0 (
         L1_1_L2_3_G1_MINI_ALU_nx540), .A1 (L1_1_L2_3_G1_MINI_ALU_nx544)) ;
    aoi22 L1_1_L2_3_G1_MINI_ALU_ix541 (.Y (L1_1_L2_3_G1_MINI_ALU_nx540), .A0 (
          L1FirstOperands_8__2), .A1 (L1SecondOperands_8__2), .B0 (
          L1_1_L2_3_G1_MINI_ALU_nx40), .B1 (L1_1_L2_3_G1_MINI_ALU_nx24)) ;
    xnor2 L1_1_L2_3_G1_MINI_ALU_ix545 (.Y (L1_1_L2_3_G1_MINI_ALU_nx544), .A0 (
          L1SecondOperands_8__3), .A1 (L1FirstOperands_8__3)) ;
    xor2 L1_1_L2_3_G1_MINI_ALU_ix71 (.Y (L1Results_8__4), .A0 (
         L1_1_L2_3_G1_MINI_ALU_nx547), .A1 (L1_1_L2_3_G1_MINI_ALU_nx551)) ;
    aoi22 L1_1_L2_3_G1_MINI_ALU_ix548 (.Y (L1_1_L2_3_G1_MINI_ALU_nx547), .A0 (
          L1FirstOperands_8__3), .A1 (L1SecondOperands_8__3), .B0 (
          L1_1_L2_3_G1_MINI_ALU_nx44), .B1 (L1_1_L2_3_G1_MINI_ALU_nx18)) ;
    xnor2 L1_1_L2_3_G1_MINI_ALU_ix552 (.Y (L1_1_L2_3_G1_MINI_ALU_nx551), .A0 (
          L1SecondOperands_8__4), .A1 (L1FirstOperands_8__4)) ;
    xor2 L1_1_L2_3_G1_MINI_ALU_ix69 (.Y (L1Results_8__5), .A0 (
         L1_1_L2_3_G1_MINI_ALU_nx554), .A1 (L1_1_L2_3_G1_MINI_ALU_nx558)) ;
    aoi22 L1_1_L2_3_G1_MINI_ALU_ix555 (.Y (L1_1_L2_3_G1_MINI_ALU_nx554), .A0 (
          L1FirstOperands_8__4), .A1 (L1SecondOperands_8__4), .B0 (
          L1_1_L2_3_G1_MINI_ALU_nx48), .B1 (L1_1_L2_3_G1_MINI_ALU_nx12)) ;
    xnor2 L1_1_L2_3_G1_MINI_ALU_ix559 (.Y (L1_1_L2_3_G1_MINI_ALU_nx558), .A0 (
          L1SecondOperands_8__5), .A1 (L1FirstOperands_8__5)) ;
    xor2 L1_1_L2_3_G1_MINI_ALU_ix67 (.Y (L1Results_8__6), .A0 (
         L1_1_L2_3_G1_MINI_ALU_nx561), .A1 (L1_1_L2_3_G1_MINI_ALU_nx565)) ;
    aoi22 L1_1_L2_3_G1_MINI_ALU_ix562 (.Y (L1_1_L2_3_G1_MINI_ALU_nx561), .A0 (
          L1FirstOperands_8__5), .A1 (L1SecondOperands_8__5), .B0 (
          L1_1_L2_3_G1_MINI_ALU_nx52), .B1 (L1_1_L2_3_G1_MINI_ALU_nx6)) ;
    xnor2 L1_1_L2_3_G1_MINI_ALU_ix566 (.Y (L1_1_L2_3_G1_MINI_ALU_nx565), .A0 (
          L1SecondOperands_8__6), .A1 (L1FirstOperands_8__6)) ;
    xnor2 L1_1_L2_3_G1_MINI_ALU_ix65 (.Y (L1Results_8__7), .A0 (
          L1_1_L2_3_G1_MINI_ALU_nx568), .A1 (L1_1_L2_3_G1_MINI_ALU_nx62)) ;
    aoi22 L1_1_L2_3_G1_MINI_ALU_ix569 (.Y (L1_1_L2_3_G1_MINI_ALU_nx568), .A0 (
          L1FirstOperands_8__6), .A1 (L1SecondOperands_8__6), .B0 (
          L1_1_L2_3_G1_MINI_ALU_nx56), .B1 (L1_1_L2_3_G1_MINI_ALU_nx0)) ;
    xor2 L1_1_L2_3_G1_MINI_ALU_ix63 (.Y (L1_1_L2_3_G1_MINI_ALU_nx62), .A0 (
         L1SecondOperands_8__7), .A1 (L1FirstOperands_8__7)) ;
    inv01 L1_1_L2_3_G1_MINI_ALU_ix155 (.Y (L1_1_L2_3_G1_MINI_ALU_nx154), .A (
          L1_1_L2_3_G1_MINI_ALU_nx383)) ;
    inv01 L1_1_L2_3_G1_MINI_ALU_ix57 (.Y (L1_1_L2_3_G1_MINI_ALU_nx56), .A (
          L1_1_L2_3_G1_MINI_ALU_nx561)) ;
    inv01 L1_1_L2_3_G1_MINI_ALU_ix53 (.Y (L1_1_L2_3_G1_MINI_ALU_nx52), .A (
          L1_1_L2_3_G1_MINI_ALU_nx554)) ;
    inv01 L1_1_L2_3_G1_MINI_ALU_ix49 (.Y (L1_1_L2_3_G1_MINI_ALU_nx48), .A (
          L1_1_L2_3_G1_MINI_ALU_nx547)) ;
    inv01 L1_1_L2_3_G1_MINI_ALU_ix45 (.Y (L1_1_L2_3_G1_MINI_ALU_nx44), .A (
          L1_1_L2_3_G1_MINI_ALU_nx540)) ;
    inv01 L1_1_L2_3_G1_MINI_ALU_ix41 (.Y (L1_1_L2_3_G1_MINI_ALU_nx40), .A (
          L1_1_L2_3_G1_MINI_ALU_nx534)) ;
    inv01 L1_1_L2_3_G1_MINI_ALU_ix31 (.Y (L1_1_L2_3_G1_MINI_ALU_nx30), .A (
          L1_1_L2_3_G1_MINI_ALU_nx531)) ;
    inv01 L1_1_L2_3_G1_MINI_ALU_ix25 (.Y (L1_1_L2_3_G1_MINI_ALU_nx24), .A (
          L1_1_L2_3_G1_MINI_ALU_nx537)) ;
    inv01 L1_1_L2_3_G1_MINI_ALU_ix19 (.Y (L1_1_L2_3_G1_MINI_ALU_nx18), .A (
          L1_1_L2_3_G1_MINI_ALU_nx544)) ;
    inv01 L1_1_L2_3_G1_MINI_ALU_ix13 (.Y (L1_1_L2_3_G1_MINI_ALU_nx12), .A (
          L1_1_L2_3_G1_MINI_ALU_nx551)) ;
    inv01 L1_1_L2_3_G1_MINI_ALU_ix7 (.Y (L1_1_L2_3_G1_MINI_ALU_nx6), .A (
          L1_1_L2_3_G1_MINI_ALU_nx558)) ;
    inv01 L1_1_L2_3_G1_MINI_ALU_ix1 (.Y (L1_1_L2_3_G1_MINI_ALU_nx0), .A (
          L1_1_L2_3_G1_MINI_ALU_nx565)) ;
    fake_gnd L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix216 (.Y (
             L1_1_L2_3_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    nor02ii L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix81 (.Y (
            L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx80), .A0 (Instr), .A1 (Start)) ;
    aoi21 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix77 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_10), .A0 (
          FilterDin_1__3__1), .A1 (FilterDin_1__3__0), .B0 (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx4)) ;
    nor02_2x L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix5 (.Y (
             L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx4), .A0 (FilterDin_1__3__0), .A1 (
             FilterDin_1__3__1)) ;
    aoi21 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix67 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_11), .A0 (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx328), .A1 (FilterDin_1__3__2), .B0 (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx8)) ;
    nor03_2x L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix9 (.Y (
             L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx8), .A0 (FilterDin_1__3__2), .A1 (
             FilterDin_1__3__0), .A2 (FilterDin_1__3__1)) ;
    xnor2 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix59 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_12), .A0 (
          FilterDin_1__3__3), .A1 (L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx8)) ;
    xnor2 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix51 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_13), .A0 (
          FilterDin_1__3__4), .A1 (L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx12)) ;
    nor04 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix13 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx12), .A0 (FilterDin_1__3__3), .A1 (
          FilterDin_1__3__2), .A2 (FilterDin_1__3__0), .A3 (FilterDin_1__3__1)
          ) ;
    xnor2 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix43 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_14), .A0 (
          FilterDin_1__3__5), .A1 (L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx16)) ;
    nor02ii L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix17 (.Y (
            L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx16), .A0 (FilterDin_1__3__4), .A1 (
            L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx12)) ;
    xnor2 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix35 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_15), .A0 (
          FilterDin_1__3__6), .A1 (L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx20)) ;
    nor02ii L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix21 (.Y (
            L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx20), .A0 (FilterDin_1__3__5), .A1 (
            L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx16)) ;
    xnor2 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix27 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_16), .A0 (
          FilterDin_1__3__7), .A1 (L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx24)) ;
    nor02ii L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix25 (.Y (
            L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx24), .A0 (FilterDin_1__3__6), .A1 (
            L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx20)) ;
    inv01 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix329 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx328), .A (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx4)) ;
    inv02 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix383 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx384), .A (
          L1_1_L2_3_G1_MINI_ALU_BoothP_0)) ;
    dff L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_0 (.Q (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_0), .QB (\$dummy [412]), 
        .D (L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .CLK (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    nor02_2x L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix567 (.Y (
             L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566), .A0 (RST), .A1 (
             L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644)) ;
    dff L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_1 (.Q (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_1), .QB (\$dummy [413]), 
        .D (L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .CLK (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_2 (.Q (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_2), .QB (\$dummy [414]), 
        .D (L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .CLK (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_3 (.Q (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_3), .QB (\$dummy [415]), 
        .D (L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .CLK (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_4 (.Q (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_4), .QB (\$dummy [416]), 
        .D (L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .CLK (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_5 (.Q (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_5), .QB (\$dummy [417]), 
        .D (L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .CLK (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_6 (.Q (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_6), .QB (\$dummy [418]), 
        .D (L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .CLK (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_7 (.Q (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_7), .QB (\$dummy [419]), 
        .D (L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .CLK (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_8 (.Q (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_8), .QB (\$dummy [420]), 
        .D (L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .CLK (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_9 (.Q (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_9), .QB (\$dummy [421]), 
        .D (L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .CLK (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_10 (.Q (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_10), .QB (\$dummy [422])
        , .D (L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .CLK (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_11 (.Q (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_11), .QB (\$dummy [423])
        , .D (L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .CLK (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_12 (.Q (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_12), .QB (\$dummy [424])
        , .D (L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .CLK (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_13 (.Q (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_13), .QB (\$dummy [425])
        , .D (L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .CLK (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_14 (.Q (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_14), .QB (\$dummy [426])
        , .D (L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .CLK (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_15 (.Q (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_15), .QB (\$dummy [427])
        , .D (L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .CLK (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_16 (.Q (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_16), .QB (\$dummy [428])
        , .D (L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .CLK (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    inv02 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix623 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624), .A (CLK)) ;
    inv02 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix625 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626), .A (CLK)) ;
    inv02 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix627 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628), .A (CLK)) ;
    inv02 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix643 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644), .A (nx7938)) ;
    dff L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_0 (.Q (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_0), .QB (\$dummy [429]), 
        .D (L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .CLK (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    nor02_2x L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix567 (.Y (
             L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566), .A0 (RST), .A1 (
             L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644)) ;
    dff L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_1 (.Q (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_1), .QB (\$dummy [430]), 
        .D (L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .CLK (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_2 (.Q (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_2), .QB (\$dummy [431]), 
        .D (L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .CLK (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_3 (.Q (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_3), .QB (\$dummy [432]), 
        .D (L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .CLK (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_4 (.Q (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_4), .QB (\$dummy [433]), 
        .D (L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .CLK (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_5 (.Q (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_5), .QB (\$dummy [434]), 
        .D (L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .CLK (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_6 (.Q (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_6), .QB (\$dummy [435]), 
        .D (L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .CLK (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_7 (.Q (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_7), .QB (\$dummy [436]), 
        .D (L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .CLK (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_8 (.Q (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_8), .QB (\$dummy [437]), 
        .D (L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .CLK (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_9 (.Q (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_9), .QB (\$dummy [438]), 
        .D (L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .CLK (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_10 (.Q (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_10), .QB (\$dummy [439])
        , .D (L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .CLK (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_11 (.Q (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_11), .QB (\$dummy [440])
        , .D (L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .CLK (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_12 (.Q (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_12), .QB (\$dummy [441])
        , .D (L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .CLK (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_13 (.Q (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_13), .QB (\$dummy [442])
        , .D (L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .CLK (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_14 (.Q (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_14), .QB (\$dummy [443])
        , .D (L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .CLK (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_15 (.Q (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_15), .QB (\$dummy [444])
        , .D (L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .CLK (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_16 (.Q (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_16), .QB (\$dummy [445])
        , .D (L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .CLK (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    inv02 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix623 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624), .A (CLK)) ;
    inv02 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix625 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626), .A (CLK)) ;
    inv02 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix627 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628), .A (CLK)) ;
    inv02 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix643 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644), .A (nx7944)) ;
    dff L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_0 (.Q (
        L1_1_L2_3_G1_MINI_ALU_BoothP_0), .QB (\$dummy [446]), .D (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .CLK (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    nor02_2x L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix567 (.Y (
             L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566), .A0 (RST), .A1 (
             L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    dff L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_1 (.Q (
        L1_1_L2_3_G1_MINI_ALU_BoothP_1), .QB (\$dummy [447]), .D (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .CLK (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_2 (.Q (
        L1_1_L2_3_G1_MINI_ALU_BoothP_2), .QB (\$dummy [448]), .D (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .CLK (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_3 (.Q (
        L1_1_L2_3_G1_MINI_ALU_BoothP_3), .QB (\$dummy [449]), .D (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .CLK (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_4 (.Q (
        L1_1_L2_3_G1_MINI_ALU_BoothP_4), .QB (\$dummy [450]), .D (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .CLK (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_5 (.Q (
        L1_1_L2_3_G1_MINI_ALU_BoothP_5), .QB (\$dummy [451]), .D (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .CLK (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_6 (.Q (
        L1_1_L2_3_G1_MINI_ALU_BoothP_6), .QB (\$dummy [452]), .D (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .CLK (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_7 (.Q (
        L1_1_L2_3_G1_MINI_ALU_BoothP_7), .QB (\$dummy [453]), .D (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .CLK (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_8 (.Q (
        L1_1_L2_3_G1_MINI_ALU_BoothP_8), .QB (\$dummy [454]), .D (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .CLK (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_9 (.Q (
        L1_1_L2_3_G1_MINI_ALU_BoothP_9), .QB (\$dummy [455]), .D (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .CLK (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_10 (.Q (
        L1_1_L2_3_G1_MINI_ALU_BoothP_10), .QB (\$dummy [456]), .D (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .CLK (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_11 (.Q (
        L1_1_L2_3_G1_MINI_ALU_BoothP_11), .QB (\$dummy [457]), .D (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .CLK (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_12 (.Q (
        L1_1_L2_3_G1_MINI_ALU_BoothP_12), .QB (\$dummy [458]), .D (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .CLK (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_13 (.Q (
        L1_1_L2_3_G1_MINI_ALU_BoothP_13), .QB (\$dummy [459]), .D (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .CLK (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_14 (.Q (
        L1_1_L2_3_G1_MINI_ALU_BoothP_14), .QB (\$dummy [460]), .D (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .CLK (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_15 (.Q (
        L1_1_L2_3_G1_MINI_ALU_BoothP_15), .QB (\$dummy [461]), .D (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .CLK (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_16 (.Q (
        L1_1_L2_3_G1_MINI_ALU_BoothP_16), .QB (\$dummy [462]), .D (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .CLK (
        L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    inv02 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix623 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624), .A (CLK)) ;
    inv02 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix625 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626), .A (CLK)) ;
    inv02 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix627 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628), .A (CLK)) ;
    inv02 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix643 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644), .A (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642)) ;
    xor2 L1_1_L2_4_G1_MINI_ALU_ix83 (.Y (L1Results_9__0), .A0 (
         L1SecondOperands_9__0), .A1 (L1FirstOperands_9__0)) ;
    xnor2 L1_1_L2_4_G1_MINI_ALU_ix380 (.Y (L1_1_L2_4_G1_MINI_ALU_nx379), .A0 (
          L1_1_L2_4_G1_MINI_ALU_nx381), .A1 (L1_1_L2_4_G1_MINI_ALU_nx383)) ;
    nand02 L1_1_L2_4_G1_MINI_ALU_ix382 (.Y (L1_1_L2_4_G1_MINI_ALU_nx381), .A0 (
           L1_1_L2_4_G1_MINI_ALU_BoothOperand_0), .A1 (nx7964)) ;
    xnor2 L1_1_L2_4_G1_MINI_ALU_ix384 (.Y (L1_1_L2_4_G1_MINI_ALU_nx383), .A0 (
          L1_1_L2_4_G1_MINI_ALU_BoothOperand_1), .A1 (
          L1_1_L2_4_G1_MINI_ALU_BoothP_1)) ;
    inv01 L1_1_L2_4_G1_MINI_ALU_ix388 (.Y (L1_1_L2_4_G1_MINI_ALU_nx387), .A (
          L1_1_L2_4_G1_MINI_ALU_BoothP_2)) ;
    xnor2 L1_1_L2_4_G1_MINI_ALU_ix390 (.Y (L1_1_L2_4_G1_MINI_ALU_nx389), .A0 (
          L1_1_L2_4_G1_MINI_ALU_nx391), .A1 (L1_1_L2_4_G1_MINI_ALU_nx395)) ;
    aoi32 L1_1_L2_4_G1_MINI_ALU_ix392 (.Y (L1_1_L2_4_G1_MINI_ALU_nx391), .A0 (
          L1_1_L2_4_G1_MINI_ALU_BoothOperand_0), .A1 (nx7964), .A2 (
          L1_1_L2_4_G1_MINI_ALU_nx154), .B0 (L1_1_L2_4_G1_MINI_ALU_BoothP_1), .B1 (
          L1_1_L2_4_G1_MINI_ALU_BoothOperand_1)) ;
    xnor2 L1_1_L2_4_G1_MINI_ALU_ix396 (.Y (L1_1_L2_4_G1_MINI_ALU_nx395), .A0 (
          L1_1_L2_4_G1_MINI_ALU_BoothOperand_2), .A1 (
          L1_1_L2_4_G1_MINI_ALU_BoothP_2)) ;
    inv01 L1_1_L2_4_G1_MINI_ALU_ix400 (.Y (L1_1_L2_4_G1_MINI_ALU_nx399), .A (
          L1_1_L2_4_G1_MINI_ALU_BoothP_3)) ;
    xnor2 L1_1_L2_4_G1_MINI_ALU_ix402 (.Y (L1_1_L2_4_G1_MINI_ALU_nx401), .A0 (
          L1_1_L2_4_G1_MINI_ALU_nx403), .A1 (L1_1_L2_4_G1_MINI_ALU_nx405)) ;
    xnor2 L1_1_L2_4_G1_MINI_ALU_ix406 (.Y (L1_1_L2_4_G1_MINI_ALU_nx405), .A0 (
          L1_1_L2_4_G1_MINI_ALU_BoothOperand_3), .A1 (
          L1_1_L2_4_G1_MINI_ALU_BoothP_3)) ;
    inv01 L1_1_L2_4_G1_MINI_ALU_ix410 (.Y (L1_1_L2_4_G1_MINI_ALU_nx409), .A (
          L1_1_L2_4_G1_MINI_ALU_BoothP_4)) ;
    xnor2 L1_1_L2_4_G1_MINI_ALU_ix412 (.Y (L1_1_L2_4_G1_MINI_ALU_nx411), .A0 (
          L1_1_L2_4_G1_MINI_ALU_nx413), .A1 (L1_1_L2_4_G1_MINI_ALU_nx415)) ;
    xnor2 L1_1_L2_4_G1_MINI_ALU_ix416 (.Y (L1_1_L2_4_G1_MINI_ALU_nx415), .A0 (
          L1_1_L2_4_G1_MINI_ALU_BoothOperand_4), .A1 (
          L1_1_L2_4_G1_MINI_ALU_BoothP_4)) ;
    inv01 L1_1_L2_4_G1_MINI_ALU_ix420 (.Y (L1_1_L2_4_G1_MINI_ALU_nx419), .A (
          L1_1_L2_4_G1_MINI_ALU_BoothP_5)) ;
    xnor2 L1_1_L2_4_G1_MINI_ALU_ix422 (.Y (L1_1_L2_4_G1_MINI_ALU_nx421), .A0 (
          L1_1_L2_4_G1_MINI_ALU_nx423), .A1 (L1_1_L2_4_G1_MINI_ALU_nx425)) ;
    xnor2 L1_1_L2_4_G1_MINI_ALU_ix426 (.Y (L1_1_L2_4_G1_MINI_ALU_nx425), .A0 (
          L1_1_L2_4_G1_MINI_ALU_BoothOperand_5), .A1 (
          L1_1_L2_4_G1_MINI_ALU_BoothP_5)) ;
    inv01 L1_1_L2_4_G1_MINI_ALU_ix430 (.Y (L1_1_L2_4_G1_MINI_ALU_nx429), .A (
          L1_1_L2_4_G1_MINI_ALU_BoothP_6)) ;
    xnor2 L1_1_L2_4_G1_MINI_ALU_ix432 (.Y (L1_1_L2_4_G1_MINI_ALU_nx431), .A0 (
          L1_1_L2_4_G1_MINI_ALU_nx433), .A1 (L1_1_L2_4_G1_MINI_ALU_nx435)) ;
    xnor2 L1_1_L2_4_G1_MINI_ALU_ix436 (.Y (L1_1_L2_4_G1_MINI_ALU_nx435), .A0 (
          L1_1_L2_4_G1_MINI_ALU_BoothOperand_6), .A1 (
          L1_1_L2_4_G1_MINI_ALU_BoothP_6)) ;
    inv01 L1_1_L2_4_G1_MINI_ALU_ix440 (.Y (L1_1_L2_4_G1_MINI_ALU_nx439), .A (
          L1_1_L2_4_G1_MINI_ALU_BoothP_7)) ;
    xnor2 L1_1_L2_4_G1_MINI_ALU_ix442 (.Y (L1_1_L2_4_G1_MINI_ALU_nx441), .A0 (
          L1_1_L2_4_G1_MINI_ALU_nx443), .A1 (L1_1_L2_4_G1_MINI_ALU_nx445)) ;
    xnor2 L1_1_L2_4_G1_MINI_ALU_ix446 (.Y (L1_1_L2_4_G1_MINI_ALU_nx445), .A0 (
          L1_1_L2_4_G1_MINI_ALU_BoothOperand_7), .A1 (
          L1_1_L2_4_G1_MINI_ALU_BoothP_7)) ;
    inv01 L1_1_L2_4_G1_MINI_ALU_ix450 (.Y (L1_1_L2_4_G1_MINI_ALU_nx449), .A (
          L1_1_L2_4_G1_MINI_ALU_BoothP_8)) ;
    xnor2 L1_1_L2_4_G1_MINI_ALU_ix452 (.Y (L1_1_L2_4_G1_MINI_ALU_nx451), .A0 (
          L1_1_L2_4_G1_MINI_ALU_nx453), .A1 (L1_1_L2_4_G1_MINI_ALU_nx455)) ;
    xnor2 L1_1_L2_4_G1_MINI_ALU_ix456 (.Y (L1_1_L2_4_G1_MINI_ALU_nx455), .A0 (
          L1_1_L2_4_G1_MINI_ALU_BoothOperand_8), .A1 (
          L1_1_L2_4_G1_MINI_ALU_BoothP_8)) ;
    xor2 L1_1_L2_4_G1_MINI_ALU_ix317 (.Y (L1_1_L2_4_G1_MINI_ALU_nx316), .A0 (
         L1_1_L2_4_G1_MINI_ALU_nx461), .A1 (L1_1_L2_4_G1_MINI_ALU_nx463)) ;
    xnor2 L1_1_L2_4_G1_MINI_ALU_ix464 (.Y (L1_1_L2_4_G1_MINI_ALU_nx463), .A0 (
          L1_1_L2_4_G1_MINI_ALU_BoothOperand_9), .A1 (
          L1_1_L2_4_G1_MINI_ALU_BoothP_9)) ;
    xor2 L1_1_L2_4_G1_MINI_ALU_ix337 (.Y (L1_1_L2_4_G1_MINI_ALU_nx336), .A0 (
         L1_1_L2_4_G1_MINI_ALU_nx467), .A1 (L1_1_L2_4_G1_MINI_ALU_nx471)) ;
    inv01 L1_1_L2_4_G1_MINI_ALU_ix470 (.Y (L1_1_L2_4_G1_MINI_ALU_nx469), .A (
          L1_1_L2_4_G1_MINI_ALU_BoothP_9)) ;
    xnor2 L1_1_L2_4_G1_MINI_ALU_ix472 (.Y (L1_1_L2_4_G1_MINI_ALU_nx471), .A0 (
          L1_1_L2_4_G1_MINI_ALU_BoothOperand_10), .A1 (
          L1_1_L2_4_G1_MINI_ALU_BoothP_10)) ;
    xor2 L1_1_L2_4_G1_MINI_ALU_ix357 (.Y (L1_1_L2_4_G1_MINI_ALU_nx356), .A0 (
         L1_1_L2_4_G1_MINI_ALU_nx475), .A1 (L1_1_L2_4_G1_MINI_ALU_nx479)) ;
    inv01 L1_1_L2_4_G1_MINI_ALU_ix478 (.Y (L1_1_L2_4_G1_MINI_ALU_nx477), .A (
          L1_1_L2_4_G1_MINI_ALU_BoothP_10)) ;
    xnor2 L1_1_L2_4_G1_MINI_ALU_ix480 (.Y (L1_1_L2_4_G1_MINI_ALU_nx479), .A0 (
          L1_1_L2_4_G1_MINI_ALU_BoothOperand_11), .A1 (
          L1_1_L2_4_G1_MINI_ALU_BoothP_11)) ;
    xor2 L1_1_L2_4_G1_MINI_ALU_ix377 (.Y (L1_1_L2_4_G1_MINI_ALU_nx376), .A0 (
         L1_1_L2_4_G1_MINI_ALU_nx483), .A1 (L1_1_L2_4_G1_MINI_ALU_nx487)) ;
    inv01 L1_1_L2_4_G1_MINI_ALU_ix486 (.Y (L1_1_L2_4_G1_MINI_ALU_nx485), .A (
          L1_1_L2_4_G1_MINI_ALU_BoothP_11)) ;
    xnor2 L1_1_L2_4_G1_MINI_ALU_ix488 (.Y (L1_1_L2_4_G1_MINI_ALU_nx487), .A0 (
          L1_1_L2_4_G1_MINI_ALU_BoothOperand_12), .A1 (
          L1_1_L2_4_G1_MINI_ALU_BoothP_12)) ;
    xor2 L1_1_L2_4_G1_MINI_ALU_ix397 (.Y (L1_1_L2_4_G1_MINI_ALU_nx396), .A0 (
         L1_1_L2_4_G1_MINI_ALU_nx491), .A1 (L1_1_L2_4_G1_MINI_ALU_nx495)) ;
    inv01 L1_1_L2_4_G1_MINI_ALU_ix494 (.Y (L1_1_L2_4_G1_MINI_ALU_nx493), .A (
          L1_1_L2_4_G1_MINI_ALU_BoothP_12)) ;
    xnor2 L1_1_L2_4_G1_MINI_ALU_ix496 (.Y (L1_1_L2_4_G1_MINI_ALU_nx495), .A0 (
          L1_1_L2_4_G1_MINI_ALU_BoothOperand_13), .A1 (
          L1_1_L2_4_G1_MINI_ALU_BoothP_13)) ;
    xor2 L1_1_L2_4_G1_MINI_ALU_ix417 (.Y (L1_1_L2_4_G1_MINI_ALU_nx416), .A0 (
         L1_1_L2_4_G1_MINI_ALU_nx499), .A1 (L1_1_L2_4_G1_MINI_ALU_nx503)) ;
    inv01 L1_1_L2_4_G1_MINI_ALU_ix502 (.Y (L1_1_L2_4_G1_MINI_ALU_nx501), .A (
          L1_1_L2_4_G1_MINI_ALU_BoothP_13)) ;
    xnor2 L1_1_L2_4_G1_MINI_ALU_ix504 (.Y (L1_1_L2_4_G1_MINI_ALU_nx503), .A0 (
          L1_1_L2_4_G1_MINI_ALU_BoothOperand_14), .A1 (
          L1_1_L2_4_G1_MINI_ALU_BoothP_14)) ;
    xor2 L1_1_L2_4_G1_MINI_ALU_ix437 (.Y (L1_1_L2_4_G1_MINI_ALU_nx436), .A0 (
         L1_1_L2_4_G1_MINI_ALU_nx507), .A1 (L1_1_L2_4_G1_MINI_ALU_nx511)) ;
    inv01 L1_1_L2_4_G1_MINI_ALU_ix510 (.Y (L1_1_L2_4_G1_MINI_ALU_nx509), .A (
          L1_1_L2_4_G1_MINI_ALU_BoothP_14)) ;
    xnor2 L1_1_L2_4_G1_MINI_ALU_ix512 (.Y (L1_1_L2_4_G1_MINI_ALU_nx511), .A0 (
          L1_1_L2_4_G1_MINI_ALU_BoothOperand_15), .A1 (
          L1_1_L2_4_G1_MINI_ALU_BoothP_15)) ;
    xnor2 L1_1_L2_4_G1_MINI_ALU_ix457 (.Y (L1_1_L2_4_G1_MINI_ALU_nx456), .A0 (
          L1_1_L2_4_G1_MINI_ALU_nx515), .A1 (L1_1_L2_4_G1_MINI_ALU_nx454)) ;
    inv01 L1_1_L2_4_G1_MINI_ALU_ix518 (.Y (L1_1_L2_4_G1_MINI_ALU_nx517), .A (
          L1_1_L2_4_G1_MINI_ALU_BoothP_15)) ;
    xor2 L1_1_L2_4_G1_MINI_ALU_ix455 (.Y (L1_1_L2_4_G1_MINI_ALU_nx454), .A0 (
         L1_1_L2_4_G1_MINI_ALU_BoothOperand_16), .A1 (
         L1_1_L2_4_G1_MINI_ALU_BoothP_16)) ;
    mux21_ni L1_1_L2_4_G1_MINI_ALU_ix91 (.Y (L1SecondOperands_9__0), .A0 (
             L1_1_L2_4_G1_MINI_ALU_BoothP_1), .A1 (WindowDin_1__4__0), .S0 (
             Instr)) ;
    mux21_ni L1_1_L2_4_G1_MINI_ALU_ix99 (.Y (L1SecondOperands_9__1), .A0 (
             L1_1_L2_4_G1_MINI_ALU_BoothP_2), .A1 (WindowDin_1__4__1), .S0 (
             Instr)) ;
    mux21_ni L1_1_L2_4_G1_MINI_ALU_ix107 (.Y (L1SecondOperands_9__2), .A0 (
             L1_1_L2_4_G1_MINI_ALU_BoothP_3), .A1 (WindowDin_1__4__2), .S0 (
             Instr)) ;
    mux21_ni L1_1_L2_4_G1_MINI_ALU_ix115 (.Y (L1SecondOperands_9__3), .A0 (
             L1_1_L2_4_G1_MINI_ALU_BoothP_4), .A1 (WindowDin_1__4__3), .S0 (
             Instr)) ;
    mux21_ni L1_1_L2_4_G1_MINI_ALU_ix123 (.Y (L1SecondOperands_9__4), .A0 (
             L1_1_L2_4_G1_MINI_ALU_BoothP_5), .A1 (WindowDin_1__4__4), .S0 (
             Instr)) ;
    mux21_ni L1_1_L2_4_G1_MINI_ALU_ix131 (.Y (L1SecondOperands_9__5), .A0 (
             L1_1_L2_4_G1_MINI_ALU_BoothP_6), .A1 (WindowDin_1__4__5), .S0 (
             Instr)) ;
    mux21_ni L1_1_L2_4_G1_MINI_ALU_ix139 (.Y (L1SecondOperands_9__6), .A0 (
             L1_1_L2_4_G1_MINI_ALU_BoothP_7), .A1 (WindowDin_1__4__6), .S0 (
             Instr)) ;
    mux21_ni L1_1_L2_4_G1_MINI_ALU_ix147 (.Y (L1SecondOperands_9__7), .A0 (
             L1_1_L2_4_G1_MINI_ALU_BoothP_8), .A1 (WindowDin_1__4__7), .S0 (
             Instr)) ;
    xor2 L1_1_L2_4_G1_MINI_ALU_ix77 (.Y (L1Results_9__1), .A0 (
         L1_1_L2_4_G1_MINI_ALU_nx529), .A1 (L1_1_L2_4_G1_MINI_ALU_nx531)) ;
    nand02 L1_1_L2_4_G1_MINI_ALU_ix530 (.Y (L1_1_L2_4_G1_MINI_ALU_nx529), .A0 (
           L1SecondOperands_9__0), .A1 (L1FirstOperands_9__0)) ;
    xnor2 L1_1_L2_4_G1_MINI_ALU_ix532 (.Y (L1_1_L2_4_G1_MINI_ALU_nx531), .A0 (
          L1SecondOperands_9__1), .A1 (L1FirstOperands_9__1)) ;
    xor2 L1_1_L2_4_G1_MINI_ALU_ix75 (.Y (L1Results_9__2), .A0 (
         L1_1_L2_4_G1_MINI_ALU_nx534), .A1 (L1_1_L2_4_G1_MINI_ALU_nx537)) ;
    aoi32 L1_1_L2_4_G1_MINI_ALU_ix535 (.Y (L1_1_L2_4_G1_MINI_ALU_nx534), .A0 (
          L1SecondOperands_9__0), .A1 (L1FirstOperands_9__0), .A2 (
          L1_1_L2_4_G1_MINI_ALU_nx30), .B0 (L1FirstOperands_9__1), .B1 (
          L1SecondOperands_9__1)) ;
    xnor2 L1_1_L2_4_G1_MINI_ALU_ix538 (.Y (L1_1_L2_4_G1_MINI_ALU_nx537), .A0 (
          L1SecondOperands_9__2), .A1 (L1FirstOperands_9__2)) ;
    xor2 L1_1_L2_4_G1_MINI_ALU_ix73 (.Y (L1Results_9__3), .A0 (
         L1_1_L2_4_G1_MINI_ALU_nx540), .A1 (L1_1_L2_4_G1_MINI_ALU_nx544)) ;
    aoi22 L1_1_L2_4_G1_MINI_ALU_ix541 (.Y (L1_1_L2_4_G1_MINI_ALU_nx540), .A0 (
          L1FirstOperands_9__2), .A1 (L1SecondOperands_9__2), .B0 (
          L1_1_L2_4_G1_MINI_ALU_nx40), .B1 (L1_1_L2_4_G1_MINI_ALU_nx24)) ;
    xnor2 L1_1_L2_4_G1_MINI_ALU_ix545 (.Y (L1_1_L2_4_G1_MINI_ALU_nx544), .A0 (
          L1SecondOperands_9__3), .A1 (L1FirstOperands_9__3)) ;
    xor2 L1_1_L2_4_G1_MINI_ALU_ix71 (.Y (L1Results_9__4), .A0 (
         L1_1_L2_4_G1_MINI_ALU_nx547), .A1 (L1_1_L2_4_G1_MINI_ALU_nx551)) ;
    aoi22 L1_1_L2_4_G1_MINI_ALU_ix548 (.Y (L1_1_L2_4_G1_MINI_ALU_nx547), .A0 (
          L1FirstOperands_9__3), .A1 (L1SecondOperands_9__3), .B0 (
          L1_1_L2_4_G1_MINI_ALU_nx44), .B1 (L1_1_L2_4_G1_MINI_ALU_nx18)) ;
    xnor2 L1_1_L2_4_G1_MINI_ALU_ix552 (.Y (L1_1_L2_4_G1_MINI_ALU_nx551), .A0 (
          L1SecondOperands_9__4), .A1 (L1FirstOperands_9__4)) ;
    xor2 L1_1_L2_4_G1_MINI_ALU_ix69 (.Y (L1Results_9__5), .A0 (
         L1_1_L2_4_G1_MINI_ALU_nx554), .A1 (L1_1_L2_4_G1_MINI_ALU_nx558)) ;
    aoi22 L1_1_L2_4_G1_MINI_ALU_ix555 (.Y (L1_1_L2_4_G1_MINI_ALU_nx554), .A0 (
          L1FirstOperands_9__4), .A1 (L1SecondOperands_9__4), .B0 (
          L1_1_L2_4_G1_MINI_ALU_nx48), .B1 (L1_1_L2_4_G1_MINI_ALU_nx12)) ;
    xnor2 L1_1_L2_4_G1_MINI_ALU_ix559 (.Y (L1_1_L2_4_G1_MINI_ALU_nx558), .A0 (
          L1SecondOperands_9__5), .A1 (L1FirstOperands_9__5)) ;
    xor2 L1_1_L2_4_G1_MINI_ALU_ix67 (.Y (L1Results_9__6), .A0 (
         L1_1_L2_4_G1_MINI_ALU_nx561), .A1 (L1_1_L2_4_G1_MINI_ALU_nx565)) ;
    aoi22 L1_1_L2_4_G1_MINI_ALU_ix562 (.Y (L1_1_L2_4_G1_MINI_ALU_nx561), .A0 (
          L1FirstOperands_9__5), .A1 (L1SecondOperands_9__5), .B0 (
          L1_1_L2_4_G1_MINI_ALU_nx52), .B1 (L1_1_L2_4_G1_MINI_ALU_nx6)) ;
    xnor2 L1_1_L2_4_G1_MINI_ALU_ix566 (.Y (L1_1_L2_4_G1_MINI_ALU_nx565), .A0 (
          L1SecondOperands_9__6), .A1 (L1FirstOperands_9__6)) ;
    xnor2 L1_1_L2_4_G1_MINI_ALU_ix65 (.Y (L1Results_9__7), .A0 (
          L1_1_L2_4_G1_MINI_ALU_nx568), .A1 (L1_1_L2_4_G1_MINI_ALU_nx62)) ;
    aoi22 L1_1_L2_4_G1_MINI_ALU_ix569 (.Y (L1_1_L2_4_G1_MINI_ALU_nx568), .A0 (
          L1FirstOperands_9__6), .A1 (L1SecondOperands_9__6), .B0 (
          L1_1_L2_4_G1_MINI_ALU_nx56), .B1 (L1_1_L2_4_G1_MINI_ALU_nx0)) ;
    xor2 L1_1_L2_4_G1_MINI_ALU_ix63 (.Y (L1_1_L2_4_G1_MINI_ALU_nx62), .A0 (
         L1SecondOperands_9__7), .A1 (L1FirstOperands_9__7)) ;
    inv01 L1_1_L2_4_G1_MINI_ALU_ix155 (.Y (L1_1_L2_4_G1_MINI_ALU_nx154), .A (
          L1_1_L2_4_G1_MINI_ALU_nx383)) ;
    inv01 L1_1_L2_4_G1_MINI_ALU_ix57 (.Y (L1_1_L2_4_G1_MINI_ALU_nx56), .A (
          L1_1_L2_4_G1_MINI_ALU_nx561)) ;
    inv01 L1_1_L2_4_G1_MINI_ALU_ix53 (.Y (L1_1_L2_4_G1_MINI_ALU_nx52), .A (
          L1_1_L2_4_G1_MINI_ALU_nx554)) ;
    inv01 L1_1_L2_4_G1_MINI_ALU_ix49 (.Y (L1_1_L2_4_G1_MINI_ALU_nx48), .A (
          L1_1_L2_4_G1_MINI_ALU_nx547)) ;
    inv01 L1_1_L2_4_G1_MINI_ALU_ix45 (.Y (L1_1_L2_4_G1_MINI_ALU_nx44), .A (
          L1_1_L2_4_G1_MINI_ALU_nx540)) ;
    inv01 L1_1_L2_4_G1_MINI_ALU_ix41 (.Y (L1_1_L2_4_G1_MINI_ALU_nx40), .A (
          L1_1_L2_4_G1_MINI_ALU_nx534)) ;
    inv01 L1_1_L2_4_G1_MINI_ALU_ix31 (.Y (L1_1_L2_4_G1_MINI_ALU_nx30), .A (
          L1_1_L2_4_G1_MINI_ALU_nx531)) ;
    inv01 L1_1_L2_4_G1_MINI_ALU_ix25 (.Y (L1_1_L2_4_G1_MINI_ALU_nx24), .A (
          L1_1_L2_4_G1_MINI_ALU_nx537)) ;
    inv01 L1_1_L2_4_G1_MINI_ALU_ix19 (.Y (L1_1_L2_4_G1_MINI_ALU_nx18), .A (
          L1_1_L2_4_G1_MINI_ALU_nx544)) ;
    inv01 L1_1_L2_4_G1_MINI_ALU_ix13 (.Y (L1_1_L2_4_G1_MINI_ALU_nx12), .A (
          L1_1_L2_4_G1_MINI_ALU_nx551)) ;
    inv01 L1_1_L2_4_G1_MINI_ALU_ix7 (.Y (L1_1_L2_4_G1_MINI_ALU_nx6), .A (
          L1_1_L2_4_G1_MINI_ALU_nx558)) ;
    inv01 L1_1_L2_4_G1_MINI_ALU_ix1 (.Y (L1_1_L2_4_G1_MINI_ALU_nx0), .A (
          L1_1_L2_4_G1_MINI_ALU_nx565)) ;
    fake_gnd L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix216 (.Y (
             L1_1_L2_4_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    nor02ii L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix81 (.Y (
            L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx80), .A0 (Instr), .A1 (Start)) ;
    aoi21 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix77 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_10), .A0 (
          FilterDin_1__4__1), .A1 (FilterDin_1__4__0), .B0 (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx4)) ;
    nor02_2x L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix5 (.Y (
             L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx4), .A0 (FilterDin_1__4__0), .A1 (
             FilterDin_1__4__1)) ;
    aoi21 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix67 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_11), .A0 (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx328), .A1 (FilterDin_1__4__2), .B0 (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx8)) ;
    nor03_2x L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix9 (.Y (
             L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx8), .A0 (FilterDin_1__4__2), .A1 (
             FilterDin_1__4__0), .A2 (FilterDin_1__4__1)) ;
    xnor2 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix59 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_12), .A0 (
          FilterDin_1__4__3), .A1 (L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx8)) ;
    xnor2 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix51 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_13), .A0 (
          FilterDin_1__4__4), .A1 (L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx12)) ;
    nor04 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix13 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx12), .A0 (FilterDin_1__4__3), .A1 (
          FilterDin_1__4__2), .A2 (FilterDin_1__4__0), .A3 (FilterDin_1__4__1)
          ) ;
    xnor2 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix43 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_14), .A0 (
          FilterDin_1__4__5), .A1 (L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx16)) ;
    nor02ii L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix17 (.Y (
            L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx16), .A0 (FilterDin_1__4__4), .A1 (
            L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx12)) ;
    xnor2 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix35 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_15), .A0 (
          FilterDin_1__4__6), .A1 (L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx20)) ;
    nor02ii L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix21 (.Y (
            L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx20), .A0 (FilterDin_1__4__5), .A1 (
            L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx16)) ;
    xnor2 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix27 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_16), .A0 (
          FilterDin_1__4__7), .A1 (L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx24)) ;
    nor02ii L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix25 (.Y (
            L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx24), .A0 (FilterDin_1__4__6), .A1 (
            L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx20)) ;
    inv01 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix329 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx328), .A (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx4)) ;
    inv02 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix383 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx384), .A (
          L1_1_L2_4_G1_MINI_ALU_BoothP_0)) ;
    dff L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_0 (.Q (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_0), .QB (\$dummy [463]), 
        .D (L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .CLK (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    nor02_2x L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix567 (.Y (
             L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566), .A0 (RST), .A1 (
             L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644)) ;
    dff L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_1 (.Q (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_1), .QB (\$dummy [464]), 
        .D (L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .CLK (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_2 (.Q (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_2), .QB (\$dummy [465]), 
        .D (L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .CLK (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_3 (.Q (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_3), .QB (\$dummy [466]), 
        .D (L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .CLK (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_4 (.Q (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_4), .QB (\$dummy [467]), 
        .D (L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .CLK (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_5 (.Q (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_5), .QB (\$dummy [468]), 
        .D (L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .CLK (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_6 (.Q (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_6), .QB (\$dummy [469]), 
        .D (L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .CLK (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_7 (.Q (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_7), .QB (\$dummy [470]), 
        .D (L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .CLK (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_8 (.Q (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_8), .QB (\$dummy [471]), 
        .D (L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .CLK (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_9 (.Q (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_9), .QB (\$dummy [472]), 
        .D (L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .CLK (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_10 (.Q (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_10), .QB (\$dummy [473])
        , .D (L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .CLK (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_11 (.Q (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_11), .QB (\$dummy [474])
        , .D (L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .CLK (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_12 (.Q (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_12), .QB (\$dummy [475])
        , .D (L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .CLK (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_13 (.Q (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_13), .QB (\$dummy [476])
        , .D (L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .CLK (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_14 (.Q (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_14), .QB (\$dummy [477])
        , .D (L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .CLK (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_15 (.Q (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_15), .QB (\$dummy [478])
        , .D (L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .CLK (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_16 (.Q (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_16), .QB (\$dummy [479])
        , .D (L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .CLK (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    inv02 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix623 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624), .A (CLK)) ;
    inv02 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix625 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626), .A (CLK)) ;
    inv02 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix627 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628), .A (CLK)) ;
    inv02 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix643 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644), .A (nx7978)) ;
    dff L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_0 (.Q (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_0), .QB (\$dummy [480]), 
        .D (L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .CLK (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    nor02_2x L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix567 (.Y (
             L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566), .A0 (RST), .A1 (
             L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644)) ;
    dff L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_1 (.Q (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_1), .QB (\$dummy [481]), 
        .D (L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .CLK (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_2 (.Q (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_2), .QB (\$dummy [482]), 
        .D (L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .CLK (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_3 (.Q (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_3), .QB (\$dummy [483]), 
        .D (L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .CLK (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_4 (.Q (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_4), .QB (\$dummy [484]), 
        .D (L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .CLK (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_5 (.Q (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_5), .QB (\$dummy [485]), 
        .D (L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .CLK (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_6 (.Q (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_6), .QB (\$dummy [486]), 
        .D (L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .CLK (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_7 (.Q (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_7), .QB (\$dummy [487]), 
        .D (L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .CLK (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_8 (.Q (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_8), .QB (\$dummy [488]), 
        .D (L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .CLK (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_9 (.Q (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_9), .QB (\$dummy [489]), 
        .D (L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .CLK (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_10 (.Q (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_10), .QB (\$dummy [490])
        , .D (L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .CLK (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_11 (.Q (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_11), .QB (\$dummy [491])
        , .D (L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .CLK (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_12 (.Q (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_12), .QB (\$dummy [492])
        , .D (L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .CLK (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_13 (.Q (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_13), .QB (\$dummy [493])
        , .D (L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .CLK (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_14 (.Q (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_14), .QB (\$dummy [494])
        , .D (L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .CLK (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_15 (.Q (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_15), .QB (\$dummy [495])
        , .D (L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .CLK (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_16 (.Q (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_16), .QB (\$dummy [496])
        , .D (L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .CLK (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    inv02 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix623 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624), .A (CLK)) ;
    inv02 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix625 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626), .A (CLK)) ;
    inv02 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix627 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628), .A (CLK)) ;
    inv02 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix643 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644), .A (nx7984)) ;
    dff L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_0 (.Q (
        L1_1_L2_4_G1_MINI_ALU_BoothP_0), .QB (\$dummy [497]), .D (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .CLK (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    nor02_2x L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix567 (.Y (
             L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566), .A0 (RST), .A1 (
             L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    dff L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_1 (.Q (
        L1_1_L2_4_G1_MINI_ALU_BoothP_1), .QB (\$dummy [498]), .D (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .CLK (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_2 (.Q (
        L1_1_L2_4_G1_MINI_ALU_BoothP_2), .QB (\$dummy [499]), .D (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .CLK (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_3 (.Q (
        L1_1_L2_4_G1_MINI_ALU_BoothP_3), .QB (\$dummy [500]), .D (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .CLK (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_4 (.Q (
        L1_1_L2_4_G1_MINI_ALU_BoothP_4), .QB (\$dummy [501]), .D (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .CLK (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_5 (.Q (
        L1_1_L2_4_G1_MINI_ALU_BoothP_5), .QB (\$dummy [502]), .D (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .CLK (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_6 (.Q (
        L1_1_L2_4_G1_MINI_ALU_BoothP_6), .QB (\$dummy [503]), .D (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .CLK (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_7 (.Q (
        L1_1_L2_4_G1_MINI_ALU_BoothP_7), .QB (\$dummy [504]), .D (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .CLK (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_8 (.Q (
        L1_1_L2_4_G1_MINI_ALU_BoothP_8), .QB (\$dummy [505]), .D (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .CLK (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_9 (.Q (
        L1_1_L2_4_G1_MINI_ALU_BoothP_9), .QB (\$dummy [506]), .D (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .CLK (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_10 (.Q (
        L1_1_L2_4_G1_MINI_ALU_BoothP_10), .QB (\$dummy [507]), .D (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .CLK (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_11 (.Q (
        L1_1_L2_4_G1_MINI_ALU_BoothP_11), .QB (\$dummy [508]), .D (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .CLK (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_12 (.Q (
        L1_1_L2_4_G1_MINI_ALU_BoothP_12), .QB (\$dummy [509]), .D (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .CLK (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_13 (.Q (
        L1_1_L2_4_G1_MINI_ALU_BoothP_13), .QB (\$dummy [510]), .D (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .CLK (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_14 (.Q (
        L1_1_L2_4_G1_MINI_ALU_BoothP_14), .QB (\$dummy [511]), .D (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .CLK (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_15 (.Q (
        L1_1_L2_4_G1_MINI_ALU_BoothP_15), .QB (\$dummy [512]), .D (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .CLK (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_16 (.Q (
        L1_1_L2_4_G1_MINI_ALU_BoothP_16), .QB (\$dummy [513]), .D (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .CLK (
        L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    inv02 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix623 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624), .A (CLK)) ;
    inv02 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix625 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626), .A (CLK)) ;
    inv02 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix627 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628), .A (CLK)) ;
    inv02 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix643 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644), .A (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642)) ;
    xor2 L1_2_L2_0_G1_MINI_ALU_ix83 (.Y (L1Results_10__0), .A0 (
         L1SecondOperands_10__0), .A1 (L1FirstOperands_10__0)) ;
    xnor2 L1_2_L2_0_G1_MINI_ALU_ix380 (.Y (L1_2_L2_0_G1_MINI_ALU_nx379), .A0 (
          L1_2_L2_0_G1_MINI_ALU_nx381), .A1 (L1_2_L2_0_G1_MINI_ALU_nx383)) ;
    nand02 L1_2_L2_0_G1_MINI_ALU_ix382 (.Y (L1_2_L2_0_G1_MINI_ALU_nx381), .A0 (
           L1_2_L2_0_G1_MINI_ALU_BoothOperand_0), .A1 (nx8004)) ;
    xnor2 L1_2_L2_0_G1_MINI_ALU_ix384 (.Y (L1_2_L2_0_G1_MINI_ALU_nx383), .A0 (
          L1_2_L2_0_G1_MINI_ALU_BoothOperand_1), .A1 (
          L1_2_L2_0_G1_MINI_ALU_BoothP_1)) ;
    inv01 L1_2_L2_0_G1_MINI_ALU_ix388 (.Y (L1_2_L2_0_G1_MINI_ALU_nx387), .A (
          L1_2_L2_0_G1_MINI_ALU_BoothP_2)) ;
    xnor2 L1_2_L2_0_G1_MINI_ALU_ix390 (.Y (L1_2_L2_0_G1_MINI_ALU_nx389), .A0 (
          L1_2_L2_0_G1_MINI_ALU_nx391), .A1 (L1_2_L2_0_G1_MINI_ALU_nx395)) ;
    aoi32 L1_2_L2_0_G1_MINI_ALU_ix392 (.Y (L1_2_L2_0_G1_MINI_ALU_nx391), .A0 (
          L1_2_L2_0_G1_MINI_ALU_BoothOperand_0), .A1 (nx8004), .A2 (
          L1_2_L2_0_G1_MINI_ALU_nx154), .B0 (L1_2_L2_0_G1_MINI_ALU_BoothP_1), .B1 (
          L1_2_L2_0_G1_MINI_ALU_BoothOperand_1)) ;
    xnor2 L1_2_L2_0_G1_MINI_ALU_ix396 (.Y (L1_2_L2_0_G1_MINI_ALU_nx395), .A0 (
          L1_2_L2_0_G1_MINI_ALU_BoothOperand_2), .A1 (
          L1_2_L2_0_G1_MINI_ALU_BoothP_2)) ;
    inv01 L1_2_L2_0_G1_MINI_ALU_ix400 (.Y (L1_2_L2_0_G1_MINI_ALU_nx399), .A (
          L1_2_L2_0_G1_MINI_ALU_BoothP_3)) ;
    xnor2 L1_2_L2_0_G1_MINI_ALU_ix402 (.Y (L1_2_L2_0_G1_MINI_ALU_nx401), .A0 (
          L1_2_L2_0_G1_MINI_ALU_nx403), .A1 (L1_2_L2_0_G1_MINI_ALU_nx405)) ;
    xnor2 L1_2_L2_0_G1_MINI_ALU_ix406 (.Y (L1_2_L2_0_G1_MINI_ALU_nx405), .A0 (
          L1_2_L2_0_G1_MINI_ALU_BoothOperand_3), .A1 (
          L1_2_L2_0_G1_MINI_ALU_BoothP_3)) ;
    inv01 L1_2_L2_0_G1_MINI_ALU_ix410 (.Y (L1_2_L2_0_G1_MINI_ALU_nx409), .A (
          L1_2_L2_0_G1_MINI_ALU_BoothP_4)) ;
    xnor2 L1_2_L2_0_G1_MINI_ALU_ix412 (.Y (L1_2_L2_0_G1_MINI_ALU_nx411), .A0 (
          L1_2_L2_0_G1_MINI_ALU_nx413), .A1 (L1_2_L2_0_G1_MINI_ALU_nx415)) ;
    xnor2 L1_2_L2_0_G1_MINI_ALU_ix416 (.Y (L1_2_L2_0_G1_MINI_ALU_nx415), .A0 (
          L1_2_L2_0_G1_MINI_ALU_BoothOperand_4), .A1 (
          L1_2_L2_0_G1_MINI_ALU_BoothP_4)) ;
    inv01 L1_2_L2_0_G1_MINI_ALU_ix420 (.Y (L1_2_L2_0_G1_MINI_ALU_nx419), .A (
          L1_2_L2_0_G1_MINI_ALU_BoothP_5)) ;
    xnor2 L1_2_L2_0_G1_MINI_ALU_ix422 (.Y (L1_2_L2_0_G1_MINI_ALU_nx421), .A0 (
          L1_2_L2_0_G1_MINI_ALU_nx423), .A1 (L1_2_L2_0_G1_MINI_ALU_nx425)) ;
    xnor2 L1_2_L2_0_G1_MINI_ALU_ix426 (.Y (L1_2_L2_0_G1_MINI_ALU_nx425), .A0 (
          L1_2_L2_0_G1_MINI_ALU_BoothOperand_5), .A1 (
          L1_2_L2_0_G1_MINI_ALU_BoothP_5)) ;
    inv01 L1_2_L2_0_G1_MINI_ALU_ix430 (.Y (L1_2_L2_0_G1_MINI_ALU_nx429), .A (
          L1_2_L2_0_G1_MINI_ALU_BoothP_6)) ;
    xnor2 L1_2_L2_0_G1_MINI_ALU_ix432 (.Y (L1_2_L2_0_G1_MINI_ALU_nx431), .A0 (
          L1_2_L2_0_G1_MINI_ALU_nx433), .A1 (L1_2_L2_0_G1_MINI_ALU_nx435)) ;
    xnor2 L1_2_L2_0_G1_MINI_ALU_ix436 (.Y (L1_2_L2_0_G1_MINI_ALU_nx435), .A0 (
          L1_2_L2_0_G1_MINI_ALU_BoothOperand_6), .A1 (
          L1_2_L2_0_G1_MINI_ALU_BoothP_6)) ;
    inv01 L1_2_L2_0_G1_MINI_ALU_ix440 (.Y (L1_2_L2_0_G1_MINI_ALU_nx439), .A (
          L1_2_L2_0_G1_MINI_ALU_BoothP_7)) ;
    xnor2 L1_2_L2_0_G1_MINI_ALU_ix442 (.Y (L1_2_L2_0_G1_MINI_ALU_nx441), .A0 (
          L1_2_L2_0_G1_MINI_ALU_nx443), .A1 (L1_2_L2_0_G1_MINI_ALU_nx445)) ;
    xnor2 L1_2_L2_0_G1_MINI_ALU_ix446 (.Y (L1_2_L2_0_G1_MINI_ALU_nx445), .A0 (
          L1_2_L2_0_G1_MINI_ALU_BoothOperand_7), .A1 (
          L1_2_L2_0_G1_MINI_ALU_BoothP_7)) ;
    inv01 L1_2_L2_0_G1_MINI_ALU_ix450 (.Y (L1_2_L2_0_G1_MINI_ALU_nx449), .A (
          L1_2_L2_0_G1_MINI_ALU_BoothP_8)) ;
    xnor2 L1_2_L2_0_G1_MINI_ALU_ix452 (.Y (L1_2_L2_0_G1_MINI_ALU_nx451), .A0 (
          L1_2_L2_0_G1_MINI_ALU_nx453), .A1 (L1_2_L2_0_G1_MINI_ALU_nx455)) ;
    xnor2 L1_2_L2_0_G1_MINI_ALU_ix456 (.Y (L1_2_L2_0_G1_MINI_ALU_nx455), .A0 (
          L1_2_L2_0_G1_MINI_ALU_BoothOperand_8), .A1 (
          L1_2_L2_0_G1_MINI_ALU_BoothP_8)) ;
    xor2 L1_2_L2_0_G1_MINI_ALU_ix317 (.Y (L1_2_L2_0_G1_MINI_ALU_nx316), .A0 (
         L1_2_L2_0_G1_MINI_ALU_nx461), .A1 (L1_2_L2_0_G1_MINI_ALU_nx463)) ;
    xnor2 L1_2_L2_0_G1_MINI_ALU_ix464 (.Y (L1_2_L2_0_G1_MINI_ALU_nx463), .A0 (
          L1_2_L2_0_G1_MINI_ALU_BoothOperand_9), .A1 (
          L1_2_L2_0_G1_MINI_ALU_BoothP_9)) ;
    xor2 L1_2_L2_0_G1_MINI_ALU_ix337 (.Y (L1_2_L2_0_G1_MINI_ALU_nx336), .A0 (
         L1_2_L2_0_G1_MINI_ALU_nx467), .A1 (L1_2_L2_0_G1_MINI_ALU_nx471)) ;
    inv01 L1_2_L2_0_G1_MINI_ALU_ix470 (.Y (L1_2_L2_0_G1_MINI_ALU_nx469), .A (
          L1_2_L2_0_G1_MINI_ALU_BoothP_9)) ;
    xnor2 L1_2_L2_0_G1_MINI_ALU_ix472 (.Y (L1_2_L2_0_G1_MINI_ALU_nx471), .A0 (
          L1_2_L2_0_G1_MINI_ALU_BoothOperand_10), .A1 (
          L1_2_L2_0_G1_MINI_ALU_BoothP_10)) ;
    xor2 L1_2_L2_0_G1_MINI_ALU_ix357 (.Y (L1_2_L2_0_G1_MINI_ALU_nx356), .A0 (
         L1_2_L2_0_G1_MINI_ALU_nx475), .A1 (L1_2_L2_0_G1_MINI_ALU_nx479)) ;
    inv01 L1_2_L2_0_G1_MINI_ALU_ix478 (.Y (L1_2_L2_0_G1_MINI_ALU_nx477), .A (
          L1_2_L2_0_G1_MINI_ALU_BoothP_10)) ;
    xnor2 L1_2_L2_0_G1_MINI_ALU_ix480 (.Y (L1_2_L2_0_G1_MINI_ALU_nx479), .A0 (
          L1_2_L2_0_G1_MINI_ALU_BoothOperand_11), .A1 (
          L1_2_L2_0_G1_MINI_ALU_BoothP_11)) ;
    xor2 L1_2_L2_0_G1_MINI_ALU_ix377 (.Y (L1_2_L2_0_G1_MINI_ALU_nx376), .A0 (
         L1_2_L2_0_G1_MINI_ALU_nx483), .A1 (L1_2_L2_0_G1_MINI_ALU_nx487)) ;
    inv01 L1_2_L2_0_G1_MINI_ALU_ix486 (.Y (L1_2_L2_0_G1_MINI_ALU_nx485), .A (
          L1_2_L2_0_G1_MINI_ALU_BoothP_11)) ;
    xnor2 L1_2_L2_0_G1_MINI_ALU_ix488 (.Y (L1_2_L2_0_G1_MINI_ALU_nx487), .A0 (
          L1_2_L2_0_G1_MINI_ALU_BoothOperand_12), .A1 (
          L1_2_L2_0_G1_MINI_ALU_BoothP_12)) ;
    xor2 L1_2_L2_0_G1_MINI_ALU_ix397 (.Y (L1_2_L2_0_G1_MINI_ALU_nx396), .A0 (
         L1_2_L2_0_G1_MINI_ALU_nx491), .A1 (L1_2_L2_0_G1_MINI_ALU_nx495)) ;
    inv01 L1_2_L2_0_G1_MINI_ALU_ix494 (.Y (L1_2_L2_0_G1_MINI_ALU_nx493), .A (
          L1_2_L2_0_G1_MINI_ALU_BoothP_12)) ;
    xnor2 L1_2_L2_0_G1_MINI_ALU_ix496 (.Y (L1_2_L2_0_G1_MINI_ALU_nx495), .A0 (
          L1_2_L2_0_G1_MINI_ALU_BoothOperand_13), .A1 (
          L1_2_L2_0_G1_MINI_ALU_BoothP_13)) ;
    xor2 L1_2_L2_0_G1_MINI_ALU_ix417 (.Y (L1_2_L2_0_G1_MINI_ALU_nx416), .A0 (
         L1_2_L2_0_G1_MINI_ALU_nx499), .A1 (L1_2_L2_0_G1_MINI_ALU_nx503)) ;
    inv01 L1_2_L2_0_G1_MINI_ALU_ix502 (.Y (L1_2_L2_0_G1_MINI_ALU_nx501), .A (
          L1_2_L2_0_G1_MINI_ALU_BoothP_13)) ;
    xnor2 L1_2_L2_0_G1_MINI_ALU_ix504 (.Y (L1_2_L2_0_G1_MINI_ALU_nx503), .A0 (
          L1_2_L2_0_G1_MINI_ALU_BoothOperand_14), .A1 (
          L1_2_L2_0_G1_MINI_ALU_BoothP_14)) ;
    xor2 L1_2_L2_0_G1_MINI_ALU_ix437 (.Y (L1_2_L2_0_G1_MINI_ALU_nx436), .A0 (
         L1_2_L2_0_G1_MINI_ALU_nx507), .A1 (L1_2_L2_0_G1_MINI_ALU_nx511)) ;
    inv01 L1_2_L2_0_G1_MINI_ALU_ix510 (.Y (L1_2_L2_0_G1_MINI_ALU_nx509), .A (
          L1_2_L2_0_G1_MINI_ALU_BoothP_14)) ;
    xnor2 L1_2_L2_0_G1_MINI_ALU_ix512 (.Y (L1_2_L2_0_G1_MINI_ALU_nx511), .A0 (
          L1_2_L2_0_G1_MINI_ALU_BoothOperand_15), .A1 (
          L1_2_L2_0_G1_MINI_ALU_BoothP_15)) ;
    xnor2 L1_2_L2_0_G1_MINI_ALU_ix457 (.Y (L1_2_L2_0_G1_MINI_ALU_nx456), .A0 (
          L1_2_L2_0_G1_MINI_ALU_nx515), .A1 (L1_2_L2_0_G1_MINI_ALU_nx454)) ;
    inv01 L1_2_L2_0_G1_MINI_ALU_ix518 (.Y (L1_2_L2_0_G1_MINI_ALU_nx517), .A (
          L1_2_L2_0_G1_MINI_ALU_BoothP_15)) ;
    xor2 L1_2_L2_0_G1_MINI_ALU_ix455 (.Y (L1_2_L2_0_G1_MINI_ALU_nx454), .A0 (
         L1_2_L2_0_G1_MINI_ALU_BoothOperand_16), .A1 (
         L1_2_L2_0_G1_MINI_ALU_BoothP_16)) ;
    mux21_ni L1_2_L2_0_G1_MINI_ALU_ix91 (.Y (L1SecondOperands_10__0), .A0 (
             L1_2_L2_0_G1_MINI_ALU_BoothP_1), .A1 (WindowDin_2__0__0), .S0 (
             Instr)) ;
    mux21_ni L1_2_L2_0_G1_MINI_ALU_ix99 (.Y (L1SecondOperands_10__1), .A0 (
             L1_2_L2_0_G1_MINI_ALU_BoothP_2), .A1 (WindowDin_2__0__1), .S0 (
             Instr)) ;
    mux21_ni L1_2_L2_0_G1_MINI_ALU_ix107 (.Y (L1SecondOperands_10__2), .A0 (
             L1_2_L2_0_G1_MINI_ALU_BoothP_3), .A1 (WindowDin_2__0__2), .S0 (
             Instr)) ;
    mux21_ni L1_2_L2_0_G1_MINI_ALU_ix115 (.Y (L1SecondOperands_10__3), .A0 (
             L1_2_L2_0_G1_MINI_ALU_BoothP_4), .A1 (WindowDin_2__0__3), .S0 (
             Instr)) ;
    mux21_ni L1_2_L2_0_G1_MINI_ALU_ix123 (.Y (L1SecondOperands_10__4), .A0 (
             L1_2_L2_0_G1_MINI_ALU_BoothP_5), .A1 (WindowDin_2__0__4), .S0 (
             Instr)) ;
    mux21_ni L1_2_L2_0_G1_MINI_ALU_ix131 (.Y (L1SecondOperands_10__5), .A0 (
             L1_2_L2_0_G1_MINI_ALU_BoothP_6), .A1 (WindowDin_2__0__5), .S0 (
             Instr)) ;
    mux21_ni L1_2_L2_0_G1_MINI_ALU_ix139 (.Y (L1SecondOperands_10__6), .A0 (
             L1_2_L2_0_G1_MINI_ALU_BoothP_7), .A1 (WindowDin_2__0__6), .S0 (
             Instr)) ;
    mux21_ni L1_2_L2_0_G1_MINI_ALU_ix147 (.Y (L1SecondOperands_10__7), .A0 (
             L1_2_L2_0_G1_MINI_ALU_BoothP_8), .A1 (WindowDin_2__0__7), .S0 (
             Instr)) ;
    xor2 L1_2_L2_0_G1_MINI_ALU_ix77 (.Y (L1Results_10__1), .A0 (
         L1_2_L2_0_G1_MINI_ALU_nx529), .A1 (L1_2_L2_0_G1_MINI_ALU_nx531)) ;
    nand02 L1_2_L2_0_G1_MINI_ALU_ix530 (.Y (L1_2_L2_0_G1_MINI_ALU_nx529), .A0 (
           L1SecondOperands_10__0), .A1 (L1FirstOperands_10__0)) ;
    xnor2 L1_2_L2_0_G1_MINI_ALU_ix532 (.Y (L1_2_L2_0_G1_MINI_ALU_nx531), .A0 (
          L1SecondOperands_10__1), .A1 (L1FirstOperands_10__1)) ;
    xor2 L1_2_L2_0_G1_MINI_ALU_ix75 (.Y (L1Results_10__2), .A0 (
         L1_2_L2_0_G1_MINI_ALU_nx534), .A1 (L1_2_L2_0_G1_MINI_ALU_nx537)) ;
    aoi32 L1_2_L2_0_G1_MINI_ALU_ix535 (.Y (L1_2_L2_0_G1_MINI_ALU_nx534), .A0 (
          L1SecondOperands_10__0), .A1 (L1FirstOperands_10__0), .A2 (
          L1_2_L2_0_G1_MINI_ALU_nx30), .B0 (L1FirstOperands_10__1), .B1 (
          L1SecondOperands_10__1)) ;
    xnor2 L1_2_L2_0_G1_MINI_ALU_ix538 (.Y (L1_2_L2_0_G1_MINI_ALU_nx537), .A0 (
          L1SecondOperands_10__2), .A1 (L1FirstOperands_10__2)) ;
    xor2 L1_2_L2_0_G1_MINI_ALU_ix73 (.Y (L1Results_10__3), .A0 (
         L1_2_L2_0_G1_MINI_ALU_nx540), .A1 (L1_2_L2_0_G1_MINI_ALU_nx544)) ;
    aoi22 L1_2_L2_0_G1_MINI_ALU_ix541 (.Y (L1_2_L2_0_G1_MINI_ALU_nx540), .A0 (
          L1FirstOperands_10__2), .A1 (L1SecondOperands_10__2), .B0 (
          L1_2_L2_0_G1_MINI_ALU_nx40), .B1 (L1_2_L2_0_G1_MINI_ALU_nx24)) ;
    xnor2 L1_2_L2_0_G1_MINI_ALU_ix545 (.Y (L1_2_L2_0_G1_MINI_ALU_nx544), .A0 (
          L1SecondOperands_10__3), .A1 (L1FirstOperands_10__3)) ;
    xor2 L1_2_L2_0_G1_MINI_ALU_ix71 (.Y (L1Results_10__4), .A0 (
         L1_2_L2_0_G1_MINI_ALU_nx547), .A1 (L1_2_L2_0_G1_MINI_ALU_nx551)) ;
    aoi22 L1_2_L2_0_G1_MINI_ALU_ix548 (.Y (L1_2_L2_0_G1_MINI_ALU_nx547), .A0 (
          L1FirstOperands_10__3), .A1 (L1SecondOperands_10__3), .B0 (
          L1_2_L2_0_G1_MINI_ALU_nx44), .B1 (L1_2_L2_0_G1_MINI_ALU_nx18)) ;
    xnor2 L1_2_L2_0_G1_MINI_ALU_ix552 (.Y (L1_2_L2_0_G1_MINI_ALU_nx551), .A0 (
          L1SecondOperands_10__4), .A1 (L1FirstOperands_10__4)) ;
    xor2 L1_2_L2_0_G1_MINI_ALU_ix69 (.Y (L1Results_10__5), .A0 (
         L1_2_L2_0_G1_MINI_ALU_nx554), .A1 (L1_2_L2_0_G1_MINI_ALU_nx558)) ;
    aoi22 L1_2_L2_0_G1_MINI_ALU_ix555 (.Y (L1_2_L2_0_G1_MINI_ALU_nx554), .A0 (
          L1FirstOperands_10__4), .A1 (L1SecondOperands_10__4), .B0 (
          L1_2_L2_0_G1_MINI_ALU_nx48), .B1 (L1_2_L2_0_G1_MINI_ALU_nx12)) ;
    xnor2 L1_2_L2_0_G1_MINI_ALU_ix559 (.Y (L1_2_L2_0_G1_MINI_ALU_nx558), .A0 (
          L1SecondOperands_10__5), .A1 (L1FirstOperands_10__5)) ;
    xor2 L1_2_L2_0_G1_MINI_ALU_ix67 (.Y (L1Results_10__6), .A0 (
         L1_2_L2_0_G1_MINI_ALU_nx561), .A1 (L1_2_L2_0_G1_MINI_ALU_nx565)) ;
    aoi22 L1_2_L2_0_G1_MINI_ALU_ix562 (.Y (L1_2_L2_0_G1_MINI_ALU_nx561), .A0 (
          L1FirstOperands_10__5), .A1 (L1SecondOperands_10__5), .B0 (
          L1_2_L2_0_G1_MINI_ALU_nx52), .B1 (L1_2_L2_0_G1_MINI_ALU_nx6)) ;
    xnor2 L1_2_L2_0_G1_MINI_ALU_ix566 (.Y (L1_2_L2_0_G1_MINI_ALU_nx565), .A0 (
          L1SecondOperands_10__6), .A1 (L1FirstOperands_10__6)) ;
    xnor2 L1_2_L2_0_G1_MINI_ALU_ix65 (.Y (L1Results_10__7), .A0 (
          L1_2_L2_0_G1_MINI_ALU_nx568), .A1 (L1_2_L2_0_G1_MINI_ALU_nx62)) ;
    aoi22 L1_2_L2_0_G1_MINI_ALU_ix569 (.Y (L1_2_L2_0_G1_MINI_ALU_nx568), .A0 (
          L1FirstOperands_10__6), .A1 (L1SecondOperands_10__6), .B0 (
          L1_2_L2_0_G1_MINI_ALU_nx56), .B1 (L1_2_L2_0_G1_MINI_ALU_nx0)) ;
    xor2 L1_2_L2_0_G1_MINI_ALU_ix63 (.Y (L1_2_L2_0_G1_MINI_ALU_nx62), .A0 (
         L1SecondOperands_10__7), .A1 (L1FirstOperands_10__7)) ;
    inv01 L1_2_L2_0_G1_MINI_ALU_ix155 (.Y (L1_2_L2_0_G1_MINI_ALU_nx154), .A (
          L1_2_L2_0_G1_MINI_ALU_nx383)) ;
    inv01 L1_2_L2_0_G1_MINI_ALU_ix57 (.Y (L1_2_L2_0_G1_MINI_ALU_nx56), .A (
          L1_2_L2_0_G1_MINI_ALU_nx561)) ;
    inv01 L1_2_L2_0_G1_MINI_ALU_ix53 (.Y (L1_2_L2_0_G1_MINI_ALU_nx52), .A (
          L1_2_L2_0_G1_MINI_ALU_nx554)) ;
    inv01 L1_2_L2_0_G1_MINI_ALU_ix49 (.Y (L1_2_L2_0_G1_MINI_ALU_nx48), .A (
          L1_2_L2_0_G1_MINI_ALU_nx547)) ;
    inv01 L1_2_L2_0_G1_MINI_ALU_ix45 (.Y (L1_2_L2_0_G1_MINI_ALU_nx44), .A (
          L1_2_L2_0_G1_MINI_ALU_nx540)) ;
    inv01 L1_2_L2_0_G1_MINI_ALU_ix41 (.Y (L1_2_L2_0_G1_MINI_ALU_nx40), .A (
          L1_2_L2_0_G1_MINI_ALU_nx534)) ;
    inv01 L1_2_L2_0_G1_MINI_ALU_ix31 (.Y (L1_2_L2_0_G1_MINI_ALU_nx30), .A (
          L1_2_L2_0_G1_MINI_ALU_nx531)) ;
    inv01 L1_2_L2_0_G1_MINI_ALU_ix25 (.Y (L1_2_L2_0_G1_MINI_ALU_nx24), .A (
          L1_2_L2_0_G1_MINI_ALU_nx537)) ;
    inv01 L1_2_L2_0_G1_MINI_ALU_ix19 (.Y (L1_2_L2_0_G1_MINI_ALU_nx18), .A (
          L1_2_L2_0_G1_MINI_ALU_nx544)) ;
    inv01 L1_2_L2_0_G1_MINI_ALU_ix13 (.Y (L1_2_L2_0_G1_MINI_ALU_nx12), .A (
          L1_2_L2_0_G1_MINI_ALU_nx551)) ;
    inv01 L1_2_L2_0_G1_MINI_ALU_ix7 (.Y (L1_2_L2_0_G1_MINI_ALU_nx6), .A (
          L1_2_L2_0_G1_MINI_ALU_nx558)) ;
    inv01 L1_2_L2_0_G1_MINI_ALU_ix1 (.Y (L1_2_L2_0_G1_MINI_ALU_nx0), .A (
          L1_2_L2_0_G1_MINI_ALU_nx565)) ;
    fake_gnd L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix216 (.Y (
             L1_2_L2_0_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    nor02ii L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix81 (.Y (
            L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx80), .A0 (Instr), .A1 (Start)) ;
    aoi21 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix77 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_10), .A0 (
          FilterDin_2__0__1), .A1 (FilterDin_2__0__0), .B0 (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx4)) ;
    nor02_2x L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix5 (.Y (
             L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx4), .A0 (FilterDin_2__0__0), .A1 (
             FilterDin_2__0__1)) ;
    aoi21 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix67 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_11), .A0 (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx328), .A1 (FilterDin_2__0__2), .B0 (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx8)) ;
    nor03_2x L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix9 (.Y (
             L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx8), .A0 (FilterDin_2__0__2), .A1 (
             FilterDin_2__0__0), .A2 (FilterDin_2__0__1)) ;
    xnor2 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix59 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_12), .A0 (
          FilterDin_2__0__3), .A1 (L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx8)) ;
    xnor2 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix51 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_13), .A0 (
          FilterDin_2__0__4), .A1 (L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx12)) ;
    nor04 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix13 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx12), .A0 (FilterDin_2__0__3), .A1 (
          FilterDin_2__0__2), .A2 (FilterDin_2__0__0), .A3 (FilterDin_2__0__1)
          ) ;
    xnor2 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix43 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_14), .A0 (
          FilterDin_2__0__5), .A1 (L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx16)) ;
    nor02ii L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix17 (.Y (
            L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx16), .A0 (FilterDin_2__0__4), .A1 (
            L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx12)) ;
    xnor2 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix35 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_15), .A0 (
          FilterDin_2__0__6), .A1 (L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx20)) ;
    nor02ii L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix21 (.Y (
            L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx20), .A0 (FilterDin_2__0__5), .A1 (
            L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx16)) ;
    xnor2 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix27 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_16), .A0 (
          FilterDin_2__0__7), .A1 (L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx24)) ;
    nor02ii L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix25 (.Y (
            L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx24), .A0 (FilterDin_2__0__6), .A1 (
            L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx20)) ;
    inv01 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix329 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx328), .A (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx4)) ;
    inv02 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix383 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx384), .A (
          L1_2_L2_0_G1_MINI_ALU_BoothP_0)) ;
    dff L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_0 (.Q (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_0), .QB (\$dummy [514]), 
        .D (L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .CLK (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    nor02_2x L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix567 (.Y (
             L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566), .A0 (RST), .A1 (
             L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644)) ;
    dff L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_1 (.Q (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_1), .QB (\$dummy [515]), 
        .D (L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .CLK (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_2 (.Q (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_2), .QB (\$dummy [516]), 
        .D (L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .CLK (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_3 (.Q (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_3), .QB (\$dummy [517]), 
        .D (L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .CLK (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_4 (.Q (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_4), .QB (\$dummy [518]), 
        .D (L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .CLK (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_5 (.Q (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_5), .QB (\$dummy [519]), 
        .D (L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .CLK (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_6 (.Q (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_6), .QB (\$dummy [520]), 
        .D (L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .CLK (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_7 (.Q (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_7), .QB (\$dummy [521]), 
        .D (L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .CLK (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_8 (.Q (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_8), .QB (\$dummy [522]), 
        .D (L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .CLK (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_9 (.Q (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_9), .QB (\$dummy [523]), 
        .D (L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .CLK (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_10 (.Q (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_10), .QB (\$dummy [524])
        , .D (L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .CLK (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_11 (.Q (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_11), .QB (\$dummy [525])
        , .D (L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .CLK (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_12 (.Q (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_12), .QB (\$dummy [526])
        , .D (L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .CLK (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_13 (.Q (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_13), .QB (\$dummy [527])
        , .D (L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .CLK (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_14 (.Q (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_14), .QB (\$dummy [528])
        , .D (L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .CLK (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_15 (.Q (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_15), .QB (\$dummy [529])
        , .D (L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .CLK (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_16 (.Q (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_16), .QB (\$dummy [530])
        , .D (L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .CLK (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    inv02 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix623 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624), .A (CLK)) ;
    inv02 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix625 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626), .A (CLK)) ;
    inv02 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix627 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628), .A (CLK)) ;
    inv02 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix643 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644), .A (nx8018)) ;
    dff L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_0 (.Q (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_0), .QB (\$dummy [531]), 
        .D (L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .CLK (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    nor02_2x L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix567 (.Y (
             L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566), .A0 (RST), .A1 (
             L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644)) ;
    dff L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_1 (.Q (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_1), .QB (\$dummy [532]), 
        .D (L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .CLK (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_2 (.Q (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_2), .QB (\$dummy [533]), 
        .D (L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .CLK (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_3 (.Q (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_3), .QB (\$dummy [534]), 
        .D (L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .CLK (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_4 (.Q (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_4), .QB (\$dummy [535]), 
        .D (L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .CLK (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_5 (.Q (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_5), .QB (\$dummy [536]), 
        .D (L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .CLK (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_6 (.Q (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_6), .QB (\$dummy [537]), 
        .D (L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .CLK (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_7 (.Q (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_7), .QB (\$dummy [538]), 
        .D (L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .CLK (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_8 (.Q (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_8), .QB (\$dummy [539]), 
        .D (L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .CLK (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_9 (.Q (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_9), .QB (\$dummy [540]), 
        .D (L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .CLK (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_10 (.Q (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_10), .QB (\$dummy [541])
        , .D (L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .CLK (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_11 (.Q (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_11), .QB (\$dummy [542])
        , .D (L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .CLK (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_12 (.Q (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_12), .QB (\$dummy [543])
        , .D (L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .CLK (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_13 (.Q (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_13), .QB (\$dummy [544])
        , .D (L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .CLK (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_14 (.Q (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_14), .QB (\$dummy [545])
        , .D (L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .CLK (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_15 (.Q (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_15), .QB (\$dummy [546])
        , .D (L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .CLK (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_16 (.Q (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_16), .QB (\$dummy [547])
        , .D (L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .CLK (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    inv02 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix623 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624), .A (CLK)) ;
    inv02 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix625 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626), .A (CLK)) ;
    inv02 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix627 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628), .A (CLK)) ;
    inv02 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix643 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644), .A (nx8024)) ;
    dff L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_0 (.Q (
        L1_2_L2_0_G1_MINI_ALU_BoothP_0), .QB (\$dummy [548]), .D (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .CLK (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    nor02_2x L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix567 (.Y (
             L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566), .A0 (RST), .A1 (
             L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    dff L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_1 (.Q (
        L1_2_L2_0_G1_MINI_ALU_BoothP_1), .QB (\$dummy [549]), .D (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .CLK (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_2 (.Q (
        L1_2_L2_0_G1_MINI_ALU_BoothP_2), .QB (\$dummy [550]), .D (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .CLK (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_3 (.Q (
        L1_2_L2_0_G1_MINI_ALU_BoothP_3), .QB (\$dummy [551]), .D (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .CLK (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_4 (.Q (
        L1_2_L2_0_G1_MINI_ALU_BoothP_4), .QB (\$dummy [552]), .D (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .CLK (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_5 (.Q (
        L1_2_L2_0_G1_MINI_ALU_BoothP_5), .QB (\$dummy [553]), .D (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .CLK (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_6 (.Q (
        L1_2_L2_0_G1_MINI_ALU_BoothP_6), .QB (\$dummy [554]), .D (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .CLK (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_7 (.Q (
        L1_2_L2_0_G1_MINI_ALU_BoothP_7), .QB (\$dummy [555]), .D (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .CLK (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_8 (.Q (
        L1_2_L2_0_G1_MINI_ALU_BoothP_8), .QB (\$dummy [556]), .D (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .CLK (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_9 (.Q (
        L1_2_L2_0_G1_MINI_ALU_BoothP_9), .QB (\$dummy [557]), .D (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .CLK (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_10 (.Q (
        L1_2_L2_0_G1_MINI_ALU_BoothP_10), .QB (\$dummy [558]), .D (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .CLK (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_11 (.Q (
        L1_2_L2_0_G1_MINI_ALU_BoothP_11), .QB (\$dummy [559]), .D (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .CLK (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_12 (.Q (
        L1_2_L2_0_G1_MINI_ALU_BoothP_12), .QB (\$dummy [560]), .D (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .CLK (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_13 (.Q (
        L1_2_L2_0_G1_MINI_ALU_BoothP_13), .QB (\$dummy [561]), .D (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .CLK (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_14 (.Q (
        L1_2_L2_0_G1_MINI_ALU_BoothP_14), .QB (\$dummy [562]), .D (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .CLK (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_15 (.Q (
        L1_2_L2_0_G1_MINI_ALU_BoothP_15), .QB (\$dummy [563]), .D (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .CLK (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_16 (.Q (
        L1_2_L2_0_G1_MINI_ALU_BoothP_16), .QB (\$dummy [564]), .D (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .CLK (
        L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    inv02 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix623 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624), .A (CLK)) ;
    inv02 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix625 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626), .A (CLK)) ;
    inv02 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix627 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628), .A (CLK)) ;
    inv02 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix643 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644), .A (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642)) ;
    xor2 L1_2_L2_1_G1_MINI_ALU_ix83 (.Y (L1Results_11__0), .A0 (
         L1SecondOperands_11__0), .A1 (L1FirstOperands_11__0)) ;
    xnor2 L1_2_L2_1_G1_MINI_ALU_ix380 (.Y (L1_2_L2_1_G1_MINI_ALU_nx379), .A0 (
          L1_2_L2_1_G1_MINI_ALU_nx381), .A1 (L1_2_L2_1_G1_MINI_ALU_nx383)) ;
    nand02 L1_2_L2_1_G1_MINI_ALU_ix382 (.Y (L1_2_L2_1_G1_MINI_ALU_nx381), .A0 (
           L1_2_L2_1_G1_MINI_ALU_BoothOperand_0), .A1 (nx8044)) ;
    xnor2 L1_2_L2_1_G1_MINI_ALU_ix384 (.Y (L1_2_L2_1_G1_MINI_ALU_nx383), .A0 (
          L1_2_L2_1_G1_MINI_ALU_BoothOperand_1), .A1 (
          L1_2_L2_1_G1_MINI_ALU_BoothP_1)) ;
    inv01 L1_2_L2_1_G1_MINI_ALU_ix388 (.Y (L1_2_L2_1_G1_MINI_ALU_nx387), .A (
          L1_2_L2_1_G1_MINI_ALU_BoothP_2)) ;
    xnor2 L1_2_L2_1_G1_MINI_ALU_ix390 (.Y (L1_2_L2_1_G1_MINI_ALU_nx389), .A0 (
          L1_2_L2_1_G1_MINI_ALU_nx391), .A1 (L1_2_L2_1_G1_MINI_ALU_nx395)) ;
    aoi32 L1_2_L2_1_G1_MINI_ALU_ix392 (.Y (L1_2_L2_1_G1_MINI_ALU_nx391), .A0 (
          L1_2_L2_1_G1_MINI_ALU_BoothOperand_0), .A1 (nx8044), .A2 (
          L1_2_L2_1_G1_MINI_ALU_nx154), .B0 (L1_2_L2_1_G1_MINI_ALU_BoothP_1), .B1 (
          L1_2_L2_1_G1_MINI_ALU_BoothOperand_1)) ;
    xnor2 L1_2_L2_1_G1_MINI_ALU_ix396 (.Y (L1_2_L2_1_G1_MINI_ALU_nx395), .A0 (
          L1_2_L2_1_G1_MINI_ALU_BoothOperand_2), .A1 (
          L1_2_L2_1_G1_MINI_ALU_BoothP_2)) ;
    inv01 L1_2_L2_1_G1_MINI_ALU_ix400 (.Y (L1_2_L2_1_G1_MINI_ALU_nx399), .A (
          L1_2_L2_1_G1_MINI_ALU_BoothP_3)) ;
    xnor2 L1_2_L2_1_G1_MINI_ALU_ix402 (.Y (L1_2_L2_1_G1_MINI_ALU_nx401), .A0 (
          L1_2_L2_1_G1_MINI_ALU_nx403), .A1 (L1_2_L2_1_G1_MINI_ALU_nx405)) ;
    xnor2 L1_2_L2_1_G1_MINI_ALU_ix406 (.Y (L1_2_L2_1_G1_MINI_ALU_nx405), .A0 (
          L1_2_L2_1_G1_MINI_ALU_BoothOperand_3), .A1 (
          L1_2_L2_1_G1_MINI_ALU_BoothP_3)) ;
    inv01 L1_2_L2_1_G1_MINI_ALU_ix410 (.Y (L1_2_L2_1_G1_MINI_ALU_nx409), .A (
          L1_2_L2_1_G1_MINI_ALU_BoothP_4)) ;
    xnor2 L1_2_L2_1_G1_MINI_ALU_ix412 (.Y (L1_2_L2_1_G1_MINI_ALU_nx411), .A0 (
          L1_2_L2_1_G1_MINI_ALU_nx413), .A1 (L1_2_L2_1_G1_MINI_ALU_nx415)) ;
    xnor2 L1_2_L2_1_G1_MINI_ALU_ix416 (.Y (L1_2_L2_1_G1_MINI_ALU_nx415), .A0 (
          L1_2_L2_1_G1_MINI_ALU_BoothOperand_4), .A1 (
          L1_2_L2_1_G1_MINI_ALU_BoothP_4)) ;
    inv01 L1_2_L2_1_G1_MINI_ALU_ix420 (.Y (L1_2_L2_1_G1_MINI_ALU_nx419), .A (
          L1_2_L2_1_G1_MINI_ALU_BoothP_5)) ;
    xnor2 L1_2_L2_1_G1_MINI_ALU_ix422 (.Y (L1_2_L2_1_G1_MINI_ALU_nx421), .A0 (
          L1_2_L2_1_G1_MINI_ALU_nx423), .A1 (L1_2_L2_1_G1_MINI_ALU_nx425)) ;
    xnor2 L1_2_L2_1_G1_MINI_ALU_ix426 (.Y (L1_2_L2_1_G1_MINI_ALU_nx425), .A0 (
          L1_2_L2_1_G1_MINI_ALU_BoothOperand_5), .A1 (
          L1_2_L2_1_G1_MINI_ALU_BoothP_5)) ;
    inv01 L1_2_L2_1_G1_MINI_ALU_ix430 (.Y (L1_2_L2_1_G1_MINI_ALU_nx429), .A (
          L1_2_L2_1_G1_MINI_ALU_BoothP_6)) ;
    xnor2 L1_2_L2_1_G1_MINI_ALU_ix432 (.Y (L1_2_L2_1_G1_MINI_ALU_nx431), .A0 (
          L1_2_L2_1_G1_MINI_ALU_nx433), .A1 (L1_2_L2_1_G1_MINI_ALU_nx435)) ;
    xnor2 L1_2_L2_1_G1_MINI_ALU_ix436 (.Y (L1_2_L2_1_G1_MINI_ALU_nx435), .A0 (
          L1_2_L2_1_G1_MINI_ALU_BoothOperand_6), .A1 (
          L1_2_L2_1_G1_MINI_ALU_BoothP_6)) ;
    inv01 L1_2_L2_1_G1_MINI_ALU_ix440 (.Y (L1_2_L2_1_G1_MINI_ALU_nx439), .A (
          L1_2_L2_1_G1_MINI_ALU_BoothP_7)) ;
    xnor2 L1_2_L2_1_G1_MINI_ALU_ix442 (.Y (L1_2_L2_1_G1_MINI_ALU_nx441), .A0 (
          L1_2_L2_1_G1_MINI_ALU_nx443), .A1 (L1_2_L2_1_G1_MINI_ALU_nx445)) ;
    xnor2 L1_2_L2_1_G1_MINI_ALU_ix446 (.Y (L1_2_L2_1_G1_MINI_ALU_nx445), .A0 (
          L1_2_L2_1_G1_MINI_ALU_BoothOperand_7), .A1 (
          L1_2_L2_1_G1_MINI_ALU_BoothP_7)) ;
    inv01 L1_2_L2_1_G1_MINI_ALU_ix450 (.Y (L1_2_L2_1_G1_MINI_ALU_nx449), .A (
          L1_2_L2_1_G1_MINI_ALU_BoothP_8)) ;
    xnor2 L1_2_L2_1_G1_MINI_ALU_ix452 (.Y (L1_2_L2_1_G1_MINI_ALU_nx451), .A0 (
          L1_2_L2_1_G1_MINI_ALU_nx453), .A1 (L1_2_L2_1_G1_MINI_ALU_nx455)) ;
    xnor2 L1_2_L2_1_G1_MINI_ALU_ix456 (.Y (L1_2_L2_1_G1_MINI_ALU_nx455), .A0 (
          L1_2_L2_1_G1_MINI_ALU_BoothOperand_8), .A1 (
          L1_2_L2_1_G1_MINI_ALU_BoothP_8)) ;
    xor2 L1_2_L2_1_G1_MINI_ALU_ix317 (.Y (L1_2_L2_1_G1_MINI_ALU_nx316), .A0 (
         L1_2_L2_1_G1_MINI_ALU_nx461), .A1 (L1_2_L2_1_G1_MINI_ALU_nx463)) ;
    xnor2 L1_2_L2_1_G1_MINI_ALU_ix464 (.Y (L1_2_L2_1_G1_MINI_ALU_nx463), .A0 (
          L1_2_L2_1_G1_MINI_ALU_BoothOperand_9), .A1 (
          L1_2_L2_1_G1_MINI_ALU_BoothP_9)) ;
    xor2 L1_2_L2_1_G1_MINI_ALU_ix337 (.Y (L1_2_L2_1_G1_MINI_ALU_nx336), .A0 (
         L1_2_L2_1_G1_MINI_ALU_nx467), .A1 (L1_2_L2_1_G1_MINI_ALU_nx471)) ;
    inv01 L1_2_L2_1_G1_MINI_ALU_ix470 (.Y (L1_2_L2_1_G1_MINI_ALU_nx469), .A (
          L1_2_L2_1_G1_MINI_ALU_BoothP_9)) ;
    xnor2 L1_2_L2_1_G1_MINI_ALU_ix472 (.Y (L1_2_L2_1_G1_MINI_ALU_nx471), .A0 (
          L1_2_L2_1_G1_MINI_ALU_BoothOperand_10), .A1 (
          L1_2_L2_1_G1_MINI_ALU_BoothP_10)) ;
    xor2 L1_2_L2_1_G1_MINI_ALU_ix357 (.Y (L1_2_L2_1_G1_MINI_ALU_nx356), .A0 (
         L1_2_L2_1_G1_MINI_ALU_nx475), .A1 (L1_2_L2_1_G1_MINI_ALU_nx479)) ;
    inv01 L1_2_L2_1_G1_MINI_ALU_ix478 (.Y (L1_2_L2_1_G1_MINI_ALU_nx477), .A (
          L1_2_L2_1_G1_MINI_ALU_BoothP_10)) ;
    xnor2 L1_2_L2_1_G1_MINI_ALU_ix480 (.Y (L1_2_L2_1_G1_MINI_ALU_nx479), .A0 (
          L1_2_L2_1_G1_MINI_ALU_BoothOperand_11), .A1 (
          L1_2_L2_1_G1_MINI_ALU_BoothP_11)) ;
    xor2 L1_2_L2_1_G1_MINI_ALU_ix377 (.Y (L1_2_L2_1_G1_MINI_ALU_nx376), .A0 (
         L1_2_L2_1_G1_MINI_ALU_nx483), .A1 (L1_2_L2_1_G1_MINI_ALU_nx487)) ;
    inv01 L1_2_L2_1_G1_MINI_ALU_ix486 (.Y (L1_2_L2_1_G1_MINI_ALU_nx485), .A (
          L1_2_L2_1_G1_MINI_ALU_BoothP_11)) ;
    xnor2 L1_2_L2_1_G1_MINI_ALU_ix488 (.Y (L1_2_L2_1_G1_MINI_ALU_nx487), .A0 (
          L1_2_L2_1_G1_MINI_ALU_BoothOperand_12), .A1 (
          L1_2_L2_1_G1_MINI_ALU_BoothP_12)) ;
    xor2 L1_2_L2_1_G1_MINI_ALU_ix397 (.Y (L1_2_L2_1_G1_MINI_ALU_nx396), .A0 (
         L1_2_L2_1_G1_MINI_ALU_nx491), .A1 (L1_2_L2_1_G1_MINI_ALU_nx495)) ;
    inv01 L1_2_L2_1_G1_MINI_ALU_ix494 (.Y (L1_2_L2_1_G1_MINI_ALU_nx493), .A (
          L1_2_L2_1_G1_MINI_ALU_BoothP_12)) ;
    xnor2 L1_2_L2_1_G1_MINI_ALU_ix496 (.Y (L1_2_L2_1_G1_MINI_ALU_nx495), .A0 (
          L1_2_L2_1_G1_MINI_ALU_BoothOperand_13), .A1 (
          L1_2_L2_1_G1_MINI_ALU_BoothP_13)) ;
    xor2 L1_2_L2_1_G1_MINI_ALU_ix417 (.Y (L1_2_L2_1_G1_MINI_ALU_nx416), .A0 (
         L1_2_L2_1_G1_MINI_ALU_nx499), .A1 (L1_2_L2_1_G1_MINI_ALU_nx503)) ;
    inv01 L1_2_L2_1_G1_MINI_ALU_ix502 (.Y (L1_2_L2_1_G1_MINI_ALU_nx501), .A (
          L1_2_L2_1_G1_MINI_ALU_BoothP_13)) ;
    xnor2 L1_2_L2_1_G1_MINI_ALU_ix504 (.Y (L1_2_L2_1_G1_MINI_ALU_nx503), .A0 (
          L1_2_L2_1_G1_MINI_ALU_BoothOperand_14), .A1 (
          L1_2_L2_1_G1_MINI_ALU_BoothP_14)) ;
    xor2 L1_2_L2_1_G1_MINI_ALU_ix437 (.Y (L1_2_L2_1_G1_MINI_ALU_nx436), .A0 (
         L1_2_L2_1_G1_MINI_ALU_nx507), .A1 (L1_2_L2_1_G1_MINI_ALU_nx511)) ;
    inv01 L1_2_L2_1_G1_MINI_ALU_ix510 (.Y (L1_2_L2_1_G1_MINI_ALU_nx509), .A (
          L1_2_L2_1_G1_MINI_ALU_BoothP_14)) ;
    xnor2 L1_2_L2_1_G1_MINI_ALU_ix512 (.Y (L1_2_L2_1_G1_MINI_ALU_nx511), .A0 (
          L1_2_L2_1_G1_MINI_ALU_BoothOperand_15), .A1 (
          L1_2_L2_1_G1_MINI_ALU_BoothP_15)) ;
    xnor2 L1_2_L2_1_G1_MINI_ALU_ix457 (.Y (L1_2_L2_1_G1_MINI_ALU_nx456), .A0 (
          L1_2_L2_1_G1_MINI_ALU_nx515), .A1 (L1_2_L2_1_G1_MINI_ALU_nx454)) ;
    inv01 L1_2_L2_1_G1_MINI_ALU_ix518 (.Y (L1_2_L2_1_G1_MINI_ALU_nx517), .A (
          L1_2_L2_1_G1_MINI_ALU_BoothP_15)) ;
    xor2 L1_2_L2_1_G1_MINI_ALU_ix455 (.Y (L1_2_L2_1_G1_MINI_ALU_nx454), .A0 (
         L1_2_L2_1_G1_MINI_ALU_BoothOperand_16), .A1 (
         L1_2_L2_1_G1_MINI_ALU_BoothP_16)) ;
    mux21_ni L1_2_L2_1_G1_MINI_ALU_ix91 (.Y (L1SecondOperands_11__0), .A0 (
             L1_2_L2_1_G1_MINI_ALU_BoothP_1), .A1 (WindowDin_2__1__0), .S0 (
             Instr)) ;
    mux21_ni L1_2_L2_1_G1_MINI_ALU_ix99 (.Y (L1SecondOperands_11__1), .A0 (
             L1_2_L2_1_G1_MINI_ALU_BoothP_2), .A1 (WindowDin_2__1__1), .S0 (
             Instr)) ;
    mux21_ni L1_2_L2_1_G1_MINI_ALU_ix107 (.Y (L1SecondOperands_11__2), .A0 (
             L1_2_L2_1_G1_MINI_ALU_BoothP_3), .A1 (WindowDin_2__1__2), .S0 (
             Instr)) ;
    mux21_ni L1_2_L2_1_G1_MINI_ALU_ix115 (.Y (L1SecondOperands_11__3), .A0 (
             L1_2_L2_1_G1_MINI_ALU_BoothP_4), .A1 (WindowDin_2__1__3), .S0 (
             Instr)) ;
    mux21_ni L1_2_L2_1_G1_MINI_ALU_ix123 (.Y (L1SecondOperands_11__4), .A0 (
             L1_2_L2_1_G1_MINI_ALU_BoothP_5), .A1 (WindowDin_2__1__4), .S0 (
             Instr)) ;
    mux21_ni L1_2_L2_1_G1_MINI_ALU_ix131 (.Y (L1SecondOperands_11__5), .A0 (
             L1_2_L2_1_G1_MINI_ALU_BoothP_6), .A1 (WindowDin_2__1__5), .S0 (
             Instr)) ;
    mux21_ni L1_2_L2_1_G1_MINI_ALU_ix139 (.Y (L1SecondOperands_11__6), .A0 (
             L1_2_L2_1_G1_MINI_ALU_BoothP_7), .A1 (WindowDin_2__1__6), .S0 (
             Instr)) ;
    mux21_ni L1_2_L2_1_G1_MINI_ALU_ix147 (.Y (L1SecondOperands_11__7), .A0 (
             L1_2_L2_1_G1_MINI_ALU_BoothP_8), .A1 (WindowDin_2__1__7), .S0 (
             Instr)) ;
    xor2 L1_2_L2_1_G1_MINI_ALU_ix77 (.Y (L1Results_11__1), .A0 (
         L1_2_L2_1_G1_MINI_ALU_nx529), .A1 (L1_2_L2_1_G1_MINI_ALU_nx531)) ;
    nand02 L1_2_L2_1_G1_MINI_ALU_ix530 (.Y (L1_2_L2_1_G1_MINI_ALU_nx529), .A0 (
           L1SecondOperands_11__0), .A1 (L1FirstOperands_11__0)) ;
    xnor2 L1_2_L2_1_G1_MINI_ALU_ix532 (.Y (L1_2_L2_1_G1_MINI_ALU_nx531), .A0 (
          L1SecondOperands_11__1), .A1 (L1FirstOperands_11__1)) ;
    xor2 L1_2_L2_1_G1_MINI_ALU_ix75 (.Y (L1Results_11__2), .A0 (
         L1_2_L2_1_G1_MINI_ALU_nx534), .A1 (L1_2_L2_1_G1_MINI_ALU_nx537)) ;
    aoi32 L1_2_L2_1_G1_MINI_ALU_ix535 (.Y (L1_2_L2_1_G1_MINI_ALU_nx534), .A0 (
          L1SecondOperands_11__0), .A1 (L1FirstOperands_11__0), .A2 (
          L1_2_L2_1_G1_MINI_ALU_nx30), .B0 (L1FirstOperands_11__1), .B1 (
          L1SecondOperands_11__1)) ;
    xnor2 L1_2_L2_1_G1_MINI_ALU_ix538 (.Y (L1_2_L2_1_G1_MINI_ALU_nx537), .A0 (
          L1SecondOperands_11__2), .A1 (L1FirstOperands_11__2)) ;
    xor2 L1_2_L2_1_G1_MINI_ALU_ix73 (.Y (L1Results_11__3), .A0 (
         L1_2_L2_1_G1_MINI_ALU_nx540), .A1 (L1_2_L2_1_G1_MINI_ALU_nx544)) ;
    aoi22 L1_2_L2_1_G1_MINI_ALU_ix541 (.Y (L1_2_L2_1_G1_MINI_ALU_nx540), .A0 (
          L1FirstOperands_11__2), .A1 (L1SecondOperands_11__2), .B0 (
          L1_2_L2_1_G1_MINI_ALU_nx40), .B1 (L1_2_L2_1_G1_MINI_ALU_nx24)) ;
    xnor2 L1_2_L2_1_G1_MINI_ALU_ix545 (.Y (L1_2_L2_1_G1_MINI_ALU_nx544), .A0 (
          L1SecondOperands_11__3), .A1 (L1FirstOperands_11__3)) ;
    xor2 L1_2_L2_1_G1_MINI_ALU_ix71 (.Y (L1Results_11__4), .A0 (
         L1_2_L2_1_G1_MINI_ALU_nx547), .A1 (L1_2_L2_1_G1_MINI_ALU_nx551)) ;
    aoi22 L1_2_L2_1_G1_MINI_ALU_ix548 (.Y (L1_2_L2_1_G1_MINI_ALU_nx547), .A0 (
          L1FirstOperands_11__3), .A1 (L1SecondOperands_11__3), .B0 (
          L1_2_L2_1_G1_MINI_ALU_nx44), .B1 (L1_2_L2_1_G1_MINI_ALU_nx18)) ;
    xnor2 L1_2_L2_1_G1_MINI_ALU_ix552 (.Y (L1_2_L2_1_G1_MINI_ALU_nx551), .A0 (
          L1SecondOperands_11__4), .A1 (L1FirstOperands_11__4)) ;
    xor2 L1_2_L2_1_G1_MINI_ALU_ix69 (.Y (L1Results_11__5), .A0 (
         L1_2_L2_1_G1_MINI_ALU_nx554), .A1 (L1_2_L2_1_G1_MINI_ALU_nx558)) ;
    aoi22 L1_2_L2_1_G1_MINI_ALU_ix555 (.Y (L1_2_L2_1_G1_MINI_ALU_nx554), .A0 (
          L1FirstOperands_11__4), .A1 (L1SecondOperands_11__4), .B0 (
          L1_2_L2_1_G1_MINI_ALU_nx48), .B1 (L1_2_L2_1_G1_MINI_ALU_nx12)) ;
    xnor2 L1_2_L2_1_G1_MINI_ALU_ix559 (.Y (L1_2_L2_1_G1_MINI_ALU_nx558), .A0 (
          L1SecondOperands_11__5), .A1 (L1FirstOperands_11__5)) ;
    xor2 L1_2_L2_1_G1_MINI_ALU_ix67 (.Y (L1Results_11__6), .A0 (
         L1_2_L2_1_G1_MINI_ALU_nx561), .A1 (L1_2_L2_1_G1_MINI_ALU_nx565)) ;
    aoi22 L1_2_L2_1_G1_MINI_ALU_ix562 (.Y (L1_2_L2_1_G1_MINI_ALU_nx561), .A0 (
          L1FirstOperands_11__5), .A1 (L1SecondOperands_11__5), .B0 (
          L1_2_L2_1_G1_MINI_ALU_nx52), .B1 (L1_2_L2_1_G1_MINI_ALU_nx6)) ;
    xnor2 L1_2_L2_1_G1_MINI_ALU_ix566 (.Y (L1_2_L2_1_G1_MINI_ALU_nx565), .A0 (
          L1SecondOperands_11__6), .A1 (L1FirstOperands_11__6)) ;
    xnor2 L1_2_L2_1_G1_MINI_ALU_ix65 (.Y (L1Results_11__7), .A0 (
          L1_2_L2_1_G1_MINI_ALU_nx568), .A1 (L1_2_L2_1_G1_MINI_ALU_nx62)) ;
    aoi22 L1_2_L2_1_G1_MINI_ALU_ix569 (.Y (L1_2_L2_1_G1_MINI_ALU_nx568), .A0 (
          L1FirstOperands_11__6), .A1 (L1SecondOperands_11__6), .B0 (
          L1_2_L2_1_G1_MINI_ALU_nx56), .B1 (L1_2_L2_1_G1_MINI_ALU_nx0)) ;
    xor2 L1_2_L2_1_G1_MINI_ALU_ix63 (.Y (L1_2_L2_1_G1_MINI_ALU_nx62), .A0 (
         L1SecondOperands_11__7), .A1 (L1FirstOperands_11__7)) ;
    inv01 L1_2_L2_1_G1_MINI_ALU_ix155 (.Y (L1_2_L2_1_G1_MINI_ALU_nx154), .A (
          L1_2_L2_1_G1_MINI_ALU_nx383)) ;
    inv01 L1_2_L2_1_G1_MINI_ALU_ix57 (.Y (L1_2_L2_1_G1_MINI_ALU_nx56), .A (
          L1_2_L2_1_G1_MINI_ALU_nx561)) ;
    inv01 L1_2_L2_1_G1_MINI_ALU_ix53 (.Y (L1_2_L2_1_G1_MINI_ALU_nx52), .A (
          L1_2_L2_1_G1_MINI_ALU_nx554)) ;
    inv01 L1_2_L2_1_G1_MINI_ALU_ix49 (.Y (L1_2_L2_1_G1_MINI_ALU_nx48), .A (
          L1_2_L2_1_G1_MINI_ALU_nx547)) ;
    inv01 L1_2_L2_1_G1_MINI_ALU_ix45 (.Y (L1_2_L2_1_G1_MINI_ALU_nx44), .A (
          L1_2_L2_1_G1_MINI_ALU_nx540)) ;
    inv01 L1_2_L2_1_G1_MINI_ALU_ix41 (.Y (L1_2_L2_1_G1_MINI_ALU_nx40), .A (
          L1_2_L2_1_G1_MINI_ALU_nx534)) ;
    inv01 L1_2_L2_1_G1_MINI_ALU_ix31 (.Y (L1_2_L2_1_G1_MINI_ALU_nx30), .A (
          L1_2_L2_1_G1_MINI_ALU_nx531)) ;
    inv01 L1_2_L2_1_G1_MINI_ALU_ix25 (.Y (L1_2_L2_1_G1_MINI_ALU_nx24), .A (
          L1_2_L2_1_G1_MINI_ALU_nx537)) ;
    inv01 L1_2_L2_1_G1_MINI_ALU_ix19 (.Y (L1_2_L2_1_G1_MINI_ALU_nx18), .A (
          L1_2_L2_1_G1_MINI_ALU_nx544)) ;
    inv01 L1_2_L2_1_G1_MINI_ALU_ix13 (.Y (L1_2_L2_1_G1_MINI_ALU_nx12), .A (
          L1_2_L2_1_G1_MINI_ALU_nx551)) ;
    inv01 L1_2_L2_1_G1_MINI_ALU_ix7 (.Y (L1_2_L2_1_G1_MINI_ALU_nx6), .A (
          L1_2_L2_1_G1_MINI_ALU_nx558)) ;
    inv01 L1_2_L2_1_G1_MINI_ALU_ix1 (.Y (L1_2_L2_1_G1_MINI_ALU_nx0), .A (
          L1_2_L2_1_G1_MINI_ALU_nx565)) ;
    fake_gnd L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix216 (.Y (
             L1_2_L2_1_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    nor02ii L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix81 (.Y (
            L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx80), .A0 (Instr), .A1 (Start)) ;
    aoi21 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix77 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_10), .A0 (
          FilterDin_2__1__1), .A1 (FilterDin_2__1__0), .B0 (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx4)) ;
    nor02_2x L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix5 (.Y (
             L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx4), .A0 (FilterDin_2__1__0), .A1 (
             FilterDin_2__1__1)) ;
    aoi21 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix67 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_11), .A0 (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx328), .A1 (FilterDin_2__1__2), .B0 (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx8)) ;
    nor03_2x L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix9 (.Y (
             L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx8), .A0 (FilterDin_2__1__2), .A1 (
             FilterDin_2__1__0), .A2 (FilterDin_2__1__1)) ;
    xnor2 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix59 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_12), .A0 (
          FilterDin_2__1__3), .A1 (L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx8)) ;
    xnor2 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix51 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_13), .A0 (
          FilterDin_2__1__4), .A1 (L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx12)) ;
    nor04 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix13 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx12), .A0 (FilterDin_2__1__3), .A1 (
          FilterDin_2__1__2), .A2 (FilterDin_2__1__0), .A3 (FilterDin_2__1__1)
          ) ;
    xnor2 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix43 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_14), .A0 (
          FilterDin_2__1__5), .A1 (L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx16)) ;
    nor02ii L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix17 (.Y (
            L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx16), .A0 (FilterDin_2__1__4), .A1 (
            L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx12)) ;
    xnor2 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix35 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_15), .A0 (
          FilterDin_2__1__6), .A1 (L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx20)) ;
    nor02ii L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix21 (.Y (
            L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx20), .A0 (FilterDin_2__1__5), .A1 (
            L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx16)) ;
    xnor2 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix27 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_16), .A0 (
          FilterDin_2__1__7), .A1 (L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx24)) ;
    nor02ii L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix25 (.Y (
            L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx24), .A0 (FilterDin_2__1__6), .A1 (
            L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx20)) ;
    inv01 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix329 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx328), .A (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx4)) ;
    inv02 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix383 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx384), .A (
          L1_2_L2_1_G1_MINI_ALU_BoothP_0)) ;
    dff L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_0 (.Q (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_0), .QB (\$dummy [565]), 
        .D (L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .CLK (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    nor02_2x L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix567 (.Y (
             L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566), .A0 (RST), .A1 (
             L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644)) ;
    dff L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_1 (.Q (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_1), .QB (\$dummy [566]), 
        .D (L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .CLK (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_2 (.Q (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_2), .QB (\$dummy [567]), 
        .D (L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .CLK (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_3 (.Q (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_3), .QB (\$dummy [568]), 
        .D (L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .CLK (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_4 (.Q (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_4), .QB (\$dummy [569]), 
        .D (L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .CLK (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_5 (.Q (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_5), .QB (\$dummy [570]), 
        .D (L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .CLK (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_6 (.Q (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_6), .QB (\$dummy [571]), 
        .D (L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .CLK (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_7 (.Q (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_7), .QB (\$dummy [572]), 
        .D (L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .CLK (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_8 (.Q (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_8), .QB (\$dummy [573]), 
        .D (L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .CLK (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_9 (.Q (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_9), .QB (\$dummy [574]), 
        .D (L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .CLK (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_10 (.Q (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_10), .QB (\$dummy [575])
        , .D (L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .CLK (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_11 (.Q (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_11), .QB (\$dummy [576])
        , .D (L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .CLK (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_12 (.Q (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_12), .QB (\$dummy [577])
        , .D (L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .CLK (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_13 (.Q (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_13), .QB (\$dummy [578])
        , .D (L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .CLK (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_14 (.Q (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_14), .QB (\$dummy [579])
        , .D (L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .CLK (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_15 (.Q (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_15), .QB (\$dummy [580])
        , .D (L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .CLK (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_16 (.Q (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_16), .QB (\$dummy [581])
        , .D (L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .CLK (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    inv02 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix623 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624), .A (CLK)) ;
    inv02 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix625 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626), .A (CLK)) ;
    inv02 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix627 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628), .A (CLK)) ;
    inv02 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix643 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644), .A (nx8058)) ;
    dff L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_0 (.Q (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_0), .QB (\$dummy [582]), 
        .D (L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .CLK (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    nor02_2x L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix567 (.Y (
             L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566), .A0 (RST), .A1 (
             L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644)) ;
    dff L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_1 (.Q (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_1), .QB (\$dummy [583]), 
        .D (L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .CLK (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_2 (.Q (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_2), .QB (\$dummy [584]), 
        .D (L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .CLK (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_3 (.Q (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_3), .QB (\$dummy [585]), 
        .D (L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .CLK (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_4 (.Q (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_4), .QB (\$dummy [586]), 
        .D (L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .CLK (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_5 (.Q (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_5), .QB (\$dummy [587]), 
        .D (L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .CLK (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_6 (.Q (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_6), .QB (\$dummy [588]), 
        .D (L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .CLK (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_7 (.Q (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_7), .QB (\$dummy [589]), 
        .D (L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .CLK (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_8 (.Q (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_8), .QB (\$dummy [590]), 
        .D (L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .CLK (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_9 (.Q (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_9), .QB (\$dummy [591]), 
        .D (L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .CLK (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_10 (.Q (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_10), .QB (\$dummy [592])
        , .D (L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .CLK (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_11 (.Q (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_11), .QB (\$dummy [593])
        , .D (L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .CLK (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_12 (.Q (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_12), .QB (\$dummy [594])
        , .D (L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .CLK (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_13 (.Q (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_13), .QB (\$dummy [595])
        , .D (L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .CLK (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_14 (.Q (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_14), .QB (\$dummy [596])
        , .D (L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .CLK (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_15 (.Q (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_15), .QB (\$dummy [597])
        , .D (L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .CLK (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_16 (.Q (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_16), .QB (\$dummy [598])
        , .D (L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .CLK (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    inv02 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix623 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624), .A (CLK)) ;
    inv02 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix625 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626), .A (CLK)) ;
    inv02 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix627 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628), .A (CLK)) ;
    inv02 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix643 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644), .A (nx8064)) ;
    dff L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_0 (.Q (
        L1_2_L2_1_G1_MINI_ALU_BoothP_0), .QB (\$dummy [599]), .D (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .CLK (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    nor02_2x L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix567 (.Y (
             L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566), .A0 (RST), .A1 (
             L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    dff L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_1 (.Q (
        L1_2_L2_1_G1_MINI_ALU_BoothP_1), .QB (\$dummy [600]), .D (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .CLK (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_2 (.Q (
        L1_2_L2_1_G1_MINI_ALU_BoothP_2), .QB (\$dummy [601]), .D (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .CLK (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_3 (.Q (
        L1_2_L2_1_G1_MINI_ALU_BoothP_3), .QB (\$dummy [602]), .D (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .CLK (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_4 (.Q (
        L1_2_L2_1_G1_MINI_ALU_BoothP_4), .QB (\$dummy [603]), .D (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .CLK (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_5 (.Q (
        L1_2_L2_1_G1_MINI_ALU_BoothP_5), .QB (\$dummy [604]), .D (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .CLK (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_6 (.Q (
        L1_2_L2_1_G1_MINI_ALU_BoothP_6), .QB (\$dummy [605]), .D (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .CLK (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_7 (.Q (
        L1_2_L2_1_G1_MINI_ALU_BoothP_7), .QB (\$dummy [606]), .D (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .CLK (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_8 (.Q (
        L1_2_L2_1_G1_MINI_ALU_BoothP_8), .QB (\$dummy [607]), .D (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .CLK (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_9 (.Q (
        L1_2_L2_1_G1_MINI_ALU_BoothP_9), .QB (\$dummy [608]), .D (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .CLK (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_10 (.Q (
        L1_2_L2_1_G1_MINI_ALU_BoothP_10), .QB (\$dummy [609]), .D (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .CLK (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_11 (.Q (
        L1_2_L2_1_G1_MINI_ALU_BoothP_11), .QB (\$dummy [610]), .D (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .CLK (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_12 (.Q (
        L1_2_L2_1_G1_MINI_ALU_BoothP_12), .QB (\$dummy [611]), .D (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .CLK (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_13 (.Q (
        L1_2_L2_1_G1_MINI_ALU_BoothP_13), .QB (\$dummy [612]), .D (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .CLK (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_14 (.Q (
        L1_2_L2_1_G1_MINI_ALU_BoothP_14), .QB (\$dummy [613]), .D (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .CLK (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_15 (.Q (
        L1_2_L2_1_G1_MINI_ALU_BoothP_15), .QB (\$dummy [614]), .D (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .CLK (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_16 (.Q (
        L1_2_L2_1_G1_MINI_ALU_BoothP_16), .QB (\$dummy [615]), .D (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .CLK (
        L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    inv02 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix623 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624), .A (CLK)) ;
    inv02 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix625 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626), .A (CLK)) ;
    inv02 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix627 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628), .A (CLK)) ;
    inv02 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix643 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644), .A (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642)) ;
    xnor2 L1_2_L2_2_G1_MINI_ALU_ix380 (.Y (L1_2_L2_2_G1_MINI_ALU_nx379), .A0 (
          L1_2_L2_2_G1_MINI_ALU_nx381), .A1 (L1_2_L2_2_G1_MINI_ALU_nx383)) ;
    nand02 L1_2_L2_2_G1_MINI_ALU_ix382 (.Y (L1_2_L2_2_G1_MINI_ALU_nx381), .A0 (
           L1_2_L2_2_G1_MINI_ALU_BoothOperand_0), .A1 (nx8084)) ;
    xnor2 L1_2_L2_2_G1_MINI_ALU_ix384 (.Y (L1_2_L2_2_G1_MINI_ALU_nx383), .A0 (
          L1_2_L2_2_G1_MINI_ALU_BoothOperand_1), .A1 (
          L1_2_L2_2_G1_MINI_ALU_BoothP_1)) ;
    inv01 L1_2_L2_2_G1_MINI_ALU_ix388 (.Y (L1_2_L2_2_G1_MINI_ALU_nx387), .A (
          L1_2_L2_2_G1_MINI_ALU_BoothP_2)) ;
    xnor2 L1_2_L2_2_G1_MINI_ALU_ix390 (.Y (L1_2_L2_2_G1_MINI_ALU_nx389), .A0 (
          L1_2_L2_2_G1_MINI_ALU_nx391), .A1 (L1_2_L2_2_G1_MINI_ALU_nx395)) ;
    aoi32 L1_2_L2_2_G1_MINI_ALU_ix392 (.Y (L1_2_L2_2_G1_MINI_ALU_nx391), .A0 (
          L1_2_L2_2_G1_MINI_ALU_BoothOperand_0), .A1 (nx8084), .A2 (
          L1_2_L2_2_G1_MINI_ALU_nx154), .B0 (L1_2_L2_2_G1_MINI_ALU_BoothP_1), .B1 (
          L1_2_L2_2_G1_MINI_ALU_BoothOperand_1)) ;
    xnor2 L1_2_L2_2_G1_MINI_ALU_ix396 (.Y (L1_2_L2_2_G1_MINI_ALU_nx395), .A0 (
          L1_2_L2_2_G1_MINI_ALU_BoothOperand_2), .A1 (
          L1_2_L2_2_G1_MINI_ALU_BoothP_2)) ;
    inv01 L1_2_L2_2_G1_MINI_ALU_ix400 (.Y (L1_2_L2_2_G1_MINI_ALU_nx399), .A (
          L1_2_L2_2_G1_MINI_ALU_BoothP_3)) ;
    xnor2 L1_2_L2_2_G1_MINI_ALU_ix402 (.Y (L1_2_L2_2_G1_MINI_ALU_nx401), .A0 (
          L1_2_L2_2_G1_MINI_ALU_nx403), .A1 (L1_2_L2_2_G1_MINI_ALU_nx405)) ;
    xnor2 L1_2_L2_2_G1_MINI_ALU_ix406 (.Y (L1_2_L2_2_G1_MINI_ALU_nx405), .A0 (
          L1_2_L2_2_G1_MINI_ALU_BoothOperand_3), .A1 (
          L1_2_L2_2_G1_MINI_ALU_BoothP_3)) ;
    inv01 L1_2_L2_2_G1_MINI_ALU_ix410 (.Y (L1_2_L2_2_G1_MINI_ALU_nx409), .A (
          L1_2_L2_2_G1_MINI_ALU_BoothP_4)) ;
    xnor2 L1_2_L2_2_G1_MINI_ALU_ix412 (.Y (L1_2_L2_2_G1_MINI_ALU_nx411), .A0 (
          L1_2_L2_2_G1_MINI_ALU_nx413), .A1 (L1_2_L2_2_G1_MINI_ALU_nx415)) ;
    xnor2 L1_2_L2_2_G1_MINI_ALU_ix416 (.Y (L1_2_L2_2_G1_MINI_ALU_nx415), .A0 (
          L1_2_L2_2_G1_MINI_ALU_BoothOperand_4), .A1 (
          L1_2_L2_2_G1_MINI_ALU_BoothP_4)) ;
    inv01 L1_2_L2_2_G1_MINI_ALU_ix420 (.Y (L1_2_L2_2_G1_MINI_ALU_nx419), .A (
          L1_2_L2_2_G1_MINI_ALU_BoothP_5)) ;
    xnor2 L1_2_L2_2_G1_MINI_ALU_ix422 (.Y (L1_2_L2_2_G1_MINI_ALU_nx421), .A0 (
          L1_2_L2_2_G1_MINI_ALU_nx423), .A1 (L1_2_L2_2_G1_MINI_ALU_nx425)) ;
    xnor2 L1_2_L2_2_G1_MINI_ALU_ix426 (.Y (L1_2_L2_2_G1_MINI_ALU_nx425), .A0 (
          L1_2_L2_2_G1_MINI_ALU_BoothOperand_5), .A1 (
          L1_2_L2_2_G1_MINI_ALU_BoothP_5)) ;
    inv01 L1_2_L2_2_G1_MINI_ALU_ix430 (.Y (L1_2_L2_2_G1_MINI_ALU_nx429), .A (
          L1_2_L2_2_G1_MINI_ALU_BoothP_6)) ;
    xnor2 L1_2_L2_2_G1_MINI_ALU_ix432 (.Y (L1_2_L2_2_G1_MINI_ALU_nx431), .A0 (
          L1_2_L2_2_G1_MINI_ALU_nx433), .A1 (L1_2_L2_2_G1_MINI_ALU_nx435)) ;
    xnor2 L1_2_L2_2_G1_MINI_ALU_ix436 (.Y (L1_2_L2_2_G1_MINI_ALU_nx435), .A0 (
          L1_2_L2_2_G1_MINI_ALU_BoothOperand_6), .A1 (
          L1_2_L2_2_G1_MINI_ALU_BoothP_6)) ;
    inv01 L1_2_L2_2_G1_MINI_ALU_ix440 (.Y (L1_2_L2_2_G1_MINI_ALU_nx439), .A (
          L1_2_L2_2_G1_MINI_ALU_BoothP_7)) ;
    xnor2 L1_2_L2_2_G1_MINI_ALU_ix442 (.Y (L1_2_L2_2_G1_MINI_ALU_nx441), .A0 (
          L1_2_L2_2_G1_MINI_ALU_nx443), .A1 (L1_2_L2_2_G1_MINI_ALU_nx445)) ;
    xnor2 L1_2_L2_2_G1_MINI_ALU_ix446 (.Y (L1_2_L2_2_G1_MINI_ALU_nx445), .A0 (
          L1_2_L2_2_G1_MINI_ALU_BoothOperand_7), .A1 (
          L1_2_L2_2_G1_MINI_ALU_BoothP_7)) ;
    inv01 L1_2_L2_2_G1_MINI_ALU_ix450 (.Y (L1_2_L2_2_G1_MINI_ALU_nx449), .A (
          L1_2_L2_2_G1_MINI_ALU_BoothP_8)) ;
    xnor2 L1_2_L2_2_G1_MINI_ALU_ix452 (.Y (L1_2_L2_2_G1_MINI_ALU_nx451), .A0 (
          L1_2_L2_2_G1_MINI_ALU_nx453), .A1 (L1_2_L2_2_G1_MINI_ALU_nx455)) ;
    xnor2 L1_2_L2_2_G1_MINI_ALU_ix456 (.Y (L1_2_L2_2_G1_MINI_ALU_nx455), .A0 (
          L1_2_L2_2_G1_MINI_ALU_BoothOperand_8), .A1 (
          L1_2_L2_2_G1_MINI_ALU_BoothP_8)) ;
    xor2 L1_2_L2_2_G1_MINI_ALU_ix317 (.Y (L1_2_L2_2_G1_MINI_ALU_nx316), .A0 (
         L1_2_L2_2_G1_MINI_ALU_nx461), .A1 (L1_2_L2_2_G1_MINI_ALU_nx463)) ;
    xnor2 L1_2_L2_2_G1_MINI_ALU_ix464 (.Y (L1_2_L2_2_G1_MINI_ALU_nx463), .A0 (
          L1_2_L2_2_G1_MINI_ALU_BoothOperand_9), .A1 (
          L1_2_L2_2_G1_MINI_ALU_BoothP_9)) ;
    xor2 L1_2_L2_2_G1_MINI_ALU_ix337 (.Y (L1_2_L2_2_G1_MINI_ALU_nx336), .A0 (
         L1_2_L2_2_G1_MINI_ALU_nx467), .A1 (L1_2_L2_2_G1_MINI_ALU_nx471)) ;
    inv01 L1_2_L2_2_G1_MINI_ALU_ix470 (.Y (L1_2_L2_2_G1_MINI_ALU_nx469), .A (
          L1_2_L2_2_G1_MINI_ALU_BoothP_9)) ;
    xnor2 L1_2_L2_2_G1_MINI_ALU_ix472 (.Y (L1_2_L2_2_G1_MINI_ALU_nx471), .A0 (
          L1_2_L2_2_G1_MINI_ALU_BoothOperand_10), .A1 (
          L1_2_L2_2_G1_MINI_ALU_BoothP_10)) ;
    xor2 L1_2_L2_2_G1_MINI_ALU_ix357 (.Y (L1_2_L2_2_G1_MINI_ALU_nx356), .A0 (
         L1_2_L2_2_G1_MINI_ALU_nx475), .A1 (L1_2_L2_2_G1_MINI_ALU_nx479)) ;
    inv01 L1_2_L2_2_G1_MINI_ALU_ix478 (.Y (L1_2_L2_2_G1_MINI_ALU_nx477), .A (
          L1_2_L2_2_G1_MINI_ALU_BoothP_10)) ;
    xnor2 L1_2_L2_2_G1_MINI_ALU_ix480 (.Y (L1_2_L2_2_G1_MINI_ALU_nx479), .A0 (
          L1_2_L2_2_G1_MINI_ALU_BoothOperand_11), .A1 (
          L1_2_L2_2_G1_MINI_ALU_BoothP_11)) ;
    xor2 L1_2_L2_2_G1_MINI_ALU_ix377 (.Y (L1_2_L2_2_G1_MINI_ALU_nx376), .A0 (
         L1_2_L2_2_G1_MINI_ALU_nx483), .A1 (L1_2_L2_2_G1_MINI_ALU_nx487)) ;
    inv01 L1_2_L2_2_G1_MINI_ALU_ix486 (.Y (L1_2_L2_2_G1_MINI_ALU_nx485), .A (
          L1_2_L2_2_G1_MINI_ALU_BoothP_11)) ;
    xnor2 L1_2_L2_2_G1_MINI_ALU_ix488 (.Y (L1_2_L2_2_G1_MINI_ALU_nx487), .A0 (
          L1_2_L2_2_G1_MINI_ALU_BoothOperand_12), .A1 (
          L1_2_L2_2_G1_MINI_ALU_BoothP_12)) ;
    xor2 L1_2_L2_2_G1_MINI_ALU_ix397 (.Y (L1_2_L2_2_G1_MINI_ALU_nx396), .A0 (
         L1_2_L2_2_G1_MINI_ALU_nx491), .A1 (L1_2_L2_2_G1_MINI_ALU_nx495)) ;
    inv01 L1_2_L2_2_G1_MINI_ALU_ix494 (.Y (L1_2_L2_2_G1_MINI_ALU_nx493), .A (
          L1_2_L2_2_G1_MINI_ALU_BoothP_12)) ;
    xnor2 L1_2_L2_2_G1_MINI_ALU_ix496 (.Y (L1_2_L2_2_G1_MINI_ALU_nx495), .A0 (
          L1_2_L2_2_G1_MINI_ALU_BoothOperand_13), .A1 (
          L1_2_L2_2_G1_MINI_ALU_BoothP_13)) ;
    xor2 L1_2_L2_2_G1_MINI_ALU_ix417 (.Y (L1_2_L2_2_G1_MINI_ALU_nx416), .A0 (
         L1_2_L2_2_G1_MINI_ALU_nx499), .A1 (L1_2_L2_2_G1_MINI_ALU_nx503)) ;
    inv01 L1_2_L2_2_G1_MINI_ALU_ix502 (.Y (L1_2_L2_2_G1_MINI_ALU_nx501), .A (
          L1_2_L2_2_G1_MINI_ALU_BoothP_13)) ;
    xnor2 L1_2_L2_2_G1_MINI_ALU_ix504 (.Y (L1_2_L2_2_G1_MINI_ALU_nx503), .A0 (
          L1_2_L2_2_G1_MINI_ALU_BoothOperand_14), .A1 (
          L1_2_L2_2_G1_MINI_ALU_BoothP_14)) ;
    xor2 L1_2_L2_2_G1_MINI_ALU_ix437 (.Y (L1_2_L2_2_G1_MINI_ALU_nx436), .A0 (
         L1_2_L2_2_G1_MINI_ALU_nx507), .A1 (L1_2_L2_2_G1_MINI_ALU_nx511)) ;
    inv01 L1_2_L2_2_G1_MINI_ALU_ix510 (.Y (L1_2_L2_2_G1_MINI_ALU_nx509), .A (
          L1_2_L2_2_G1_MINI_ALU_BoothP_14)) ;
    xnor2 L1_2_L2_2_G1_MINI_ALU_ix512 (.Y (L1_2_L2_2_G1_MINI_ALU_nx511), .A0 (
          L1_2_L2_2_G1_MINI_ALU_BoothOperand_15), .A1 (
          L1_2_L2_2_G1_MINI_ALU_BoothP_15)) ;
    xnor2 L1_2_L2_2_G1_MINI_ALU_ix457 (.Y (L1_2_L2_2_G1_MINI_ALU_nx456), .A0 (
          L1_2_L2_2_G1_MINI_ALU_nx515), .A1 (L1_2_L2_2_G1_MINI_ALU_nx454)) ;
    inv01 L1_2_L2_2_G1_MINI_ALU_ix518 (.Y (L1_2_L2_2_G1_MINI_ALU_nx517), .A (
          L1_2_L2_2_G1_MINI_ALU_BoothP_15)) ;
    xor2 L1_2_L2_2_G1_MINI_ALU_ix455 (.Y (L1_2_L2_2_G1_MINI_ALU_nx454), .A0 (
         L1_2_L2_2_G1_MINI_ALU_BoothOperand_16), .A1 (
         L1_2_L2_2_G1_MINI_ALU_BoothP_16)) ;
    mux21_ni L1_2_L2_2_G1_MINI_ALU_ix91 (.Y (L1FirstOperands_11__0), .A0 (
             L1_2_L2_2_G1_MINI_ALU_BoothP_1), .A1 (WindowDin_2__2__0), .S0 (
             Instr)) ;
    mux21_ni L1_2_L2_2_G1_MINI_ALU_ix99 (.Y (L1FirstOperands_11__1), .A0 (
             L1_2_L2_2_G1_MINI_ALU_BoothP_2), .A1 (WindowDin_2__2__1), .S0 (
             Instr)) ;
    mux21_ni L1_2_L2_2_G1_MINI_ALU_ix107 (.Y (L1FirstOperands_11__2), .A0 (
             L1_2_L2_2_G1_MINI_ALU_BoothP_3), .A1 (WindowDin_2__2__2), .S0 (
             Instr)) ;
    mux21_ni L1_2_L2_2_G1_MINI_ALU_ix115 (.Y (L1FirstOperands_11__3), .A0 (
             L1_2_L2_2_G1_MINI_ALU_BoothP_4), .A1 (WindowDin_2__2__3), .S0 (
             Instr)) ;
    mux21_ni L1_2_L2_2_G1_MINI_ALU_ix123 (.Y (L1FirstOperands_11__4), .A0 (
             L1_2_L2_2_G1_MINI_ALU_BoothP_5), .A1 (WindowDin_2__2__4), .S0 (
             Instr)) ;
    mux21_ni L1_2_L2_2_G1_MINI_ALU_ix131 (.Y (L1FirstOperands_11__5), .A0 (
             L1_2_L2_2_G1_MINI_ALU_BoothP_6), .A1 (WindowDin_2__2__5), .S0 (
             Instr)) ;
    mux21_ni L1_2_L2_2_G1_MINI_ALU_ix139 (.Y (L1FirstOperands_11__6), .A0 (
             L1_2_L2_2_G1_MINI_ALU_BoothP_7), .A1 (WindowDin_2__2__6), .S0 (
             Instr)) ;
    mux21_ni L1_2_L2_2_G1_MINI_ALU_ix147 (.Y (L1FirstOperands_11__7), .A0 (
             L1_2_L2_2_G1_MINI_ALU_BoothP_8), .A1 (WindowDin_2__2__7), .S0 (
             Instr)) ;
    inv01 L1_2_L2_2_G1_MINI_ALU_ix155 (.Y (L1_2_L2_2_G1_MINI_ALU_nx154), .A (
          L1_2_L2_2_G1_MINI_ALU_nx383)) ;
    fake_gnd L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix216 (.Y (
             L1_2_L2_2_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    nor02ii L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix81 (.Y (
            L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx80), .A0 (Instr), .A1 (Start)) ;
    aoi21 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix77 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_10), .A0 (
          FilterDin_2__2__1), .A1 (FilterDin_2__2__0), .B0 (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx4)) ;
    nor02_2x L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix5 (.Y (
             L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx4), .A0 (FilterDin_2__2__0), .A1 (
             FilterDin_2__2__1)) ;
    aoi21 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix67 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_11), .A0 (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx328), .A1 (FilterDin_2__2__2), .B0 (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx8)) ;
    nor03_2x L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix9 (.Y (
             L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx8), .A0 (FilterDin_2__2__2), .A1 (
             FilterDin_2__2__0), .A2 (FilterDin_2__2__1)) ;
    xnor2 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix59 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_12), .A0 (
          FilterDin_2__2__3), .A1 (L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx8)) ;
    xnor2 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix51 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_13), .A0 (
          FilterDin_2__2__4), .A1 (L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx12)) ;
    nor04 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix13 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx12), .A0 (FilterDin_2__2__3), .A1 (
          FilterDin_2__2__2), .A2 (FilterDin_2__2__0), .A3 (FilterDin_2__2__1)
          ) ;
    xnor2 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix43 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_14), .A0 (
          FilterDin_2__2__5), .A1 (L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx16)) ;
    nor02ii L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix17 (.Y (
            L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx16), .A0 (FilterDin_2__2__4), .A1 (
            L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx12)) ;
    xnor2 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix35 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_15), .A0 (
          FilterDin_2__2__6), .A1 (L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx20)) ;
    nor02ii L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix21 (.Y (
            L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx20), .A0 (FilterDin_2__2__5), .A1 (
            L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx16)) ;
    xnor2 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix27 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_16), .A0 (
          FilterDin_2__2__7), .A1 (L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx24)) ;
    nor02ii L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix25 (.Y (
            L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx24), .A0 (FilterDin_2__2__6), .A1 (
            L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx20)) ;
    inv01 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix329 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx328), .A (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx4)) ;
    inv02 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix383 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx384), .A (
          L1_2_L2_2_G1_MINI_ALU_BoothP_0)) ;
    dff L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_0 (.Q (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_0), .QB (\$dummy [616]), 
        .D (L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .CLK (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    nor02_2x L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix567 (.Y (
             L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566), .A0 (RST), .A1 (
             L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644)) ;
    dff L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_1 (.Q (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_1), .QB (\$dummy [617]), 
        .D (L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .CLK (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_2 (.Q (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_2), .QB (\$dummy [618]), 
        .D (L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .CLK (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_3 (.Q (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_3), .QB (\$dummy [619]), 
        .D (L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .CLK (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_4 (.Q (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_4), .QB (\$dummy [620]), 
        .D (L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .CLK (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_5 (.Q (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_5), .QB (\$dummy [621]), 
        .D (L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .CLK (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_6 (.Q (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_6), .QB (\$dummy [622]), 
        .D (L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .CLK (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_7 (.Q (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_7), .QB (\$dummy [623]), 
        .D (L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .CLK (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_8 (.Q (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_8), .QB (\$dummy [624]), 
        .D (L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .CLK (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_9 (.Q (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_9), .QB (\$dummy [625]), 
        .D (L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .CLK (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_10 (.Q (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_10), .QB (\$dummy [626])
        , .D (L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .CLK (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_11 (.Q (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_11), .QB (\$dummy [627])
        , .D (L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .CLK (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_12 (.Q (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_12), .QB (\$dummy [628])
        , .D (L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .CLK (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_13 (.Q (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_13), .QB (\$dummy [629])
        , .D (L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .CLK (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_14 (.Q (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_14), .QB (\$dummy [630])
        , .D (L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .CLK (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_15 (.Q (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_15), .QB (\$dummy [631])
        , .D (L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .CLK (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_16 (.Q (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_16), .QB (\$dummy [632])
        , .D (L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .CLK (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    inv02 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix623 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624), .A (CLK)) ;
    inv02 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix625 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626), .A (CLK)) ;
    inv02 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix627 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628), .A (CLK)) ;
    inv02 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix643 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644), .A (nx8098)) ;
    dff L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_0 (.Q (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_0), .QB (\$dummy [633]), 
        .D (L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .CLK (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    nor02_2x L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix567 (.Y (
             L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566), .A0 (RST), .A1 (
             L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644)) ;
    dff L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_1 (.Q (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_1), .QB (\$dummy [634]), 
        .D (L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .CLK (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_2 (.Q (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_2), .QB (\$dummy [635]), 
        .D (L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .CLK (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_3 (.Q (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_3), .QB (\$dummy [636]), 
        .D (L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .CLK (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_4 (.Q (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_4), .QB (\$dummy [637]), 
        .D (L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .CLK (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_5 (.Q (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_5), .QB (\$dummy [638]), 
        .D (L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .CLK (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_6 (.Q (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_6), .QB (\$dummy [639]), 
        .D (L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .CLK (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_7 (.Q (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_7), .QB (\$dummy [640]), 
        .D (L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .CLK (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_8 (.Q (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_8), .QB (\$dummy [641]), 
        .D (L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .CLK (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_9 (.Q (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_9), .QB (\$dummy [642]), 
        .D (L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .CLK (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_10 (.Q (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_10), .QB (\$dummy [643])
        , .D (L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .CLK (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_11 (.Q (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_11), .QB (\$dummy [644])
        , .D (L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .CLK (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_12 (.Q (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_12), .QB (\$dummy [645])
        , .D (L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .CLK (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_13 (.Q (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_13), .QB (\$dummy [646])
        , .D (L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .CLK (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_14 (.Q (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_14), .QB (\$dummy [647])
        , .D (L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .CLK (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_15 (.Q (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_15), .QB (\$dummy [648])
        , .D (L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .CLK (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_16 (.Q (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_16), .QB (\$dummy [649])
        , .D (L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .CLK (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    inv02 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix623 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624), .A (CLK)) ;
    inv02 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix625 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626), .A (CLK)) ;
    inv02 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix627 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628), .A (CLK)) ;
    inv02 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix643 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644), .A (nx8104)) ;
    dff L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_0 (.Q (
        L1_2_L2_2_G1_MINI_ALU_BoothP_0), .QB (\$dummy [650]), .D (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .CLK (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    nor02_2x L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix567 (.Y (
             L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566), .A0 (RST), .A1 (
             L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    dff L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_1 (.Q (
        L1_2_L2_2_G1_MINI_ALU_BoothP_1), .QB (\$dummy [651]), .D (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .CLK (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_2 (.Q (
        L1_2_L2_2_G1_MINI_ALU_BoothP_2), .QB (\$dummy [652]), .D (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .CLK (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_3 (.Q (
        L1_2_L2_2_G1_MINI_ALU_BoothP_3), .QB (\$dummy [653]), .D (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .CLK (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_4 (.Q (
        L1_2_L2_2_G1_MINI_ALU_BoothP_4), .QB (\$dummy [654]), .D (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .CLK (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_5 (.Q (
        L1_2_L2_2_G1_MINI_ALU_BoothP_5), .QB (\$dummy [655]), .D (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .CLK (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_6 (.Q (
        L1_2_L2_2_G1_MINI_ALU_BoothP_6), .QB (\$dummy [656]), .D (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .CLK (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_7 (.Q (
        L1_2_L2_2_G1_MINI_ALU_BoothP_7), .QB (\$dummy [657]), .D (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .CLK (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_8 (.Q (
        L1_2_L2_2_G1_MINI_ALU_BoothP_8), .QB (\$dummy [658]), .D (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .CLK (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_9 (.Q (
        L1_2_L2_2_G1_MINI_ALU_BoothP_9), .QB (\$dummy [659]), .D (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .CLK (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_10 (.Q (
        L1_2_L2_2_G1_MINI_ALU_BoothP_10), .QB (\$dummy [660]), .D (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .CLK (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_11 (.Q (
        L1_2_L2_2_G1_MINI_ALU_BoothP_11), .QB (\$dummy [661]), .D (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .CLK (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_12 (.Q (
        L1_2_L2_2_G1_MINI_ALU_BoothP_12), .QB (\$dummy [662]), .D (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .CLK (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_13 (.Q (
        L1_2_L2_2_G1_MINI_ALU_BoothP_13), .QB (\$dummy [663]), .D (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .CLK (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_14 (.Q (
        L1_2_L2_2_G1_MINI_ALU_BoothP_14), .QB (\$dummy [664]), .D (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .CLK (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_15 (.Q (
        L1_2_L2_2_G1_MINI_ALU_BoothP_15), .QB (\$dummy [665]), .D (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .CLK (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_16 (.Q (
        L1_2_L2_2_G1_MINI_ALU_BoothP_16), .QB (\$dummy [666]), .D (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .CLK (
        L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    inv02 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix623 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624), .A (CLK)) ;
    inv02 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix625 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626), .A (CLK)) ;
    inv02 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix627 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628), .A (CLK)) ;
    inv02 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix643 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644), .A (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642)) ;
    xor2 L1_2_L2_3_G2_MINI_ALU_ix83 (.Y (L2Results_0__0), .A0 (L1Results_1__0), 
         .A1 (L1Results_0__0)) ;
    xnor2 L1_2_L2_3_G2_MINI_ALU_ix380 (.Y (L1_2_L2_3_G2_MINI_ALU_nx379), .A0 (
          L1_2_L2_3_G2_MINI_ALU_nx381), .A1 (L1_2_L2_3_G2_MINI_ALU_nx383)) ;
    nand02 L1_2_L2_3_G2_MINI_ALU_ix382 (.Y (L1_2_L2_3_G2_MINI_ALU_nx381), .A0 (
           L1_2_L2_3_G2_MINI_ALU_BoothOperand_0), .A1 (nx8124)) ;
    xnor2 L1_2_L2_3_G2_MINI_ALU_ix384 (.Y (L1_2_L2_3_G2_MINI_ALU_nx383), .A0 (
          L1_2_L2_3_G2_MINI_ALU_BoothOperand_1), .A1 (
          L1_2_L2_3_G2_MINI_ALU_BoothP_1)) ;
    inv01 L1_2_L2_3_G2_MINI_ALU_ix388 (.Y (L1_2_L2_3_G2_MINI_ALU_nx387), .A (
          L1_2_L2_3_G2_MINI_ALU_BoothP_2)) ;
    xnor2 L1_2_L2_3_G2_MINI_ALU_ix390 (.Y (L1_2_L2_3_G2_MINI_ALU_nx389), .A0 (
          L1_2_L2_3_G2_MINI_ALU_nx391), .A1 (L1_2_L2_3_G2_MINI_ALU_nx395)) ;
    aoi32 L1_2_L2_3_G2_MINI_ALU_ix392 (.Y (L1_2_L2_3_G2_MINI_ALU_nx391), .A0 (
          L1_2_L2_3_G2_MINI_ALU_BoothOperand_0), .A1 (nx8124), .A2 (
          L1_2_L2_3_G2_MINI_ALU_nx154), .B0 (L1_2_L2_3_G2_MINI_ALU_BoothP_1), .B1 (
          L1_2_L2_3_G2_MINI_ALU_BoothOperand_1)) ;
    xnor2 L1_2_L2_3_G2_MINI_ALU_ix396 (.Y (L1_2_L2_3_G2_MINI_ALU_nx395), .A0 (
          L1_2_L2_3_G2_MINI_ALU_BoothOperand_2), .A1 (
          L1_2_L2_3_G2_MINI_ALU_BoothP_2)) ;
    inv01 L1_2_L2_3_G2_MINI_ALU_ix400 (.Y (L1_2_L2_3_G2_MINI_ALU_nx399), .A (
          L1_2_L2_3_G2_MINI_ALU_BoothP_3)) ;
    xnor2 L1_2_L2_3_G2_MINI_ALU_ix402 (.Y (L1_2_L2_3_G2_MINI_ALU_nx401), .A0 (
          L1_2_L2_3_G2_MINI_ALU_nx403), .A1 (L1_2_L2_3_G2_MINI_ALU_nx405)) ;
    xnor2 L1_2_L2_3_G2_MINI_ALU_ix406 (.Y (L1_2_L2_3_G2_MINI_ALU_nx405), .A0 (
          L1_2_L2_3_G2_MINI_ALU_BoothOperand_3), .A1 (
          L1_2_L2_3_G2_MINI_ALU_BoothP_3)) ;
    inv01 L1_2_L2_3_G2_MINI_ALU_ix410 (.Y (L1_2_L2_3_G2_MINI_ALU_nx409), .A (
          L1_2_L2_3_G2_MINI_ALU_BoothP_4)) ;
    xnor2 L1_2_L2_3_G2_MINI_ALU_ix412 (.Y (L1_2_L2_3_G2_MINI_ALU_nx411), .A0 (
          L1_2_L2_3_G2_MINI_ALU_nx413), .A1 (L1_2_L2_3_G2_MINI_ALU_nx415)) ;
    xnor2 L1_2_L2_3_G2_MINI_ALU_ix416 (.Y (L1_2_L2_3_G2_MINI_ALU_nx415), .A0 (
          L1_2_L2_3_G2_MINI_ALU_BoothOperand_4), .A1 (
          L1_2_L2_3_G2_MINI_ALU_BoothP_4)) ;
    inv01 L1_2_L2_3_G2_MINI_ALU_ix420 (.Y (L1_2_L2_3_G2_MINI_ALU_nx419), .A (
          L1_2_L2_3_G2_MINI_ALU_BoothP_5)) ;
    xnor2 L1_2_L2_3_G2_MINI_ALU_ix422 (.Y (L1_2_L2_3_G2_MINI_ALU_nx421), .A0 (
          L1_2_L2_3_G2_MINI_ALU_nx423), .A1 (L1_2_L2_3_G2_MINI_ALU_nx425)) ;
    xnor2 L1_2_L2_3_G2_MINI_ALU_ix426 (.Y (L1_2_L2_3_G2_MINI_ALU_nx425), .A0 (
          L1_2_L2_3_G2_MINI_ALU_BoothOperand_5), .A1 (
          L1_2_L2_3_G2_MINI_ALU_BoothP_5)) ;
    inv01 L1_2_L2_3_G2_MINI_ALU_ix430 (.Y (L1_2_L2_3_G2_MINI_ALU_nx429), .A (
          L1_2_L2_3_G2_MINI_ALU_BoothP_6)) ;
    xnor2 L1_2_L2_3_G2_MINI_ALU_ix432 (.Y (L1_2_L2_3_G2_MINI_ALU_nx431), .A0 (
          L1_2_L2_3_G2_MINI_ALU_nx433), .A1 (L1_2_L2_3_G2_MINI_ALU_nx435)) ;
    xnor2 L1_2_L2_3_G2_MINI_ALU_ix436 (.Y (L1_2_L2_3_G2_MINI_ALU_nx435), .A0 (
          L1_2_L2_3_G2_MINI_ALU_BoothOperand_6), .A1 (
          L1_2_L2_3_G2_MINI_ALU_BoothP_6)) ;
    inv01 L1_2_L2_3_G2_MINI_ALU_ix440 (.Y (L1_2_L2_3_G2_MINI_ALU_nx439), .A (
          L1_2_L2_3_G2_MINI_ALU_BoothP_7)) ;
    xnor2 L1_2_L2_3_G2_MINI_ALU_ix442 (.Y (L1_2_L2_3_G2_MINI_ALU_nx441), .A0 (
          L1_2_L2_3_G2_MINI_ALU_nx443), .A1 (L1_2_L2_3_G2_MINI_ALU_nx445)) ;
    xnor2 L1_2_L2_3_G2_MINI_ALU_ix446 (.Y (L1_2_L2_3_G2_MINI_ALU_nx445), .A0 (
          L1_2_L2_3_G2_MINI_ALU_BoothOperand_7), .A1 (
          L1_2_L2_3_G2_MINI_ALU_BoothP_7)) ;
    inv01 L1_2_L2_3_G2_MINI_ALU_ix450 (.Y (L1_2_L2_3_G2_MINI_ALU_nx449), .A (
          L1_2_L2_3_G2_MINI_ALU_BoothP_8)) ;
    xnor2 L1_2_L2_3_G2_MINI_ALU_ix452 (.Y (L1_2_L2_3_G2_MINI_ALU_nx451), .A0 (
          L1_2_L2_3_G2_MINI_ALU_nx453), .A1 (L1_2_L2_3_G2_MINI_ALU_nx455)) ;
    xnor2 L1_2_L2_3_G2_MINI_ALU_ix456 (.Y (L1_2_L2_3_G2_MINI_ALU_nx455), .A0 (
          L1_2_L2_3_G2_MINI_ALU_BoothOperand_8), .A1 (
          L1_2_L2_3_G2_MINI_ALU_BoothP_8)) ;
    xor2 L1_2_L2_3_G2_MINI_ALU_ix317 (.Y (L1_2_L2_3_G2_MINI_ALU_nx316), .A0 (
         L1_2_L2_3_G2_MINI_ALU_nx461), .A1 (L1_2_L2_3_G2_MINI_ALU_nx463)) ;
    xnor2 L1_2_L2_3_G2_MINI_ALU_ix464 (.Y (L1_2_L2_3_G2_MINI_ALU_nx463), .A0 (
          L1_2_L2_3_G2_MINI_ALU_BoothOperand_9), .A1 (
          L1_2_L2_3_G2_MINI_ALU_BoothP_9)) ;
    xor2 L1_2_L2_3_G2_MINI_ALU_ix337 (.Y (L1_2_L2_3_G2_MINI_ALU_nx336), .A0 (
         L1_2_L2_3_G2_MINI_ALU_nx467), .A1 (L1_2_L2_3_G2_MINI_ALU_nx471)) ;
    inv01 L1_2_L2_3_G2_MINI_ALU_ix470 (.Y (L1_2_L2_3_G2_MINI_ALU_nx469), .A (
          L1_2_L2_3_G2_MINI_ALU_BoothP_9)) ;
    xnor2 L1_2_L2_3_G2_MINI_ALU_ix472 (.Y (L1_2_L2_3_G2_MINI_ALU_nx471), .A0 (
          L1_2_L2_3_G2_MINI_ALU_BoothOperand_10), .A1 (
          L1_2_L2_3_G2_MINI_ALU_BoothP_10)) ;
    xor2 L1_2_L2_3_G2_MINI_ALU_ix357 (.Y (L1_2_L2_3_G2_MINI_ALU_nx356), .A0 (
         L1_2_L2_3_G2_MINI_ALU_nx475), .A1 (L1_2_L2_3_G2_MINI_ALU_nx479)) ;
    inv01 L1_2_L2_3_G2_MINI_ALU_ix478 (.Y (L1_2_L2_3_G2_MINI_ALU_nx477), .A (
          L1_2_L2_3_G2_MINI_ALU_BoothP_10)) ;
    xnor2 L1_2_L2_3_G2_MINI_ALU_ix480 (.Y (L1_2_L2_3_G2_MINI_ALU_nx479), .A0 (
          L1_2_L2_3_G2_MINI_ALU_BoothOperand_11), .A1 (
          L1_2_L2_3_G2_MINI_ALU_BoothP_11)) ;
    xor2 L1_2_L2_3_G2_MINI_ALU_ix377 (.Y (L1_2_L2_3_G2_MINI_ALU_nx376), .A0 (
         L1_2_L2_3_G2_MINI_ALU_nx483), .A1 (L1_2_L2_3_G2_MINI_ALU_nx487)) ;
    inv01 L1_2_L2_3_G2_MINI_ALU_ix486 (.Y (L1_2_L2_3_G2_MINI_ALU_nx485), .A (
          L1_2_L2_3_G2_MINI_ALU_BoothP_11)) ;
    xnor2 L1_2_L2_3_G2_MINI_ALU_ix488 (.Y (L1_2_L2_3_G2_MINI_ALU_nx487), .A0 (
          L1_2_L2_3_G2_MINI_ALU_BoothOperand_12), .A1 (
          L1_2_L2_3_G2_MINI_ALU_BoothP_12)) ;
    xor2 L1_2_L2_3_G2_MINI_ALU_ix397 (.Y (L1_2_L2_3_G2_MINI_ALU_nx396), .A0 (
         L1_2_L2_3_G2_MINI_ALU_nx491), .A1 (L1_2_L2_3_G2_MINI_ALU_nx495)) ;
    inv01 L1_2_L2_3_G2_MINI_ALU_ix494 (.Y (L1_2_L2_3_G2_MINI_ALU_nx493), .A (
          L1_2_L2_3_G2_MINI_ALU_BoothP_12)) ;
    xnor2 L1_2_L2_3_G2_MINI_ALU_ix496 (.Y (L1_2_L2_3_G2_MINI_ALU_nx495), .A0 (
          L1_2_L2_3_G2_MINI_ALU_BoothOperand_13), .A1 (
          L1_2_L2_3_G2_MINI_ALU_BoothP_13)) ;
    xor2 L1_2_L2_3_G2_MINI_ALU_ix417 (.Y (L1_2_L2_3_G2_MINI_ALU_nx416), .A0 (
         L1_2_L2_3_G2_MINI_ALU_nx499), .A1 (L1_2_L2_3_G2_MINI_ALU_nx503)) ;
    inv01 L1_2_L2_3_G2_MINI_ALU_ix502 (.Y (L1_2_L2_3_G2_MINI_ALU_nx501), .A (
          L1_2_L2_3_G2_MINI_ALU_BoothP_13)) ;
    xnor2 L1_2_L2_3_G2_MINI_ALU_ix504 (.Y (L1_2_L2_3_G2_MINI_ALU_nx503), .A0 (
          L1_2_L2_3_G2_MINI_ALU_BoothOperand_14), .A1 (
          L1_2_L2_3_G2_MINI_ALU_BoothP_14)) ;
    xor2 L1_2_L2_3_G2_MINI_ALU_ix437 (.Y (L1_2_L2_3_G2_MINI_ALU_nx436), .A0 (
         L1_2_L2_3_G2_MINI_ALU_nx507), .A1 (L1_2_L2_3_G2_MINI_ALU_nx511)) ;
    inv01 L1_2_L2_3_G2_MINI_ALU_ix510 (.Y (L1_2_L2_3_G2_MINI_ALU_nx509), .A (
          L1_2_L2_3_G2_MINI_ALU_BoothP_14)) ;
    xnor2 L1_2_L2_3_G2_MINI_ALU_ix512 (.Y (L1_2_L2_3_G2_MINI_ALU_nx511), .A0 (
          L1_2_L2_3_G2_MINI_ALU_BoothOperand_15), .A1 (
          L1_2_L2_3_G2_MINI_ALU_BoothP_15)) ;
    xnor2 L1_2_L2_3_G2_MINI_ALU_ix457 (.Y (L1_2_L2_3_G2_MINI_ALU_nx456), .A0 (
          L1_2_L2_3_G2_MINI_ALU_nx515), .A1 (L1_2_L2_3_G2_MINI_ALU_nx454)) ;
    inv01 L1_2_L2_3_G2_MINI_ALU_ix518 (.Y (L1_2_L2_3_G2_MINI_ALU_nx517), .A (
          L1_2_L2_3_G2_MINI_ALU_BoothP_15)) ;
    xor2 L1_2_L2_3_G2_MINI_ALU_ix455 (.Y (L1_2_L2_3_G2_MINI_ALU_nx454), .A0 (
         L1_2_L2_3_G2_MINI_ALU_BoothOperand_16), .A1 (
         L1_2_L2_3_G2_MINI_ALU_BoothP_16)) ;
    mux21_ni L1_2_L2_3_G2_MINI_ALU_ix91 (.Y (L1FirstOperands_0__0), .A0 (
             L1_2_L2_3_G2_MINI_ALU_BoothP_1), .A1 (WindowDin_2__3__0), .S0 (
             Instr)) ;
    mux21_ni L1_2_L2_3_G2_MINI_ALU_ix99 (.Y (L1FirstOperands_0__1), .A0 (
             L1_2_L2_3_G2_MINI_ALU_BoothP_2), .A1 (WindowDin_2__3__1), .S0 (
             Instr)) ;
    mux21_ni L1_2_L2_3_G2_MINI_ALU_ix107 (.Y (L1FirstOperands_0__2), .A0 (
             L1_2_L2_3_G2_MINI_ALU_BoothP_3), .A1 (WindowDin_2__3__2), .S0 (
             Instr)) ;
    mux21_ni L1_2_L2_3_G2_MINI_ALU_ix115 (.Y (L1FirstOperands_0__3), .A0 (
             L1_2_L2_3_G2_MINI_ALU_BoothP_4), .A1 (WindowDin_2__3__3), .S0 (
             Instr)) ;
    mux21_ni L1_2_L2_3_G2_MINI_ALU_ix123 (.Y (L1FirstOperands_0__4), .A0 (
             L1_2_L2_3_G2_MINI_ALU_BoothP_5), .A1 (WindowDin_2__3__4), .S0 (
             Instr)) ;
    mux21_ni L1_2_L2_3_G2_MINI_ALU_ix131 (.Y (L1FirstOperands_0__5), .A0 (
             L1_2_L2_3_G2_MINI_ALU_BoothP_6), .A1 (WindowDin_2__3__5), .S0 (
             Instr)) ;
    mux21_ni L1_2_L2_3_G2_MINI_ALU_ix139 (.Y (L1FirstOperands_0__6), .A0 (
             L1_2_L2_3_G2_MINI_ALU_BoothP_7), .A1 (WindowDin_2__3__6), .S0 (
             Instr)) ;
    mux21_ni L1_2_L2_3_G2_MINI_ALU_ix147 (.Y (L1FirstOperands_0__7), .A0 (
             L1_2_L2_3_G2_MINI_ALU_BoothP_8), .A1 (WindowDin_2__3__7), .S0 (
             Instr)) ;
    xor2 L1_2_L2_3_G2_MINI_ALU_ix77 (.Y (L2Results_0__1), .A0 (
         L1_2_L2_3_G2_MINI_ALU_nx529), .A1 (L1_2_L2_3_G2_MINI_ALU_nx531)) ;
    nand02 L1_2_L2_3_G2_MINI_ALU_ix530 (.Y (L1_2_L2_3_G2_MINI_ALU_nx529), .A0 (
           L1Results_1__0), .A1 (L1Results_0__0)) ;
    xnor2 L1_2_L2_3_G2_MINI_ALU_ix532 (.Y (L1_2_L2_3_G2_MINI_ALU_nx531), .A0 (
          L1Results_1__1), .A1 (L1Results_0__1)) ;
    xor2 L1_2_L2_3_G2_MINI_ALU_ix75 (.Y (L2Results_0__2), .A0 (
         L1_2_L2_3_G2_MINI_ALU_nx534), .A1 (L1_2_L2_3_G2_MINI_ALU_nx537)) ;
    aoi32 L1_2_L2_3_G2_MINI_ALU_ix535 (.Y (L1_2_L2_3_G2_MINI_ALU_nx534), .A0 (
          L1Results_1__0), .A1 (L1Results_0__0), .A2 (L1_2_L2_3_G2_MINI_ALU_nx30
          ), .B0 (L1Results_0__1), .B1 (L1Results_1__1)) ;
    xnor2 L1_2_L2_3_G2_MINI_ALU_ix538 (.Y (L1_2_L2_3_G2_MINI_ALU_nx537), .A0 (
          L1Results_1__2), .A1 (L1Results_0__2)) ;
    xor2 L1_2_L2_3_G2_MINI_ALU_ix73 (.Y (L2Results_0__3), .A0 (
         L1_2_L2_3_G2_MINI_ALU_nx540), .A1 (L1_2_L2_3_G2_MINI_ALU_nx544)) ;
    aoi22 L1_2_L2_3_G2_MINI_ALU_ix541 (.Y (L1_2_L2_3_G2_MINI_ALU_nx540), .A0 (
          L1Results_0__2), .A1 (L1Results_1__2), .B0 (L1_2_L2_3_G2_MINI_ALU_nx40
          ), .B1 (L1_2_L2_3_G2_MINI_ALU_nx24)) ;
    xnor2 L1_2_L2_3_G2_MINI_ALU_ix545 (.Y (L1_2_L2_3_G2_MINI_ALU_nx544), .A0 (
          L1Results_1__3), .A1 (L1Results_0__3)) ;
    xor2 L1_2_L2_3_G2_MINI_ALU_ix71 (.Y (L2Results_0__4), .A0 (
         L1_2_L2_3_G2_MINI_ALU_nx547), .A1 (L1_2_L2_3_G2_MINI_ALU_nx551)) ;
    aoi22 L1_2_L2_3_G2_MINI_ALU_ix548 (.Y (L1_2_L2_3_G2_MINI_ALU_nx547), .A0 (
          L1Results_0__3), .A1 (L1Results_1__3), .B0 (L1_2_L2_3_G2_MINI_ALU_nx44
          ), .B1 (L1_2_L2_3_G2_MINI_ALU_nx18)) ;
    xnor2 L1_2_L2_3_G2_MINI_ALU_ix552 (.Y (L1_2_L2_3_G2_MINI_ALU_nx551), .A0 (
          L1Results_1__4), .A1 (L1Results_0__4)) ;
    xor2 L1_2_L2_3_G2_MINI_ALU_ix69 (.Y (L2Results_0__5), .A0 (
         L1_2_L2_3_G2_MINI_ALU_nx554), .A1 (L1_2_L2_3_G2_MINI_ALU_nx558)) ;
    aoi22 L1_2_L2_3_G2_MINI_ALU_ix555 (.Y (L1_2_L2_3_G2_MINI_ALU_nx554), .A0 (
          L1Results_0__4), .A1 (L1Results_1__4), .B0 (L1_2_L2_3_G2_MINI_ALU_nx48
          ), .B1 (L1_2_L2_3_G2_MINI_ALU_nx12)) ;
    xnor2 L1_2_L2_3_G2_MINI_ALU_ix559 (.Y (L1_2_L2_3_G2_MINI_ALU_nx558), .A0 (
          L1Results_1__5), .A1 (L1Results_0__5)) ;
    xor2 L1_2_L2_3_G2_MINI_ALU_ix67 (.Y (L2Results_0__6), .A0 (
         L1_2_L2_3_G2_MINI_ALU_nx561), .A1 (L1_2_L2_3_G2_MINI_ALU_nx565)) ;
    aoi22 L1_2_L2_3_G2_MINI_ALU_ix562 (.Y (L1_2_L2_3_G2_MINI_ALU_nx561), .A0 (
          L1Results_0__5), .A1 (L1Results_1__5), .B0 (L1_2_L2_3_G2_MINI_ALU_nx52
          ), .B1 (L1_2_L2_3_G2_MINI_ALU_nx6)) ;
    xnor2 L1_2_L2_3_G2_MINI_ALU_ix566 (.Y (L1_2_L2_3_G2_MINI_ALU_nx565), .A0 (
          L1Results_1__6), .A1 (L1Results_0__6)) ;
    xnor2 L1_2_L2_3_G2_MINI_ALU_ix65 (.Y (L2Results_0__7), .A0 (
          L1_2_L2_3_G2_MINI_ALU_nx568), .A1 (L1_2_L2_3_G2_MINI_ALU_nx62)) ;
    aoi22 L1_2_L2_3_G2_MINI_ALU_ix569 (.Y (L1_2_L2_3_G2_MINI_ALU_nx568), .A0 (
          L1Results_0__6), .A1 (L1Results_1__6), .B0 (L1_2_L2_3_G2_MINI_ALU_nx56
          ), .B1 (L1_2_L2_3_G2_MINI_ALU_nx0)) ;
    xor2 L1_2_L2_3_G2_MINI_ALU_ix63 (.Y (L1_2_L2_3_G2_MINI_ALU_nx62), .A0 (
         L1Results_1__7), .A1 (L1Results_0__7)) ;
    inv01 L1_2_L2_3_G2_MINI_ALU_ix155 (.Y (L1_2_L2_3_G2_MINI_ALU_nx154), .A (
          L1_2_L2_3_G2_MINI_ALU_nx383)) ;
    inv01 L1_2_L2_3_G2_MINI_ALU_ix57 (.Y (L1_2_L2_3_G2_MINI_ALU_nx56), .A (
          L1_2_L2_3_G2_MINI_ALU_nx561)) ;
    inv01 L1_2_L2_3_G2_MINI_ALU_ix53 (.Y (L1_2_L2_3_G2_MINI_ALU_nx52), .A (
          L1_2_L2_3_G2_MINI_ALU_nx554)) ;
    inv01 L1_2_L2_3_G2_MINI_ALU_ix49 (.Y (L1_2_L2_3_G2_MINI_ALU_nx48), .A (
          L1_2_L2_3_G2_MINI_ALU_nx547)) ;
    inv01 L1_2_L2_3_G2_MINI_ALU_ix45 (.Y (L1_2_L2_3_G2_MINI_ALU_nx44), .A (
          L1_2_L2_3_G2_MINI_ALU_nx540)) ;
    inv01 L1_2_L2_3_G2_MINI_ALU_ix41 (.Y (L1_2_L2_3_G2_MINI_ALU_nx40), .A (
          L1_2_L2_3_G2_MINI_ALU_nx534)) ;
    inv01 L1_2_L2_3_G2_MINI_ALU_ix31 (.Y (L1_2_L2_3_G2_MINI_ALU_nx30), .A (
          L1_2_L2_3_G2_MINI_ALU_nx531)) ;
    inv01 L1_2_L2_3_G2_MINI_ALU_ix25 (.Y (L1_2_L2_3_G2_MINI_ALU_nx24), .A (
          L1_2_L2_3_G2_MINI_ALU_nx537)) ;
    inv01 L1_2_L2_3_G2_MINI_ALU_ix19 (.Y (L1_2_L2_3_G2_MINI_ALU_nx18), .A (
          L1_2_L2_3_G2_MINI_ALU_nx544)) ;
    inv01 L1_2_L2_3_G2_MINI_ALU_ix13 (.Y (L1_2_L2_3_G2_MINI_ALU_nx12), .A (
          L1_2_L2_3_G2_MINI_ALU_nx551)) ;
    inv01 L1_2_L2_3_G2_MINI_ALU_ix7 (.Y (L1_2_L2_3_G2_MINI_ALU_nx6), .A (
          L1_2_L2_3_G2_MINI_ALU_nx558)) ;
    inv01 L1_2_L2_3_G2_MINI_ALU_ix1 (.Y (L1_2_L2_3_G2_MINI_ALU_nx0), .A (
          L1_2_L2_3_G2_MINI_ALU_nx565)) ;
    fake_gnd L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix216 (.Y (
             L1_2_L2_3_G2_MINI_ALU_WindowCellShiftedLeft_16)) ;
    nor02ii L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix81 (.Y (
            L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx80), .A0 (Instr), .A1 (Start)) ;
    aoi21 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix77 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_10), .A0 (
          FilterDin_2__3__1), .A1 (FilterDin_2__3__0), .B0 (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx4)) ;
    nor02_2x L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix5 (.Y (
             L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx4), .A0 (FilterDin_2__3__0), .A1 (
             FilterDin_2__3__1)) ;
    aoi21 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix67 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_11), .A0 (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx328), .A1 (FilterDin_2__3__2), .B0 (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx8)) ;
    nor03_2x L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix9 (.Y (
             L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx8), .A0 (FilterDin_2__3__2), .A1 (
             FilterDin_2__3__0), .A2 (FilterDin_2__3__1)) ;
    xnor2 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix59 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_12), .A0 (
          FilterDin_2__3__3), .A1 (L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx8)) ;
    xnor2 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix51 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_13), .A0 (
          FilterDin_2__3__4), .A1 (L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx12)) ;
    nor04 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix13 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx12), .A0 (FilterDin_2__3__3), .A1 (
          FilterDin_2__3__2), .A2 (FilterDin_2__3__0), .A3 (FilterDin_2__3__1)
          ) ;
    xnor2 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix43 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_14), .A0 (
          FilterDin_2__3__5), .A1 (L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx16)) ;
    nor02ii L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix17 (.Y (
            L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx16), .A0 (FilterDin_2__3__4), .A1 (
            L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx12)) ;
    xnor2 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix35 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_15), .A0 (
          FilterDin_2__3__6), .A1 (L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx20)) ;
    nor02ii L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix21 (.Y (
            L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx20), .A0 (FilterDin_2__3__5), .A1 (
            L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx16)) ;
    xnor2 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix27 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_16), .A0 (
          FilterDin_2__3__7), .A1 (L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx24)) ;
    nor02ii L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix25 (.Y (
            L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx24), .A0 (FilterDin_2__3__6), .A1 (
            L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx20)) ;
    inv01 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix329 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx328), .A (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx4)) ;
    inv02 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix383 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx384), .A (
          L1_2_L2_3_G2_MINI_ALU_BoothP_0)) ;
    dff L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_0 (.Q (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_0), .QB (\$dummy [667]), 
        .D (L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .CLK (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    nor02_2x L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix567 (.Y (
             L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566), .A0 (RST), .A1 (
             L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644)) ;
    dff L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_1 (.Q (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_1), .QB (\$dummy [668]), 
        .D (L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .CLK (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_2 (.Q (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_2), .QB (\$dummy [669]), 
        .D (L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .CLK (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_3 (.Q (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_3), .QB (\$dummy [670]), 
        .D (L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .CLK (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_4 (.Q (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_4), .QB (\$dummy [671]), 
        .D (L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .CLK (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_5 (.Q (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_5), .QB (\$dummy [672]), 
        .D (L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .CLK (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_6 (.Q (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_6), .QB (\$dummy [673]), 
        .D (L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .CLK (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_7 (.Q (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_7), .QB (\$dummy [674]), 
        .D (L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .CLK (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_8 (.Q (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_8), .QB (\$dummy [675]), 
        .D (L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .CLK (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_9 (.Q (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_9), .QB (\$dummy [676]), 
        .D (L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .CLK (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_10 (.Q (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_10), .QB (\$dummy [677])
        , .D (L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .CLK (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_11 (.Q (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_11), .QB (\$dummy [678])
        , .D (L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .CLK (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_12 (.Q (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_12), .QB (\$dummy [679])
        , .D (L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .CLK (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_13 (.Q (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_13), .QB (\$dummy [680])
        , .D (L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .CLK (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_14 (.Q (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_14), .QB (\$dummy [681])
        , .D (L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .CLK (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_15 (.Q (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_15), .QB (\$dummy [682])
        , .D (L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .CLK (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_16 (.Q (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_16), .QB (\$dummy [683])
        , .D (L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .CLK (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    inv02 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix623 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624), .A (CLK)) ;
    inv02 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix625 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626), .A (CLK)) ;
    inv02 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix627 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628), .A (CLK)) ;
    inv02 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix643 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644), .A (nx8138)) ;
    dff L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_0 (.Q (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_0), .QB (\$dummy [684]), 
        .D (L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .CLK (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    nor02_2x L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix567 (.Y (
             L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566), .A0 (RST), .A1 (
             L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644)) ;
    dff L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_1 (.Q (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_1), .QB (\$dummy [685]), 
        .D (L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .CLK (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_2 (.Q (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_2), .QB (\$dummy [686]), 
        .D (L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .CLK (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_3 (.Q (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_3), .QB (\$dummy [687]), 
        .D (L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .CLK (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_4 (.Q (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_4), .QB (\$dummy [688]), 
        .D (L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .CLK (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_5 (.Q (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_5), .QB (\$dummy [689]), 
        .D (L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .CLK (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_6 (.Q (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_6), .QB (\$dummy [690]), 
        .D (L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .CLK (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_7 (.Q (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_7), .QB (\$dummy [691]), 
        .D (L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .CLK (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_8 (.Q (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_8), .QB (\$dummy [692]), 
        .D (L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .CLK (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_9 (.Q (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_9), .QB (\$dummy [693]), 
        .D (L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .CLK (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_10 (.Q (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_10), .QB (\$dummy [694])
        , .D (L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .CLK (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_11 (.Q (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_11), .QB (\$dummy [695])
        , .D (L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .CLK (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_12 (.Q (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_12), .QB (\$dummy [696])
        , .D (L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .CLK (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_13 (.Q (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_13), .QB (\$dummy [697])
        , .D (L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .CLK (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_14 (.Q (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_14), .QB (\$dummy [698])
        , .D (L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .CLK (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_15 (.Q (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_15), .QB (\$dummy [699])
        , .D (L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .CLK (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_16 (.Q (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_16), .QB (\$dummy [700])
        , .D (L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .CLK (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    inv02 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix623 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624), .A (CLK)) ;
    inv02 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix625 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626), .A (CLK)) ;
    inv02 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix627 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628), .A (CLK)) ;
    inv02 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix643 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644), .A (nx8144)) ;
    dff L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_0 (.Q (
        L1_2_L2_3_G2_MINI_ALU_BoothP_0), .QB (\$dummy [701]), .D (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .CLK (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    nor02_2x L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix567 (.Y (
             L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566), .A0 (RST), .A1 (
             L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    dff L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_1 (.Q (
        L1_2_L2_3_G2_MINI_ALU_BoothP_1), .QB (\$dummy [702]), .D (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .CLK (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_2 (.Q (
        L1_2_L2_3_G2_MINI_ALU_BoothP_2), .QB (\$dummy [703]), .D (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .CLK (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_3 (.Q (
        L1_2_L2_3_G2_MINI_ALU_BoothP_3), .QB (\$dummy [704]), .D (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .CLK (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_4 (.Q (
        L1_2_L2_3_G2_MINI_ALU_BoothP_4), .QB (\$dummy [705]), .D (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .CLK (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_5 (.Q (
        L1_2_L2_3_G2_MINI_ALU_BoothP_5), .QB (\$dummy [706]), .D (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .CLK (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_6 (.Q (
        L1_2_L2_3_G2_MINI_ALU_BoothP_6), .QB (\$dummy [707]), .D (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .CLK (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_7 (.Q (
        L1_2_L2_3_G2_MINI_ALU_BoothP_7), .QB (\$dummy [708]), .D (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .CLK (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_8 (.Q (
        L1_2_L2_3_G2_MINI_ALU_BoothP_8), .QB (\$dummy [709]), .D (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .CLK (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_9 (.Q (
        L1_2_L2_3_G2_MINI_ALU_BoothP_9), .QB (\$dummy [710]), .D (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .CLK (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_10 (.Q (
        L1_2_L2_3_G2_MINI_ALU_BoothP_10), .QB (\$dummy [711]), .D (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .CLK (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_11 (.Q (
        L1_2_L2_3_G2_MINI_ALU_BoothP_11), .QB (\$dummy [712]), .D (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .CLK (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_12 (.Q (
        L1_2_L2_3_G2_MINI_ALU_BoothP_12), .QB (\$dummy [713]), .D (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .CLK (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_13 (.Q (
        L1_2_L2_3_G2_MINI_ALU_BoothP_13), .QB (\$dummy [714]), .D (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .CLK (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_14 (.Q (
        L1_2_L2_3_G2_MINI_ALU_BoothP_14), .QB (\$dummy [715]), .D (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .CLK (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_15 (.Q (
        L1_2_L2_3_G2_MINI_ALU_BoothP_15), .QB (\$dummy [716]), .D (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .CLK (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_16 (.Q (
        L1_2_L2_3_G2_MINI_ALU_BoothP_16), .QB (\$dummy [717]), .D (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .CLK (
        L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    inv02 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix623 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624), .A (CLK)) ;
    inv02 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix625 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626), .A (CLK)) ;
    inv02 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix627 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628), .A (CLK)) ;
    inv02 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix643 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644), .A (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642)) ;
    xor2 L1_2_L2_4_G2_MINI_ALU_ix83 (.Y (L2Results_1__0), .A0 (L1Results_3__0), 
         .A1 (L1Results_2__0)) ;
    xnor2 L1_2_L2_4_G2_MINI_ALU_ix380 (.Y (L1_2_L2_4_G2_MINI_ALU_nx379), .A0 (
          L1_2_L2_4_G2_MINI_ALU_nx381), .A1 (L1_2_L2_4_G2_MINI_ALU_nx383)) ;
    nand02 L1_2_L2_4_G2_MINI_ALU_ix382 (.Y (L1_2_L2_4_G2_MINI_ALU_nx381), .A0 (
           L1_2_L2_4_G2_MINI_ALU_BoothOperand_0), .A1 (nx8164)) ;
    xnor2 L1_2_L2_4_G2_MINI_ALU_ix384 (.Y (L1_2_L2_4_G2_MINI_ALU_nx383), .A0 (
          L1_2_L2_4_G2_MINI_ALU_BoothOperand_1), .A1 (
          L1_2_L2_4_G2_MINI_ALU_BoothP_1)) ;
    inv01 L1_2_L2_4_G2_MINI_ALU_ix388 (.Y (L1_2_L2_4_G2_MINI_ALU_nx387), .A (
          L1_2_L2_4_G2_MINI_ALU_BoothP_2)) ;
    xnor2 L1_2_L2_4_G2_MINI_ALU_ix390 (.Y (L1_2_L2_4_G2_MINI_ALU_nx389), .A0 (
          L1_2_L2_4_G2_MINI_ALU_nx391), .A1 (L1_2_L2_4_G2_MINI_ALU_nx395)) ;
    aoi32 L1_2_L2_4_G2_MINI_ALU_ix392 (.Y (L1_2_L2_4_G2_MINI_ALU_nx391), .A0 (
          L1_2_L2_4_G2_MINI_ALU_BoothOperand_0), .A1 (nx8164), .A2 (
          L1_2_L2_4_G2_MINI_ALU_nx154), .B0 (L1_2_L2_4_G2_MINI_ALU_BoothP_1), .B1 (
          L1_2_L2_4_G2_MINI_ALU_BoothOperand_1)) ;
    xnor2 L1_2_L2_4_G2_MINI_ALU_ix396 (.Y (L1_2_L2_4_G2_MINI_ALU_nx395), .A0 (
          L1_2_L2_4_G2_MINI_ALU_BoothOperand_2), .A1 (
          L1_2_L2_4_G2_MINI_ALU_BoothP_2)) ;
    inv01 L1_2_L2_4_G2_MINI_ALU_ix400 (.Y (L1_2_L2_4_G2_MINI_ALU_nx399), .A (
          L1_2_L2_4_G2_MINI_ALU_BoothP_3)) ;
    xnor2 L1_2_L2_4_G2_MINI_ALU_ix402 (.Y (L1_2_L2_4_G2_MINI_ALU_nx401), .A0 (
          L1_2_L2_4_G2_MINI_ALU_nx403), .A1 (L1_2_L2_4_G2_MINI_ALU_nx405)) ;
    xnor2 L1_2_L2_4_G2_MINI_ALU_ix406 (.Y (L1_2_L2_4_G2_MINI_ALU_nx405), .A0 (
          L1_2_L2_4_G2_MINI_ALU_BoothOperand_3), .A1 (
          L1_2_L2_4_G2_MINI_ALU_BoothP_3)) ;
    inv01 L1_2_L2_4_G2_MINI_ALU_ix410 (.Y (L1_2_L2_4_G2_MINI_ALU_nx409), .A (
          L1_2_L2_4_G2_MINI_ALU_BoothP_4)) ;
    xnor2 L1_2_L2_4_G2_MINI_ALU_ix412 (.Y (L1_2_L2_4_G2_MINI_ALU_nx411), .A0 (
          L1_2_L2_4_G2_MINI_ALU_nx413), .A1 (L1_2_L2_4_G2_MINI_ALU_nx415)) ;
    xnor2 L1_2_L2_4_G2_MINI_ALU_ix416 (.Y (L1_2_L2_4_G2_MINI_ALU_nx415), .A0 (
          L1_2_L2_4_G2_MINI_ALU_BoothOperand_4), .A1 (
          L1_2_L2_4_G2_MINI_ALU_BoothP_4)) ;
    inv01 L1_2_L2_4_G2_MINI_ALU_ix420 (.Y (L1_2_L2_4_G2_MINI_ALU_nx419), .A (
          L1_2_L2_4_G2_MINI_ALU_BoothP_5)) ;
    xnor2 L1_2_L2_4_G2_MINI_ALU_ix422 (.Y (L1_2_L2_4_G2_MINI_ALU_nx421), .A0 (
          L1_2_L2_4_G2_MINI_ALU_nx423), .A1 (L1_2_L2_4_G2_MINI_ALU_nx425)) ;
    xnor2 L1_2_L2_4_G2_MINI_ALU_ix426 (.Y (L1_2_L2_4_G2_MINI_ALU_nx425), .A0 (
          L1_2_L2_4_G2_MINI_ALU_BoothOperand_5), .A1 (
          L1_2_L2_4_G2_MINI_ALU_BoothP_5)) ;
    inv01 L1_2_L2_4_G2_MINI_ALU_ix430 (.Y (L1_2_L2_4_G2_MINI_ALU_nx429), .A (
          L1_2_L2_4_G2_MINI_ALU_BoothP_6)) ;
    xnor2 L1_2_L2_4_G2_MINI_ALU_ix432 (.Y (L1_2_L2_4_G2_MINI_ALU_nx431), .A0 (
          L1_2_L2_4_G2_MINI_ALU_nx433), .A1 (L1_2_L2_4_G2_MINI_ALU_nx435)) ;
    xnor2 L1_2_L2_4_G2_MINI_ALU_ix436 (.Y (L1_2_L2_4_G2_MINI_ALU_nx435), .A0 (
          L1_2_L2_4_G2_MINI_ALU_BoothOperand_6), .A1 (
          L1_2_L2_4_G2_MINI_ALU_BoothP_6)) ;
    inv01 L1_2_L2_4_G2_MINI_ALU_ix440 (.Y (L1_2_L2_4_G2_MINI_ALU_nx439), .A (
          L1_2_L2_4_G2_MINI_ALU_BoothP_7)) ;
    xnor2 L1_2_L2_4_G2_MINI_ALU_ix442 (.Y (L1_2_L2_4_G2_MINI_ALU_nx441), .A0 (
          L1_2_L2_4_G2_MINI_ALU_nx443), .A1 (L1_2_L2_4_G2_MINI_ALU_nx445)) ;
    xnor2 L1_2_L2_4_G2_MINI_ALU_ix446 (.Y (L1_2_L2_4_G2_MINI_ALU_nx445), .A0 (
          L1_2_L2_4_G2_MINI_ALU_BoothOperand_7), .A1 (
          L1_2_L2_4_G2_MINI_ALU_BoothP_7)) ;
    inv01 L1_2_L2_4_G2_MINI_ALU_ix450 (.Y (L1_2_L2_4_G2_MINI_ALU_nx449), .A (
          L1_2_L2_4_G2_MINI_ALU_BoothP_8)) ;
    xnor2 L1_2_L2_4_G2_MINI_ALU_ix452 (.Y (L1_2_L2_4_G2_MINI_ALU_nx451), .A0 (
          L1_2_L2_4_G2_MINI_ALU_nx453), .A1 (L1_2_L2_4_G2_MINI_ALU_nx455)) ;
    xnor2 L1_2_L2_4_G2_MINI_ALU_ix456 (.Y (L1_2_L2_4_G2_MINI_ALU_nx455), .A0 (
          L1_2_L2_4_G2_MINI_ALU_BoothOperand_8), .A1 (
          L1_2_L2_4_G2_MINI_ALU_BoothP_8)) ;
    xor2 L1_2_L2_4_G2_MINI_ALU_ix317 (.Y (L1_2_L2_4_G2_MINI_ALU_nx316), .A0 (
         L1_2_L2_4_G2_MINI_ALU_nx461), .A1 (L1_2_L2_4_G2_MINI_ALU_nx463)) ;
    xnor2 L1_2_L2_4_G2_MINI_ALU_ix464 (.Y (L1_2_L2_4_G2_MINI_ALU_nx463), .A0 (
          L1_2_L2_4_G2_MINI_ALU_BoothOperand_9), .A1 (
          L1_2_L2_4_G2_MINI_ALU_BoothP_9)) ;
    xor2 L1_2_L2_4_G2_MINI_ALU_ix337 (.Y (L1_2_L2_4_G2_MINI_ALU_nx336), .A0 (
         L1_2_L2_4_G2_MINI_ALU_nx467), .A1 (L1_2_L2_4_G2_MINI_ALU_nx471)) ;
    inv01 L1_2_L2_4_G2_MINI_ALU_ix470 (.Y (L1_2_L2_4_G2_MINI_ALU_nx469), .A (
          L1_2_L2_4_G2_MINI_ALU_BoothP_9)) ;
    xnor2 L1_2_L2_4_G2_MINI_ALU_ix472 (.Y (L1_2_L2_4_G2_MINI_ALU_nx471), .A0 (
          L1_2_L2_4_G2_MINI_ALU_BoothOperand_10), .A1 (
          L1_2_L2_4_G2_MINI_ALU_BoothP_10)) ;
    xor2 L1_2_L2_4_G2_MINI_ALU_ix357 (.Y (L1_2_L2_4_G2_MINI_ALU_nx356), .A0 (
         L1_2_L2_4_G2_MINI_ALU_nx475), .A1 (L1_2_L2_4_G2_MINI_ALU_nx479)) ;
    inv01 L1_2_L2_4_G2_MINI_ALU_ix478 (.Y (L1_2_L2_4_G2_MINI_ALU_nx477), .A (
          L1_2_L2_4_G2_MINI_ALU_BoothP_10)) ;
    xnor2 L1_2_L2_4_G2_MINI_ALU_ix480 (.Y (L1_2_L2_4_G2_MINI_ALU_nx479), .A0 (
          L1_2_L2_4_G2_MINI_ALU_BoothOperand_11), .A1 (
          L1_2_L2_4_G2_MINI_ALU_BoothP_11)) ;
    xor2 L1_2_L2_4_G2_MINI_ALU_ix377 (.Y (L1_2_L2_4_G2_MINI_ALU_nx376), .A0 (
         L1_2_L2_4_G2_MINI_ALU_nx483), .A1 (L1_2_L2_4_G2_MINI_ALU_nx487)) ;
    inv01 L1_2_L2_4_G2_MINI_ALU_ix486 (.Y (L1_2_L2_4_G2_MINI_ALU_nx485), .A (
          L1_2_L2_4_G2_MINI_ALU_BoothP_11)) ;
    xnor2 L1_2_L2_4_G2_MINI_ALU_ix488 (.Y (L1_2_L2_4_G2_MINI_ALU_nx487), .A0 (
          L1_2_L2_4_G2_MINI_ALU_BoothOperand_12), .A1 (
          L1_2_L2_4_G2_MINI_ALU_BoothP_12)) ;
    xor2 L1_2_L2_4_G2_MINI_ALU_ix397 (.Y (L1_2_L2_4_G2_MINI_ALU_nx396), .A0 (
         L1_2_L2_4_G2_MINI_ALU_nx491), .A1 (L1_2_L2_4_G2_MINI_ALU_nx495)) ;
    inv01 L1_2_L2_4_G2_MINI_ALU_ix494 (.Y (L1_2_L2_4_G2_MINI_ALU_nx493), .A (
          L1_2_L2_4_G2_MINI_ALU_BoothP_12)) ;
    xnor2 L1_2_L2_4_G2_MINI_ALU_ix496 (.Y (L1_2_L2_4_G2_MINI_ALU_nx495), .A0 (
          L1_2_L2_4_G2_MINI_ALU_BoothOperand_13), .A1 (
          L1_2_L2_4_G2_MINI_ALU_BoothP_13)) ;
    xor2 L1_2_L2_4_G2_MINI_ALU_ix417 (.Y (L1_2_L2_4_G2_MINI_ALU_nx416), .A0 (
         L1_2_L2_4_G2_MINI_ALU_nx499), .A1 (L1_2_L2_4_G2_MINI_ALU_nx503)) ;
    inv01 L1_2_L2_4_G2_MINI_ALU_ix502 (.Y (L1_2_L2_4_G2_MINI_ALU_nx501), .A (
          L1_2_L2_4_G2_MINI_ALU_BoothP_13)) ;
    xnor2 L1_2_L2_4_G2_MINI_ALU_ix504 (.Y (L1_2_L2_4_G2_MINI_ALU_nx503), .A0 (
          L1_2_L2_4_G2_MINI_ALU_BoothOperand_14), .A1 (
          L1_2_L2_4_G2_MINI_ALU_BoothP_14)) ;
    xor2 L1_2_L2_4_G2_MINI_ALU_ix437 (.Y (L1_2_L2_4_G2_MINI_ALU_nx436), .A0 (
         L1_2_L2_4_G2_MINI_ALU_nx507), .A1 (L1_2_L2_4_G2_MINI_ALU_nx511)) ;
    inv01 L1_2_L2_4_G2_MINI_ALU_ix510 (.Y (L1_2_L2_4_G2_MINI_ALU_nx509), .A (
          L1_2_L2_4_G2_MINI_ALU_BoothP_14)) ;
    xnor2 L1_2_L2_4_G2_MINI_ALU_ix512 (.Y (L1_2_L2_4_G2_MINI_ALU_nx511), .A0 (
          L1_2_L2_4_G2_MINI_ALU_BoothOperand_15), .A1 (
          L1_2_L2_4_G2_MINI_ALU_BoothP_15)) ;
    xnor2 L1_2_L2_4_G2_MINI_ALU_ix457 (.Y (L1_2_L2_4_G2_MINI_ALU_nx456), .A0 (
          L1_2_L2_4_G2_MINI_ALU_nx515), .A1 (L1_2_L2_4_G2_MINI_ALU_nx454)) ;
    inv01 L1_2_L2_4_G2_MINI_ALU_ix518 (.Y (L1_2_L2_4_G2_MINI_ALU_nx517), .A (
          L1_2_L2_4_G2_MINI_ALU_BoothP_15)) ;
    xor2 L1_2_L2_4_G2_MINI_ALU_ix455 (.Y (L1_2_L2_4_G2_MINI_ALU_nx454), .A0 (
         L1_2_L2_4_G2_MINI_ALU_BoothOperand_16), .A1 (
         L1_2_L2_4_G2_MINI_ALU_BoothP_16)) ;
    mux21_ni L1_2_L2_4_G2_MINI_ALU_ix91 (.Y (L1FirstOperands_2__0), .A0 (
             L1_2_L2_4_G2_MINI_ALU_BoothP_1), .A1 (WindowDin_2__4__0), .S0 (
             Instr)) ;
    mux21_ni L1_2_L2_4_G2_MINI_ALU_ix99 (.Y (L1FirstOperands_2__1), .A0 (
             L1_2_L2_4_G2_MINI_ALU_BoothP_2), .A1 (WindowDin_2__4__1), .S0 (
             Instr)) ;
    mux21_ni L1_2_L2_4_G2_MINI_ALU_ix107 (.Y (L1FirstOperands_2__2), .A0 (
             L1_2_L2_4_G2_MINI_ALU_BoothP_3), .A1 (WindowDin_2__4__2), .S0 (
             Instr)) ;
    mux21_ni L1_2_L2_4_G2_MINI_ALU_ix115 (.Y (L1FirstOperands_2__3), .A0 (
             L1_2_L2_4_G2_MINI_ALU_BoothP_4), .A1 (WindowDin_2__4__3), .S0 (
             Instr)) ;
    mux21_ni L1_2_L2_4_G2_MINI_ALU_ix123 (.Y (L1FirstOperands_2__4), .A0 (
             L1_2_L2_4_G2_MINI_ALU_BoothP_5), .A1 (WindowDin_2__4__4), .S0 (
             Instr)) ;
    mux21_ni L1_2_L2_4_G2_MINI_ALU_ix131 (.Y (L1FirstOperands_2__5), .A0 (
             L1_2_L2_4_G2_MINI_ALU_BoothP_6), .A1 (WindowDin_2__4__5), .S0 (
             Instr)) ;
    mux21_ni L1_2_L2_4_G2_MINI_ALU_ix139 (.Y (L1FirstOperands_2__6), .A0 (
             L1_2_L2_4_G2_MINI_ALU_BoothP_7), .A1 (WindowDin_2__4__6), .S0 (
             Instr)) ;
    mux21_ni L1_2_L2_4_G2_MINI_ALU_ix147 (.Y (L1FirstOperands_2__7), .A0 (
             L1_2_L2_4_G2_MINI_ALU_BoothP_8), .A1 (WindowDin_2__4__7), .S0 (
             Instr)) ;
    xor2 L1_2_L2_4_G2_MINI_ALU_ix77 (.Y (L2Results_1__1), .A0 (
         L1_2_L2_4_G2_MINI_ALU_nx529), .A1 (L1_2_L2_4_G2_MINI_ALU_nx531)) ;
    nand02 L1_2_L2_4_G2_MINI_ALU_ix530 (.Y (L1_2_L2_4_G2_MINI_ALU_nx529), .A0 (
           L1Results_3__0), .A1 (L1Results_2__0)) ;
    xnor2 L1_2_L2_4_G2_MINI_ALU_ix532 (.Y (L1_2_L2_4_G2_MINI_ALU_nx531), .A0 (
          L1Results_3__1), .A1 (L1Results_2__1)) ;
    xor2 L1_2_L2_4_G2_MINI_ALU_ix75 (.Y (L2Results_1__2), .A0 (
         L1_2_L2_4_G2_MINI_ALU_nx534), .A1 (L1_2_L2_4_G2_MINI_ALU_nx537)) ;
    aoi32 L1_2_L2_4_G2_MINI_ALU_ix535 (.Y (L1_2_L2_4_G2_MINI_ALU_nx534), .A0 (
          L1Results_3__0), .A1 (L1Results_2__0), .A2 (L1_2_L2_4_G2_MINI_ALU_nx30
          ), .B0 (L1Results_2__1), .B1 (L1Results_3__1)) ;
    xnor2 L1_2_L2_4_G2_MINI_ALU_ix538 (.Y (L1_2_L2_4_G2_MINI_ALU_nx537), .A0 (
          L1Results_3__2), .A1 (L1Results_2__2)) ;
    xor2 L1_2_L2_4_G2_MINI_ALU_ix73 (.Y (L2Results_1__3), .A0 (
         L1_2_L2_4_G2_MINI_ALU_nx540), .A1 (L1_2_L2_4_G2_MINI_ALU_nx544)) ;
    aoi22 L1_2_L2_4_G2_MINI_ALU_ix541 (.Y (L1_2_L2_4_G2_MINI_ALU_nx540), .A0 (
          L1Results_2__2), .A1 (L1Results_3__2), .B0 (L1_2_L2_4_G2_MINI_ALU_nx40
          ), .B1 (L1_2_L2_4_G2_MINI_ALU_nx24)) ;
    xnor2 L1_2_L2_4_G2_MINI_ALU_ix545 (.Y (L1_2_L2_4_G2_MINI_ALU_nx544), .A0 (
          L1Results_3__3), .A1 (L1Results_2__3)) ;
    xor2 L1_2_L2_4_G2_MINI_ALU_ix71 (.Y (L2Results_1__4), .A0 (
         L1_2_L2_4_G2_MINI_ALU_nx547), .A1 (L1_2_L2_4_G2_MINI_ALU_nx551)) ;
    aoi22 L1_2_L2_4_G2_MINI_ALU_ix548 (.Y (L1_2_L2_4_G2_MINI_ALU_nx547), .A0 (
          L1Results_2__3), .A1 (L1Results_3__3), .B0 (L1_2_L2_4_G2_MINI_ALU_nx44
          ), .B1 (L1_2_L2_4_G2_MINI_ALU_nx18)) ;
    xnor2 L1_2_L2_4_G2_MINI_ALU_ix552 (.Y (L1_2_L2_4_G2_MINI_ALU_nx551), .A0 (
          L1Results_3__4), .A1 (L1Results_2__4)) ;
    xor2 L1_2_L2_4_G2_MINI_ALU_ix69 (.Y (L2Results_1__5), .A0 (
         L1_2_L2_4_G2_MINI_ALU_nx554), .A1 (L1_2_L2_4_G2_MINI_ALU_nx558)) ;
    aoi22 L1_2_L2_4_G2_MINI_ALU_ix555 (.Y (L1_2_L2_4_G2_MINI_ALU_nx554), .A0 (
          L1Results_2__4), .A1 (L1Results_3__4), .B0 (L1_2_L2_4_G2_MINI_ALU_nx48
          ), .B1 (L1_2_L2_4_G2_MINI_ALU_nx12)) ;
    xnor2 L1_2_L2_4_G2_MINI_ALU_ix559 (.Y (L1_2_L2_4_G2_MINI_ALU_nx558), .A0 (
          L1Results_3__5), .A1 (L1Results_2__5)) ;
    xor2 L1_2_L2_4_G2_MINI_ALU_ix67 (.Y (L2Results_1__6), .A0 (
         L1_2_L2_4_G2_MINI_ALU_nx561), .A1 (L1_2_L2_4_G2_MINI_ALU_nx565)) ;
    aoi22 L1_2_L2_4_G2_MINI_ALU_ix562 (.Y (L1_2_L2_4_G2_MINI_ALU_nx561), .A0 (
          L1Results_2__5), .A1 (L1Results_3__5), .B0 (L1_2_L2_4_G2_MINI_ALU_nx52
          ), .B1 (L1_2_L2_4_G2_MINI_ALU_nx6)) ;
    xnor2 L1_2_L2_4_G2_MINI_ALU_ix566 (.Y (L1_2_L2_4_G2_MINI_ALU_nx565), .A0 (
          L1Results_3__6), .A1 (L1Results_2__6)) ;
    xnor2 L1_2_L2_4_G2_MINI_ALU_ix65 (.Y (L2Results_1__7), .A0 (
          L1_2_L2_4_G2_MINI_ALU_nx568), .A1 (L1_2_L2_4_G2_MINI_ALU_nx62)) ;
    aoi22 L1_2_L2_4_G2_MINI_ALU_ix569 (.Y (L1_2_L2_4_G2_MINI_ALU_nx568), .A0 (
          L1Results_2__6), .A1 (L1Results_3__6), .B0 (L1_2_L2_4_G2_MINI_ALU_nx56
          ), .B1 (L1_2_L2_4_G2_MINI_ALU_nx0)) ;
    xor2 L1_2_L2_4_G2_MINI_ALU_ix63 (.Y (L1_2_L2_4_G2_MINI_ALU_nx62), .A0 (
         L1Results_3__7), .A1 (L1Results_2__7)) ;
    inv01 L1_2_L2_4_G2_MINI_ALU_ix155 (.Y (L1_2_L2_4_G2_MINI_ALU_nx154), .A (
          L1_2_L2_4_G2_MINI_ALU_nx383)) ;
    inv01 L1_2_L2_4_G2_MINI_ALU_ix57 (.Y (L1_2_L2_4_G2_MINI_ALU_nx56), .A (
          L1_2_L2_4_G2_MINI_ALU_nx561)) ;
    inv01 L1_2_L2_4_G2_MINI_ALU_ix53 (.Y (L1_2_L2_4_G2_MINI_ALU_nx52), .A (
          L1_2_L2_4_G2_MINI_ALU_nx554)) ;
    inv01 L1_2_L2_4_G2_MINI_ALU_ix49 (.Y (L1_2_L2_4_G2_MINI_ALU_nx48), .A (
          L1_2_L2_4_G2_MINI_ALU_nx547)) ;
    inv01 L1_2_L2_4_G2_MINI_ALU_ix45 (.Y (L1_2_L2_4_G2_MINI_ALU_nx44), .A (
          L1_2_L2_4_G2_MINI_ALU_nx540)) ;
    inv01 L1_2_L2_4_G2_MINI_ALU_ix41 (.Y (L1_2_L2_4_G2_MINI_ALU_nx40), .A (
          L1_2_L2_4_G2_MINI_ALU_nx534)) ;
    inv01 L1_2_L2_4_G2_MINI_ALU_ix31 (.Y (L1_2_L2_4_G2_MINI_ALU_nx30), .A (
          L1_2_L2_4_G2_MINI_ALU_nx531)) ;
    inv01 L1_2_L2_4_G2_MINI_ALU_ix25 (.Y (L1_2_L2_4_G2_MINI_ALU_nx24), .A (
          L1_2_L2_4_G2_MINI_ALU_nx537)) ;
    inv01 L1_2_L2_4_G2_MINI_ALU_ix19 (.Y (L1_2_L2_4_G2_MINI_ALU_nx18), .A (
          L1_2_L2_4_G2_MINI_ALU_nx544)) ;
    inv01 L1_2_L2_4_G2_MINI_ALU_ix13 (.Y (L1_2_L2_4_G2_MINI_ALU_nx12), .A (
          L1_2_L2_4_G2_MINI_ALU_nx551)) ;
    inv01 L1_2_L2_4_G2_MINI_ALU_ix7 (.Y (L1_2_L2_4_G2_MINI_ALU_nx6), .A (
          L1_2_L2_4_G2_MINI_ALU_nx558)) ;
    inv01 L1_2_L2_4_G2_MINI_ALU_ix1 (.Y (L1_2_L2_4_G2_MINI_ALU_nx0), .A (
          L1_2_L2_4_G2_MINI_ALU_nx565)) ;
    fake_gnd L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix216 (.Y (
             L1_2_L2_4_G2_MINI_ALU_WindowCellShiftedLeft_16)) ;
    nor02ii L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix81 (.Y (
            L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_nx80), .A0 (Instr), .A1 (Start)) ;
    aoi21 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix77 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_10), .A0 (
          FilterDin_2__4__1), .A1 (FilterDin_2__4__0), .B0 (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_nx4)) ;
    nor02_2x L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix5 (.Y (
             L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_nx4), .A0 (FilterDin_2__4__0), .A1 (
             FilterDin_2__4__1)) ;
    aoi21 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix67 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_11), .A0 (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_nx328), .A1 (FilterDin_2__4__2), .B0 (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_nx8)) ;
    nor03_2x L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix9 (.Y (
             L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_nx8), .A0 (FilterDin_2__4__2), .A1 (
             FilterDin_2__4__0), .A2 (FilterDin_2__4__1)) ;
    xnor2 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix59 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_12), .A0 (
          FilterDin_2__4__3), .A1 (L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_nx8)) ;
    xnor2 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix51 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_13), .A0 (
          FilterDin_2__4__4), .A1 (L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_nx12)) ;
    nor04 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix13 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_nx12), .A0 (FilterDin_2__4__3), .A1 (
          FilterDin_2__4__2), .A2 (FilterDin_2__4__0), .A3 (FilterDin_2__4__1)
          ) ;
    xnor2 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix43 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_14), .A0 (
          FilterDin_2__4__5), .A1 (L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_nx16)) ;
    nor02ii L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix17 (.Y (
            L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_nx16), .A0 (FilterDin_2__4__4), .A1 (
            L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_nx12)) ;
    xnor2 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix35 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_15), .A0 (
          FilterDin_2__4__6), .A1 (L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_nx20)) ;
    nor02ii L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix21 (.Y (
            L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_nx20), .A0 (FilterDin_2__4__5), .A1 (
            L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_nx16)) ;
    xnor2 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix27 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_16), .A0 (
          FilterDin_2__4__7), .A1 (L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_nx24)) ;
    nor02ii L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix25 (.Y (
            L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_nx24), .A0 (FilterDin_2__4__6), .A1 (
            L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_nx20)) ;
    inv01 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix329 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_nx328), .A (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_nx4)) ;
    inv02 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix383 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_nx384), .A (
          L1_2_L2_4_G2_MINI_ALU_BoothP_0)) ;
    dff L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_0 (.Q (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_0), .QB (\$dummy [718]), 
        .D (L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .CLK (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    nor02_2x L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix567 (.Y (
             L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566), .A0 (RST), .A1 (
             L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644)) ;
    dff L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_1 (.Q (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_1), .QB (\$dummy [719]), 
        .D (L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .CLK (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_2 (.Q (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_2), .QB (\$dummy [720]), 
        .D (L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .CLK (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_3 (.Q (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_3), .QB (\$dummy [721]), 
        .D (L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .CLK (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_4 (.Q (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_4), .QB (\$dummy [722]), 
        .D (L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .CLK (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_5 (.Q (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_5), .QB (\$dummy [723]), 
        .D (L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .CLK (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_6 (.Q (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_6), .QB (\$dummy [724]), 
        .D (L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .CLK (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_7 (.Q (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_7), .QB (\$dummy [725]), 
        .D (L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .CLK (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_8 (.Q (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_8), .QB (\$dummy [726]), 
        .D (L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .CLK (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_9 (.Q (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_9), .QB (\$dummy [727]), 
        .D (L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .CLK (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_10 (.Q (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_10), .QB (\$dummy [728])
        , .D (L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .CLK (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_11 (.Q (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_11), .QB (\$dummy [729])
        , .D (L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .CLK (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_12 (.Q (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_12), .QB (\$dummy [730])
        , .D (L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .CLK (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_13 (.Q (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_13), .QB (\$dummy [731])
        , .D (L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .CLK (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_14 (.Q (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_14), .QB (\$dummy [732])
        , .D (L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .CLK (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_15 (.Q (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_15), .QB (\$dummy [733])
        , .D (L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .CLK (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_16 (.Q (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_16), .QB (\$dummy [734])
        , .D (L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .CLK (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    inv02 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix623 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624), .A (CLK)) ;
    inv02 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix625 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626), .A (CLK)) ;
    inv02 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix627 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628), .A (CLK)) ;
    inv02 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix643 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644), .A (nx8178)) ;
    dff L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_0 (.Q (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_0), .QB (\$dummy [735]), 
        .D (L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .CLK (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    nor02_2x L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix567 (.Y (
             L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566), .A0 (RST), .A1 (
             L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644)) ;
    dff L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_1 (.Q (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_1), .QB (\$dummy [736]), 
        .D (L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .CLK (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_2 (.Q (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_2), .QB (\$dummy [737]), 
        .D (L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .CLK (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_3 (.Q (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_3), .QB (\$dummy [738]), 
        .D (L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .CLK (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_4 (.Q (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_4), .QB (\$dummy [739]), 
        .D (L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .CLK (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_5 (.Q (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_5), .QB (\$dummy [740]), 
        .D (L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .CLK (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_6 (.Q (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_6), .QB (\$dummy [741]), 
        .D (L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .CLK (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_7 (.Q (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_7), .QB (\$dummy [742]), 
        .D (L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .CLK (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_8 (.Q (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_8), .QB (\$dummy [743]), 
        .D (L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .CLK (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_9 (.Q (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_9), .QB (\$dummy [744]), 
        .D (L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .CLK (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_10 (.Q (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_10), .QB (\$dummy [745])
        , .D (L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .CLK (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_11 (.Q (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_11), .QB (\$dummy [746])
        , .D (L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .CLK (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_12 (.Q (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_12), .QB (\$dummy [747])
        , .D (L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .CLK (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_13 (.Q (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_13), .QB (\$dummy [748])
        , .D (L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .CLK (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_14 (.Q (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_14), .QB (\$dummy [749])
        , .D (L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .CLK (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_15 (.Q (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_15), .QB (\$dummy [750])
        , .D (L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .CLK (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_16 (.Q (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_16), .QB (\$dummy [751])
        , .D (L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .CLK (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    inv02 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix623 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624), .A (CLK)) ;
    inv02 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix625 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626), .A (CLK)) ;
    inv02 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix627 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628), .A (CLK)) ;
    inv02 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix643 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644), .A (nx8184)) ;
    dff L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_0 (.Q (
        L1_2_L2_4_G2_MINI_ALU_BoothP_0), .QB (\$dummy [752]), .D (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .CLK (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    nor02_2x L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix567 (.Y (
             L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566), .A0 (RST), .A1 (
             L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    dff L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_1 (.Q (
        L1_2_L2_4_G2_MINI_ALU_BoothP_1), .QB (\$dummy [753]), .D (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .CLK (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_2 (.Q (
        L1_2_L2_4_G2_MINI_ALU_BoothP_2), .QB (\$dummy [754]), .D (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .CLK (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_3 (.Q (
        L1_2_L2_4_G2_MINI_ALU_BoothP_3), .QB (\$dummy [755]), .D (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .CLK (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_4 (.Q (
        L1_2_L2_4_G2_MINI_ALU_BoothP_4), .QB (\$dummy [756]), .D (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .CLK (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_5 (.Q (
        L1_2_L2_4_G2_MINI_ALU_BoothP_5), .QB (\$dummy [757]), .D (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .CLK (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_6 (.Q (
        L1_2_L2_4_G2_MINI_ALU_BoothP_6), .QB (\$dummy [758]), .D (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .CLK (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_7 (.Q (
        L1_2_L2_4_G2_MINI_ALU_BoothP_7), .QB (\$dummy [759]), .D (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .CLK (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_8 (.Q (
        L1_2_L2_4_G2_MINI_ALU_BoothP_8), .QB (\$dummy [760]), .D (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .CLK (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_9 (.Q (
        L1_2_L2_4_G2_MINI_ALU_BoothP_9), .QB (\$dummy [761]), .D (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .CLK (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_10 (.Q (
        L1_2_L2_4_G2_MINI_ALU_BoothP_10), .QB (\$dummy [762]), .D (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .CLK (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_11 (.Q (
        L1_2_L2_4_G2_MINI_ALU_BoothP_11), .QB (\$dummy [763]), .D (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .CLK (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_12 (.Q (
        L1_2_L2_4_G2_MINI_ALU_BoothP_12), .QB (\$dummy [764]), .D (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .CLK (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_13 (.Q (
        L1_2_L2_4_G2_MINI_ALU_BoothP_13), .QB (\$dummy [765]), .D (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .CLK (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_14 (.Q (
        L1_2_L2_4_G2_MINI_ALU_BoothP_14), .QB (\$dummy [766]), .D (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .CLK (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_15 (.Q (
        L1_2_L2_4_G2_MINI_ALU_BoothP_15), .QB (\$dummy [767]), .D (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .CLK (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_16 (.Q (
        L1_2_L2_4_G2_MINI_ALU_BoothP_16), .QB (\$dummy [768]), .D (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .CLK (
        L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    inv02 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix623 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624), .A (CLK)) ;
    inv02 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix625 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626), .A (CLK)) ;
    inv02 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix627 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628), .A (CLK)) ;
    inv02 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix643 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644), .A (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642)) ;
    xor2 L1_3_L2_0_G2_MINI_ALU_ix83 (.Y (L2Results_2__0), .A0 (L1Results_5__0), 
         .A1 (L1Results_4__0)) ;
    xnor2 L1_3_L2_0_G2_MINI_ALU_ix380 (.Y (L1_3_L2_0_G2_MINI_ALU_nx379), .A0 (
          L1_3_L2_0_G2_MINI_ALU_nx381), .A1 (L1_3_L2_0_G2_MINI_ALU_nx383)) ;
    nand02 L1_3_L2_0_G2_MINI_ALU_ix382 (.Y (L1_3_L2_0_G2_MINI_ALU_nx381), .A0 (
           L1_3_L2_0_G2_MINI_ALU_BoothOperand_0), .A1 (nx8204)) ;
    xnor2 L1_3_L2_0_G2_MINI_ALU_ix384 (.Y (L1_3_L2_0_G2_MINI_ALU_nx383), .A0 (
          L1_3_L2_0_G2_MINI_ALU_BoothOperand_1), .A1 (
          L1_3_L2_0_G2_MINI_ALU_BoothP_1)) ;
    inv01 L1_3_L2_0_G2_MINI_ALU_ix388 (.Y (L1_3_L2_0_G2_MINI_ALU_nx387), .A (
          L1_3_L2_0_G2_MINI_ALU_BoothP_2)) ;
    xnor2 L1_3_L2_0_G2_MINI_ALU_ix390 (.Y (L1_3_L2_0_G2_MINI_ALU_nx389), .A0 (
          L1_3_L2_0_G2_MINI_ALU_nx391), .A1 (L1_3_L2_0_G2_MINI_ALU_nx395)) ;
    aoi32 L1_3_L2_0_G2_MINI_ALU_ix392 (.Y (L1_3_L2_0_G2_MINI_ALU_nx391), .A0 (
          L1_3_L2_0_G2_MINI_ALU_BoothOperand_0), .A1 (nx8204), .A2 (
          L1_3_L2_0_G2_MINI_ALU_nx154), .B0 (L1_3_L2_0_G2_MINI_ALU_BoothP_1), .B1 (
          L1_3_L2_0_G2_MINI_ALU_BoothOperand_1)) ;
    xnor2 L1_3_L2_0_G2_MINI_ALU_ix396 (.Y (L1_3_L2_0_G2_MINI_ALU_nx395), .A0 (
          L1_3_L2_0_G2_MINI_ALU_BoothOperand_2), .A1 (
          L1_3_L2_0_G2_MINI_ALU_BoothP_2)) ;
    inv01 L1_3_L2_0_G2_MINI_ALU_ix400 (.Y (L1_3_L2_0_G2_MINI_ALU_nx399), .A (
          L1_3_L2_0_G2_MINI_ALU_BoothP_3)) ;
    xnor2 L1_3_L2_0_G2_MINI_ALU_ix402 (.Y (L1_3_L2_0_G2_MINI_ALU_nx401), .A0 (
          L1_3_L2_0_G2_MINI_ALU_nx403), .A1 (L1_3_L2_0_G2_MINI_ALU_nx405)) ;
    xnor2 L1_3_L2_0_G2_MINI_ALU_ix406 (.Y (L1_3_L2_0_G2_MINI_ALU_nx405), .A0 (
          L1_3_L2_0_G2_MINI_ALU_BoothOperand_3), .A1 (
          L1_3_L2_0_G2_MINI_ALU_BoothP_3)) ;
    inv01 L1_3_L2_0_G2_MINI_ALU_ix410 (.Y (L1_3_L2_0_G2_MINI_ALU_nx409), .A (
          L1_3_L2_0_G2_MINI_ALU_BoothP_4)) ;
    xnor2 L1_3_L2_0_G2_MINI_ALU_ix412 (.Y (L1_3_L2_0_G2_MINI_ALU_nx411), .A0 (
          L1_3_L2_0_G2_MINI_ALU_nx413), .A1 (L1_3_L2_0_G2_MINI_ALU_nx415)) ;
    xnor2 L1_3_L2_0_G2_MINI_ALU_ix416 (.Y (L1_3_L2_0_G2_MINI_ALU_nx415), .A0 (
          L1_3_L2_0_G2_MINI_ALU_BoothOperand_4), .A1 (
          L1_3_L2_0_G2_MINI_ALU_BoothP_4)) ;
    inv01 L1_3_L2_0_G2_MINI_ALU_ix420 (.Y (L1_3_L2_0_G2_MINI_ALU_nx419), .A (
          L1_3_L2_0_G2_MINI_ALU_BoothP_5)) ;
    xnor2 L1_3_L2_0_G2_MINI_ALU_ix422 (.Y (L1_3_L2_0_G2_MINI_ALU_nx421), .A0 (
          L1_3_L2_0_G2_MINI_ALU_nx423), .A1 (L1_3_L2_0_G2_MINI_ALU_nx425)) ;
    xnor2 L1_3_L2_0_G2_MINI_ALU_ix426 (.Y (L1_3_L2_0_G2_MINI_ALU_nx425), .A0 (
          L1_3_L2_0_G2_MINI_ALU_BoothOperand_5), .A1 (
          L1_3_L2_0_G2_MINI_ALU_BoothP_5)) ;
    inv01 L1_3_L2_0_G2_MINI_ALU_ix430 (.Y (L1_3_L2_0_G2_MINI_ALU_nx429), .A (
          L1_3_L2_0_G2_MINI_ALU_BoothP_6)) ;
    xnor2 L1_3_L2_0_G2_MINI_ALU_ix432 (.Y (L1_3_L2_0_G2_MINI_ALU_nx431), .A0 (
          L1_3_L2_0_G2_MINI_ALU_nx433), .A1 (L1_3_L2_0_G2_MINI_ALU_nx435)) ;
    xnor2 L1_3_L2_0_G2_MINI_ALU_ix436 (.Y (L1_3_L2_0_G2_MINI_ALU_nx435), .A0 (
          L1_3_L2_0_G2_MINI_ALU_BoothOperand_6), .A1 (
          L1_3_L2_0_G2_MINI_ALU_BoothP_6)) ;
    inv01 L1_3_L2_0_G2_MINI_ALU_ix440 (.Y (L1_3_L2_0_G2_MINI_ALU_nx439), .A (
          L1_3_L2_0_G2_MINI_ALU_BoothP_7)) ;
    xnor2 L1_3_L2_0_G2_MINI_ALU_ix442 (.Y (L1_3_L2_0_G2_MINI_ALU_nx441), .A0 (
          L1_3_L2_0_G2_MINI_ALU_nx443), .A1 (L1_3_L2_0_G2_MINI_ALU_nx445)) ;
    xnor2 L1_3_L2_0_G2_MINI_ALU_ix446 (.Y (L1_3_L2_0_G2_MINI_ALU_nx445), .A0 (
          L1_3_L2_0_G2_MINI_ALU_BoothOperand_7), .A1 (
          L1_3_L2_0_G2_MINI_ALU_BoothP_7)) ;
    inv01 L1_3_L2_0_G2_MINI_ALU_ix450 (.Y (L1_3_L2_0_G2_MINI_ALU_nx449), .A (
          L1_3_L2_0_G2_MINI_ALU_BoothP_8)) ;
    xnor2 L1_3_L2_0_G2_MINI_ALU_ix452 (.Y (L1_3_L2_0_G2_MINI_ALU_nx451), .A0 (
          L1_3_L2_0_G2_MINI_ALU_nx453), .A1 (L1_3_L2_0_G2_MINI_ALU_nx455)) ;
    xnor2 L1_3_L2_0_G2_MINI_ALU_ix456 (.Y (L1_3_L2_0_G2_MINI_ALU_nx455), .A0 (
          L1_3_L2_0_G2_MINI_ALU_BoothOperand_8), .A1 (
          L1_3_L2_0_G2_MINI_ALU_BoothP_8)) ;
    xor2 L1_3_L2_0_G2_MINI_ALU_ix317 (.Y (L1_3_L2_0_G2_MINI_ALU_nx316), .A0 (
         L1_3_L2_0_G2_MINI_ALU_nx461), .A1 (L1_3_L2_0_G2_MINI_ALU_nx463)) ;
    xnor2 L1_3_L2_0_G2_MINI_ALU_ix464 (.Y (L1_3_L2_0_G2_MINI_ALU_nx463), .A0 (
          L1_3_L2_0_G2_MINI_ALU_BoothOperand_9), .A1 (
          L1_3_L2_0_G2_MINI_ALU_BoothP_9)) ;
    xor2 L1_3_L2_0_G2_MINI_ALU_ix337 (.Y (L1_3_L2_0_G2_MINI_ALU_nx336), .A0 (
         L1_3_L2_0_G2_MINI_ALU_nx467), .A1 (L1_3_L2_0_G2_MINI_ALU_nx471)) ;
    inv01 L1_3_L2_0_G2_MINI_ALU_ix470 (.Y (L1_3_L2_0_G2_MINI_ALU_nx469), .A (
          L1_3_L2_0_G2_MINI_ALU_BoothP_9)) ;
    xnor2 L1_3_L2_0_G2_MINI_ALU_ix472 (.Y (L1_3_L2_0_G2_MINI_ALU_nx471), .A0 (
          L1_3_L2_0_G2_MINI_ALU_BoothOperand_10), .A1 (
          L1_3_L2_0_G2_MINI_ALU_BoothP_10)) ;
    xor2 L1_3_L2_0_G2_MINI_ALU_ix357 (.Y (L1_3_L2_0_G2_MINI_ALU_nx356), .A0 (
         L1_3_L2_0_G2_MINI_ALU_nx475), .A1 (L1_3_L2_0_G2_MINI_ALU_nx479)) ;
    inv01 L1_3_L2_0_G2_MINI_ALU_ix478 (.Y (L1_3_L2_0_G2_MINI_ALU_nx477), .A (
          L1_3_L2_0_G2_MINI_ALU_BoothP_10)) ;
    xnor2 L1_3_L2_0_G2_MINI_ALU_ix480 (.Y (L1_3_L2_0_G2_MINI_ALU_nx479), .A0 (
          L1_3_L2_0_G2_MINI_ALU_BoothOperand_11), .A1 (
          L1_3_L2_0_G2_MINI_ALU_BoothP_11)) ;
    xor2 L1_3_L2_0_G2_MINI_ALU_ix377 (.Y (L1_3_L2_0_G2_MINI_ALU_nx376), .A0 (
         L1_3_L2_0_G2_MINI_ALU_nx483), .A1 (L1_3_L2_0_G2_MINI_ALU_nx487)) ;
    inv01 L1_3_L2_0_G2_MINI_ALU_ix486 (.Y (L1_3_L2_0_G2_MINI_ALU_nx485), .A (
          L1_3_L2_0_G2_MINI_ALU_BoothP_11)) ;
    xnor2 L1_3_L2_0_G2_MINI_ALU_ix488 (.Y (L1_3_L2_0_G2_MINI_ALU_nx487), .A0 (
          L1_3_L2_0_G2_MINI_ALU_BoothOperand_12), .A1 (
          L1_3_L2_0_G2_MINI_ALU_BoothP_12)) ;
    xor2 L1_3_L2_0_G2_MINI_ALU_ix397 (.Y (L1_3_L2_0_G2_MINI_ALU_nx396), .A0 (
         L1_3_L2_0_G2_MINI_ALU_nx491), .A1 (L1_3_L2_0_G2_MINI_ALU_nx495)) ;
    inv01 L1_3_L2_0_G2_MINI_ALU_ix494 (.Y (L1_3_L2_0_G2_MINI_ALU_nx493), .A (
          L1_3_L2_0_G2_MINI_ALU_BoothP_12)) ;
    xnor2 L1_3_L2_0_G2_MINI_ALU_ix496 (.Y (L1_3_L2_0_G2_MINI_ALU_nx495), .A0 (
          L1_3_L2_0_G2_MINI_ALU_BoothOperand_13), .A1 (
          L1_3_L2_0_G2_MINI_ALU_BoothP_13)) ;
    xor2 L1_3_L2_0_G2_MINI_ALU_ix417 (.Y (L1_3_L2_0_G2_MINI_ALU_nx416), .A0 (
         L1_3_L2_0_G2_MINI_ALU_nx499), .A1 (L1_3_L2_0_G2_MINI_ALU_nx503)) ;
    inv01 L1_3_L2_0_G2_MINI_ALU_ix502 (.Y (L1_3_L2_0_G2_MINI_ALU_nx501), .A (
          L1_3_L2_0_G2_MINI_ALU_BoothP_13)) ;
    xnor2 L1_3_L2_0_G2_MINI_ALU_ix504 (.Y (L1_3_L2_0_G2_MINI_ALU_nx503), .A0 (
          L1_3_L2_0_G2_MINI_ALU_BoothOperand_14), .A1 (
          L1_3_L2_0_G2_MINI_ALU_BoothP_14)) ;
    xor2 L1_3_L2_0_G2_MINI_ALU_ix437 (.Y (L1_3_L2_0_G2_MINI_ALU_nx436), .A0 (
         L1_3_L2_0_G2_MINI_ALU_nx507), .A1 (L1_3_L2_0_G2_MINI_ALU_nx511)) ;
    inv01 L1_3_L2_0_G2_MINI_ALU_ix510 (.Y (L1_3_L2_0_G2_MINI_ALU_nx509), .A (
          L1_3_L2_0_G2_MINI_ALU_BoothP_14)) ;
    xnor2 L1_3_L2_0_G2_MINI_ALU_ix512 (.Y (L1_3_L2_0_G2_MINI_ALU_nx511), .A0 (
          L1_3_L2_0_G2_MINI_ALU_BoothOperand_15), .A1 (
          L1_3_L2_0_G2_MINI_ALU_BoothP_15)) ;
    xnor2 L1_3_L2_0_G2_MINI_ALU_ix457 (.Y (L1_3_L2_0_G2_MINI_ALU_nx456), .A0 (
          L1_3_L2_0_G2_MINI_ALU_nx515), .A1 (L1_3_L2_0_G2_MINI_ALU_nx454)) ;
    inv01 L1_3_L2_0_G2_MINI_ALU_ix518 (.Y (L1_3_L2_0_G2_MINI_ALU_nx517), .A (
          L1_3_L2_0_G2_MINI_ALU_BoothP_15)) ;
    xor2 L1_3_L2_0_G2_MINI_ALU_ix455 (.Y (L1_3_L2_0_G2_MINI_ALU_nx454), .A0 (
         L1_3_L2_0_G2_MINI_ALU_BoothOperand_16), .A1 (
         L1_3_L2_0_G2_MINI_ALU_BoothP_16)) ;
    mux21_ni L1_3_L2_0_G2_MINI_ALU_ix91 (.Y (L1FirstOperands_4__0), .A0 (
             L1_3_L2_0_G2_MINI_ALU_BoothP_1), .A1 (WindowDin_3__0__0), .S0 (
             Instr)) ;
    mux21_ni L1_3_L2_0_G2_MINI_ALU_ix99 (.Y (L1FirstOperands_4__1), .A0 (
             L1_3_L2_0_G2_MINI_ALU_BoothP_2), .A1 (WindowDin_3__0__1), .S0 (
             Instr)) ;
    mux21_ni L1_3_L2_0_G2_MINI_ALU_ix107 (.Y (L1FirstOperands_4__2), .A0 (
             L1_3_L2_0_G2_MINI_ALU_BoothP_3), .A1 (WindowDin_3__0__2), .S0 (
             Instr)) ;
    mux21_ni L1_3_L2_0_G2_MINI_ALU_ix115 (.Y (L1FirstOperands_4__3), .A0 (
             L1_3_L2_0_G2_MINI_ALU_BoothP_4), .A1 (WindowDin_3__0__3), .S0 (
             Instr)) ;
    mux21_ni L1_3_L2_0_G2_MINI_ALU_ix123 (.Y (L1FirstOperands_4__4), .A0 (
             L1_3_L2_0_G2_MINI_ALU_BoothP_5), .A1 (WindowDin_3__0__4), .S0 (
             Instr)) ;
    mux21_ni L1_3_L2_0_G2_MINI_ALU_ix131 (.Y (L1FirstOperands_4__5), .A0 (
             L1_3_L2_0_G2_MINI_ALU_BoothP_6), .A1 (WindowDin_3__0__5), .S0 (
             Instr)) ;
    mux21_ni L1_3_L2_0_G2_MINI_ALU_ix139 (.Y (L1FirstOperands_4__6), .A0 (
             L1_3_L2_0_G2_MINI_ALU_BoothP_7), .A1 (WindowDin_3__0__6), .S0 (
             Instr)) ;
    mux21_ni L1_3_L2_0_G2_MINI_ALU_ix147 (.Y (L1FirstOperands_4__7), .A0 (
             L1_3_L2_0_G2_MINI_ALU_BoothP_8), .A1 (WindowDin_3__0__7), .S0 (
             Instr)) ;
    xor2 L1_3_L2_0_G2_MINI_ALU_ix77 (.Y (L2Results_2__1), .A0 (
         L1_3_L2_0_G2_MINI_ALU_nx529), .A1 (L1_3_L2_0_G2_MINI_ALU_nx531)) ;
    nand02 L1_3_L2_0_G2_MINI_ALU_ix530 (.Y (L1_3_L2_0_G2_MINI_ALU_nx529), .A0 (
           L1Results_5__0), .A1 (L1Results_4__0)) ;
    xnor2 L1_3_L2_0_G2_MINI_ALU_ix532 (.Y (L1_3_L2_0_G2_MINI_ALU_nx531), .A0 (
          L1Results_5__1), .A1 (L1Results_4__1)) ;
    xor2 L1_3_L2_0_G2_MINI_ALU_ix75 (.Y (L2Results_2__2), .A0 (
         L1_3_L2_0_G2_MINI_ALU_nx534), .A1 (L1_3_L2_0_G2_MINI_ALU_nx537)) ;
    aoi32 L1_3_L2_0_G2_MINI_ALU_ix535 (.Y (L1_3_L2_0_G2_MINI_ALU_nx534), .A0 (
          L1Results_5__0), .A1 (L1Results_4__0), .A2 (L1_3_L2_0_G2_MINI_ALU_nx30
          ), .B0 (L1Results_4__1), .B1 (L1Results_5__1)) ;
    xnor2 L1_3_L2_0_G2_MINI_ALU_ix538 (.Y (L1_3_L2_0_G2_MINI_ALU_nx537), .A0 (
          L1Results_5__2), .A1 (L1Results_4__2)) ;
    xor2 L1_3_L2_0_G2_MINI_ALU_ix73 (.Y (L2Results_2__3), .A0 (
         L1_3_L2_0_G2_MINI_ALU_nx540), .A1 (L1_3_L2_0_G2_MINI_ALU_nx544)) ;
    aoi22 L1_3_L2_0_G2_MINI_ALU_ix541 (.Y (L1_3_L2_0_G2_MINI_ALU_nx540), .A0 (
          L1Results_4__2), .A1 (L1Results_5__2), .B0 (L1_3_L2_0_G2_MINI_ALU_nx40
          ), .B1 (L1_3_L2_0_G2_MINI_ALU_nx24)) ;
    xnor2 L1_3_L2_0_G2_MINI_ALU_ix545 (.Y (L1_3_L2_0_G2_MINI_ALU_nx544), .A0 (
          L1Results_5__3), .A1 (L1Results_4__3)) ;
    xor2 L1_3_L2_0_G2_MINI_ALU_ix71 (.Y (L2Results_2__4), .A0 (
         L1_3_L2_0_G2_MINI_ALU_nx547), .A1 (L1_3_L2_0_G2_MINI_ALU_nx551)) ;
    aoi22 L1_3_L2_0_G2_MINI_ALU_ix548 (.Y (L1_3_L2_0_G2_MINI_ALU_nx547), .A0 (
          L1Results_4__3), .A1 (L1Results_5__3), .B0 (L1_3_L2_0_G2_MINI_ALU_nx44
          ), .B1 (L1_3_L2_0_G2_MINI_ALU_nx18)) ;
    xnor2 L1_3_L2_0_G2_MINI_ALU_ix552 (.Y (L1_3_L2_0_G2_MINI_ALU_nx551), .A0 (
          L1Results_5__4), .A1 (L1Results_4__4)) ;
    xor2 L1_3_L2_0_G2_MINI_ALU_ix69 (.Y (L2Results_2__5), .A0 (
         L1_3_L2_0_G2_MINI_ALU_nx554), .A1 (L1_3_L2_0_G2_MINI_ALU_nx558)) ;
    aoi22 L1_3_L2_0_G2_MINI_ALU_ix555 (.Y (L1_3_L2_0_G2_MINI_ALU_nx554), .A0 (
          L1Results_4__4), .A1 (L1Results_5__4), .B0 (L1_3_L2_0_G2_MINI_ALU_nx48
          ), .B1 (L1_3_L2_0_G2_MINI_ALU_nx12)) ;
    xnor2 L1_3_L2_0_G2_MINI_ALU_ix559 (.Y (L1_3_L2_0_G2_MINI_ALU_nx558), .A0 (
          L1Results_5__5), .A1 (L1Results_4__5)) ;
    xor2 L1_3_L2_0_G2_MINI_ALU_ix67 (.Y (L2Results_2__6), .A0 (
         L1_3_L2_0_G2_MINI_ALU_nx561), .A1 (L1_3_L2_0_G2_MINI_ALU_nx565)) ;
    aoi22 L1_3_L2_0_G2_MINI_ALU_ix562 (.Y (L1_3_L2_0_G2_MINI_ALU_nx561), .A0 (
          L1Results_4__5), .A1 (L1Results_5__5), .B0 (L1_3_L2_0_G2_MINI_ALU_nx52
          ), .B1 (L1_3_L2_0_G2_MINI_ALU_nx6)) ;
    xnor2 L1_3_L2_0_G2_MINI_ALU_ix566 (.Y (L1_3_L2_0_G2_MINI_ALU_nx565), .A0 (
          L1Results_5__6), .A1 (L1Results_4__6)) ;
    xnor2 L1_3_L2_0_G2_MINI_ALU_ix65 (.Y (L2Results_2__7), .A0 (
          L1_3_L2_0_G2_MINI_ALU_nx568), .A1 (L1_3_L2_0_G2_MINI_ALU_nx62)) ;
    aoi22 L1_3_L2_0_G2_MINI_ALU_ix569 (.Y (L1_3_L2_0_G2_MINI_ALU_nx568), .A0 (
          L1Results_4__6), .A1 (L1Results_5__6), .B0 (L1_3_L2_0_G2_MINI_ALU_nx56
          ), .B1 (L1_3_L2_0_G2_MINI_ALU_nx0)) ;
    xor2 L1_3_L2_0_G2_MINI_ALU_ix63 (.Y (L1_3_L2_0_G2_MINI_ALU_nx62), .A0 (
         L1Results_5__7), .A1 (L1Results_4__7)) ;
    inv01 L1_3_L2_0_G2_MINI_ALU_ix155 (.Y (L1_3_L2_0_G2_MINI_ALU_nx154), .A (
          L1_3_L2_0_G2_MINI_ALU_nx383)) ;
    inv01 L1_3_L2_0_G2_MINI_ALU_ix57 (.Y (L1_3_L2_0_G2_MINI_ALU_nx56), .A (
          L1_3_L2_0_G2_MINI_ALU_nx561)) ;
    inv01 L1_3_L2_0_G2_MINI_ALU_ix53 (.Y (L1_3_L2_0_G2_MINI_ALU_nx52), .A (
          L1_3_L2_0_G2_MINI_ALU_nx554)) ;
    inv01 L1_3_L2_0_G2_MINI_ALU_ix49 (.Y (L1_3_L2_0_G2_MINI_ALU_nx48), .A (
          L1_3_L2_0_G2_MINI_ALU_nx547)) ;
    inv01 L1_3_L2_0_G2_MINI_ALU_ix45 (.Y (L1_3_L2_0_G2_MINI_ALU_nx44), .A (
          L1_3_L2_0_G2_MINI_ALU_nx540)) ;
    inv01 L1_3_L2_0_G2_MINI_ALU_ix41 (.Y (L1_3_L2_0_G2_MINI_ALU_nx40), .A (
          L1_3_L2_0_G2_MINI_ALU_nx534)) ;
    inv01 L1_3_L2_0_G2_MINI_ALU_ix31 (.Y (L1_3_L2_0_G2_MINI_ALU_nx30), .A (
          L1_3_L2_0_G2_MINI_ALU_nx531)) ;
    inv01 L1_3_L2_0_G2_MINI_ALU_ix25 (.Y (L1_3_L2_0_G2_MINI_ALU_nx24), .A (
          L1_3_L2_0_G2_MINI_ALU_nx537)) ;
    inv01 L1_3_L2_0_G2_MINI_ALU_ix19 (.Y (L1_3_L2_0_G2_MINI_ALU_nx18), .A (
          L1_3_L2_0_G2_MINI_ALU_nx544)) ;
    inv01 L1_3_L2_0_G2_MINI_ALU_ix13 (.Y (L1_3_L2_0_G2_MINI_ALU_nx12), .A (
          L1_3_L2_0_G2_MINI_ALU_nx551)) ;
    inv01 L1_3_L2_0_G2_MINI_ALU_ix7 (.Y (L1_3_L2_0_G2_MINI_ALU_nx6), .A (
          L1_3_L2_0_G2_MINI_ALU_nx558)) ;
    inv01 L1_3_L2_0_G2_MINI_ALU_ix1 (.Y (L1_3_L2_0_G2_MINI_ALU_nx0), .A (
          L1_3_L2_0_G2_MINI_ALU_nx565)) ;
    fake_gnd L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix216 (.Y (
             L1_3_L2_0_G2_MINI_ALU_WindowCellShiftedLeft_16)) ;
    nor02ii L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix81 (.Y (
            L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_nx80), .A0 (Instr), .A1 (Start)) ;
    aoi21 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix77 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_10), .A0 (
          FilterDin_3__0__1), .A1 (FilterDin_3__0__0), .B0 (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_nx4)) ;
    nor02_2x L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix5 (.Y (
             L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_nx4), .A0 (FilterDin_3__0__0), .A1 (
             FilterDin_3__0__1)) ;
    aoi21 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix67 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_11), .A0 (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_nx328), .A1 (FilterDin_3__0__2), .B0 (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_nx8)) ;
    nor03_2x L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix9 (.Y (
             L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_nx8), .A0 (FilterDin_3__0__2), .A1 (
             FilterDin_3__0__0), .A2 (FilterDin_3__0__1)) ;
    xnor2 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix59 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_12), .A0 (
          FilterDin_3__0__3), .A1 (L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_nx8)) ;
    xnor2 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix51 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_13), .A0 (
          FilterDin_3__0__4), .A1 (L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_nx12)) ;
    nor04 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix13 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_nx12), .A0 (FilterDin_3__0__3), .A1 (
          FilterDin_3__0__2), .A2 (FilterDin_3__0__0), .A3 (FilterDin_3__0__1)
          ) ;
    xnor2 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix43 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_14), .A0 (
          FilterDin_3__0__5), .A1 (L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_nx16)) ;
    nor02ii L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix17 (.Y (
            L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_nx16), .A0 (FilterDin_3__0__4), .A1 (
            L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_nx12)) ;
    xnor2 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix35 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_15), .A0 (
          FilterDin_3__0__6), .A1 (L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_nx20)) ;
    nor02ii L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix21 (.Y (
            L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_nx20), .A0 (FilterDin_3__0__5), .A1 (
            L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_nx16)) ;
    xnor2 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix27 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_16), .A0 (
          FilterDin_3__0__7), .A1 (L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_nx24)) ;
    nor02ii L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix25 (.Y (
            L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_nx24), .A0 (FilterDin_3__0__6), .A1 (
            L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_nx20)) ;
    inv01 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix329 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_nx328), .A (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_nx4)) ;
    inv02 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix383 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_nx384), .A (
          L1_3_L2_0_G2_MINI_ALU_BoothP_0)) ;
    dff L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_0 (.Q (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_0), .QB (\$dummy [769]), 
        .D (L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .CLK (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    nor02_2x L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix567 (.Y (
             L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566), .A0 (RST), .A1 (
             L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644)) ;
    dff L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_1 (.Q (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_1), .QB (\$dummy [770]), 
        .D (L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .CLK (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_2 (.Q (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_2), .QB (\$dummy [771]), 
        .D (L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .CLK (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_3 (.Q (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_3), .QB (\$dummy [772]), 
        .D (L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .CLK (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_4 (.Q (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_4), .QB (\$dummy [773]), 
        .D (L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .CLK (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_5 (.Q (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_5), .QB (\$dummy [774]), 
        .D (L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .CLK (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_6 (.Q (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_6), .QB (\$dummy [775]), 
        .D (L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .CLK (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_7 (.Q (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_7), .QB (\$dummy [776]), 
        .D (L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .CLK (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_8 (.Q (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_8), .QB (\$dummy [777]), 
        .D (L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .CLK (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_9 (.Q (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_9), .QB (\$dummy [778]), 
        .D (L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .CLK (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_10 (.Q (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_10), .QB (\$dummy [779])
        , .D (L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .CLK (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_11 (.Q (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_11), .QB (\$dummy [780])
        , .D (L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .CLK (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_12 (.Q (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_12), .QB (\$dummy [781])
        , .D (L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .CLK (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_13 (.Q (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_13), .QB (\$dummy [782])
        , .D (L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .CLK (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_14 (.Q (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_14), .QB (\$dummy [783])
        , .D (L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .CLK (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_15 (.Q (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_15), .QB (\$dummy [784])
        , .D (L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .CLK (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_16 (.Q (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_16), .QB (\$dummy [785])
        , .D (L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .CLK (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    inv02 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix623 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624), .A (CLK)) ;
    inv02 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix625 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626), .A (CLK)) ;
    inv02 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix627 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628), .A (CLK)) ;
    inv02 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix643 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644), .A (nx8218)) ;
    dff L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_0 (.Q (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_0), .QB (\$dummy [786]), 
        .D (L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .CLK (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    nor02_2x L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix567 (.Y (
             L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566), .A0 (RST), .A1 (
             L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644)) ;
    dff L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_1 (.Q (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_1), .QB (\$dummy [787]), 
        .D (L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .CLK (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_2 (.Q (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_2), .QB (\$dummy [788]), 
        .D (L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .CLK (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_3 (.Q (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_3), .QB (\$dummy [789]), 
        .D (L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .CLK (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_4 (.Q (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_4), .QB (\$dummy [790]), 
        .D (L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .CLK (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_5 (.Q (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_5), .QB (\$dummy [791]), 
        .D (L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .CLK (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_6 (.Q (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_6), .QB (\$dummy [792]), 
        .D (L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .CLK (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_7 (.Q (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_7), .QB (\$dummy [793]), 
        .D (L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .CLK (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_8 (.Q (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_8), .QB (\$dummy [794]), 
        .D (L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .CLK (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_9 (.Q (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_9), .QB (\$dummy [795]), 
        .D (L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .CLK (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_10 (.Q (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_10), .QB (\$dummy [796])
        , .D (L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .CLK (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_11 (.Q (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_11), .QB (\$dummy [797])
        , .D (L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .CLK (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_12 (.Q (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_12), .QB (\$dummy [798])
        , .D (L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .CLK (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_13 (.Q (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_13), .QB (\$dummy [799])
        , .D (L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .CLK (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_14 (.Q (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_14), .QB (\$dummy [800])
        , .D (L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .CLK (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_15 (.Q (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_15), .QB (\$dummy [801])
        , .D (L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .CLK (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_16 (.Q (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_16), .QB (\$dummy [802])
        , .D (L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .CLK (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    inv02 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix623 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624), .A (CLK)) ;
    inv02 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix625 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626), .A (CLK)) ;
    inv02 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix627 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628), .A (CLK)) ;
    inv02 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix643 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644), .A (nx8224)) ;
    dff L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_0 (.Q (
        L1_3_L2_0_G2_MINI_ALU_BoothP_0), .QB (\$dummy [803]), .D (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .CLK (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    nor02_2x L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix567 (.Y (
             L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566), .A0 (RST), .A1 (
             L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    dff L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_1 (.Q (
        L1_3_L2_0_G2_MINI_ALU_BoothP_1), .QB (\$dummy [804]), .D (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .CLK (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_2 (.Q (
        L1_3_L2_0_G2_MINI_ALU_BoothP_2), .QB (\$dummy [805]), .D (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .CLK (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_3 (.Q (
        L1_3_L2_0_G2_MINI_ALU_BoothP_3), .QB (\$dummy [806]), .D (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .CLK (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_4 (.Q (
        L1_3_L2_0_G2_MINI_ALU_BoothP_4), .QB (\$dummy [807]), .D (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .CLK (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_5 (.Q (
        L1_3_L2_0_G2_MINI_ALU_BoothP_5), .QB (\$dummy [808]), .D (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .CLK (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_6 (.Q (
        L1_3_L2_0_G2_MINI_ALU_BoothP_6), .QB (\$dummy [809]), .D (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .CLK (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_7 (.Q (
        L1_3_L2_0_G2_MINI_ALU_BoothP_7), .QB (\$dummy [810]), .D (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .CLK (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_8 (.Q (
        L1_3_L2_0_G2_MINI_ALU_BoothP_8), .QB (\$dummy [811]), .D (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .CLK (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_9 (.Q (
        L1_3_L2_0_G2_MINI_ALU_BoothP_9), .QB (\$dummy [812]), .D (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .CLK (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_10 (.Q (
        L1_3_L2_0_G2_MINI_ALU_BoothP_10), .QB (\$dummy [813]), .D (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .CLK (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_11 (.Q (
        L1_3_L2_0_G2_MINI_ALU_BoothP_11), .QB (\$dummy [814]), .D (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .CLK (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_12 (.Q (
        L1_3_L2_0_G2_MINI_ALU_BoothP_12), .QB (\$dummy [815]), .D (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .CLK (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_13 (.Q (
        L1_3_L2_0_G2_MINI_ALU_BoothP_13), .QB (\$dummy [816]), .D (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .CLK (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_14 (.Q (
        L1_3_L2_0_G2_MINI_ALU_BoothP_14), .QB (\$dummy [817]), .D (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .CLK (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_15 (.Q (
        L1_3_L2_0_G2_MINI_ALU_BoothP_15), .QB (\$dummy [818]), .D (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .CLK (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_16 (.Q (
        L1_3_L2_0_G2_MINI_ALU_BoothP_16), .QB (\$dummy [819]), .D (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .CLK (
        L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    inv02 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix623 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624), .A (CLK)) ;
    inv02 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix625 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626), .A (CLK)) ;
    inv02 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix627 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628), .A (CLK)) ;
    inv02 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix643 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644), .A (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642)) ;
    xor2 L1_3_L2_1_G2_MINI_ALU_ix83 (.Y (L2Results_3__0), .A0 (L1Results_7__0), 
         .A1 (L1Results_6__0)) ;
    xnor2 L1_3_L2_1_G2_MINI_ALU_ix380 (.Y (L1_3_L2_1_G2_MINI_ALU_nx379), .A0 (
          L1_3_L2_1_G2_MINI_ALU_nx381), .A1 (L1_3_L2_1_G2_MINI_ALU_nx383)) ;
    nand02 L1_3_L2_1_G2_MINI_ALU_ix382 (.Y (L1_3_L2_1_G2_MINI_ALU_nx381), .A0 (
           L1_3_L2_1_G2_MINI_ALU_BoothOperand_0), .A1 (nx8244)) ;
    xnor2 L1_3_L2_1_G2_MINI_ALU_ix384 (.Y (L1_3_L2_1_G2_MINI_ALU_nx383), .A0 (
          L1_3_L2_1_G2_MINI_ALU_BoothOperand_1), .A1 (
          L1_3_L2_1_G2_MINI_ALU_BoothP_1)) ;
    inv01 L1_3_L2_1_G2_MINI_ALU_ix388 (.Y (L1_3_L2_1_G2_MINI_ALU_nx387), .A (
          L1_3_L2_1_G2_MINI_ALU_BoothP_2)) ;
    xnor2 L1_3_L2_1_G2_MINI_ALU_ix390 (.Y (L1_3_L2_1_G2_MINI_ALU_nx389), .A0 (
          L1_3_L2_1_G2_MINI_ALU_nx391), .A1 (L1_3_L2_1_G2_MINI_ALU_nx395)) ;
    aoi32 L1_3_L2_1_G2_MINI_ALU_ix392 (.Y (L1_3_L2_1_G2_MINI_ALU_nx391), .A0 (
          L1_3_L2_1_G2_MINI_ALU_BoothOperand_0), .A1 (nx8244), .A2 (
          L1_3_L2_1_G2_MINI_ALU_nx154), .B0 (L1_3_L2_1_G2_MINI_ALU_BoothP_1), .B1 (
          L1_3_L2_1_G2_MINI_ALU_BoothOperand_1)) ;
    xnor2 L1_3_L2_1_G2_MINI_ALU_ix396 (.Y (L1_3_L2_1_G2_MINI_ALU_nx395), .A0 (
          L1_3_L2_1_G2_MINI_ALU_BoothOperand_2), .A1 (
          L1_3_L2_1_G2_MINI_ALU_BoothP_2)) ;
    inv01 L1_3_L2_1_G2_MINI_ALU_ix400 (.Y (L1_3_L2_1_G2_MINI_ALU_nx399), .A (
          L1_3_L2_1_G2_MINI_ALU_BoothP_3)) ;
    xnor2 L1_3_L2_1_G2_MINI_ALU_ix402 (.Y (L1_3_L2_1_G2_MINI_ALU_nx401), .A0 (
          L1_3_L2_1_G2_MINI_ALU_nx403), .A1 (L1_3_L2_1_G2_MINI_ALU_nx405)) ;
    xnor2 L1_3_L2_1_G2_MINI_ALU_ix406 (.Y (L1_3_L2_1_G2_MINI_ALU_nx405), .A0 (
          L1_3_L2_1_G2_MINI_ALU_BoothOperand_3), .A1 (
          L1_3_L2_1_G2_MINI_ALU_BoothP_3)) ;
    inv01 L1_3_L2_1_G2_MINI_ALU_ix410 (.Y (L1_3_L2_1_G2_MINI_ALU_nx409), .A (
          L1_3_L2_1_G2_MINI_ALU_BoothP_4)) ;
    xnor2 L1_3_L2_1_G2_MINI_ALU_ix412 (.Y (L1_3_L2_1_G2_MINI_ALU_nx411), .A0 (
          L1_3_L2_1_G2_MINI_ALU_nx413), .A1 (L1_3_L2_1_G2_MINI_ALU_nx415)) ;
    xnor2 L1_3_L2_1_G2_MINI_ALU_ix416 (.Y (L1_3_L2_1_G2_MINI_ALU_nx415), .A0 (
          L1_3_L2_1_G2_MINI_ALU_BoothOperand_4), .A1 (
          L1_3_L2_1_G2_MINI_ALU_BoothP_4)) ;
    inv01 L1_3_L2_1_G2_MINI_ALU_ix420 (.Y (L1_3_L2_1_G2_MINI_ALU_nx419), .A (
          L1_3_L2_1_G2_MINI_ALU_BoothP_5)) ;
    xnor2 L1_3_L2_1_G2_MINI_ALU_ix422 (.Y (L1_3_L2_1_G2_MINI_ALU_nx421), .A0 (
          L1_3_L2_1_G2_MINI_ALU_nx423), .A1 (L1_3_L2_1_G2_MINI_ALU_nx425)) ;
    xnor2 L1_3_L2_1_G2_MINI_ALU_ix426 (.Y (L1_3_L2_1_G2_MINI_ALU_nx425), .A0 (
          L1_3_L2_1_G2_MINI_ALU_BoothOperand_5), .A1 (
          L1_3_L2_1_G2_MINI_ALU_BoothP_5)) ;
    inv01 L1_3_L2_1_G2_MINI_ALU_ix430 (.Y (L1_3_L2_1_G2_MINI_ALU_nx429), .A (
          L1_3_L2_1_G2_MINI_ALU_BoothP_6)) ;
    xnor2 L1_3_L2_1_G2_MINI_ALU_ix432 (.Y (L1_3_L2_1_G2_MINI_ALU_nx431), .A0 (
          L1_3_L2_1_G2_MINI_ALU_nx433), .A1 (L1_3_L2_1_G2_MINI_ALU_nx435)) ;
    xnor2 L1_3_L2_1_G2_MINI_ALU_ix436 (.Y (L1_3_L2_1_G2_MINI_ALU_nx435), .A0 (
          L1_3_L2_1_G2_MINI_ALU_BoothOperand_6), .A1 (
          L1_3_L2_1_G2_MINI_ALU_BoothP_6)) ;
    inv01 L1_3_L2_1_G2_MINI_ALU_ix440 (.Y (L1_3_L2_1_G2_MINI_ALU_nx439), .A (
          L1_3_L2_1_G2_MINI_ALU_BoothP_7)) ;
    xnor2 L1_3_L2_1_G2_MINI_ALU_ix442 (.Y (L1_3_L2_1_G2_MINI_ALU_nx441), .A0 (
          L1_3_L2_1_G2_MINI_ALU_nx443), .A1 (L1_3_L2_1_G2_MINI_ALU_nx445)) ;
    xnor2 L1_3_L2_1_G2_MINI_ALU_ix446 (.Y (L1_3_L2_1_G2_MINI_ALU_nx445), .A0 (
          L1_3_L2_1_G2_MINI_ALU_BoothOperand_7), .A1 (
          L1_3_L2_1_G2_MINI_ALU_BoothP_7)) ;
    inv01 L1_3_L2_1_G2_MINI_ALU_ix450 (.Y (L1_3_L2_1_G2_MINI_ALU_nx449), .A (
          L1_3_L2_1_G2_MINI_ALU_BoothP_8)) ;
    xnor2 L1_3_L2_1_G2_MINI_ALU_ix452 (.Y (L1_3_L2_1_G2_MINI_ALU_nx451), .A0 (
          L1_3_L2_1_G2_MINI_ALU_nx453), .A1 (L1_3_L2_1_G2_MINI_ALU_nx455)) ;
    xnor2 L1_3_L2_1_G2_MINI_ALU_ix456 (.Y (L1_3_L2_1_G2_MINI_ALU_nx455), .A0 (
          L1_3_L2_1_G2_MINI_ALU_BoothOperand_8), .A1 (
          L1_3_L2_1_G2_MINI_ALU_BoothP_8)) ;
    xor2 L1_3_L2_1_G2_MINI_ALU_ix317 (.Y (L1_3_L2_1_G2_MINI_ALU_nx316), .A0 (
         L1_3_L2_1_G2_MINI_ALU_nx461), .A1 (L1_3_L2_1_G2_MINI_ALU_nx463)) ;
    xnor2 L1_3_L2_1_G2_MINI_ALU_ix464 (.Y (L1_3_L2_1_G2_MINI_ALU_nx463), .A0 (
          L1_3_L2_1_G2_MINI_ALU_BoothOperand_9), .A1 (
          L1_3_L2_1_G2_MINI_ALU_BoothP_9)) ;
    xor2 L1_3_L2_1_G2_MINI_ALU_ix337 (.Y (L1_3_L2_1_G2_MINI_ALU_nx336), .A0 (
         L1_3_L2_1_G2_MINI_ALU_nx467), .A1 (L1_3_L2_1_G2_MINI_ALU_nx471)) ;
    inv01 L1_3_L2_1_G2_MINI_ALU_ix470 (.Y (L1_3_L2_1_G2_MINI_ALU_nx469), .A (
          L1_3_L2_1_G2_MINI_ALU_BoothP_9)) ;
    xnor2 L1_3_L2_1_G2_MINI_ALU_ix472 (.Y (L1_3_L2_1_G2_MINI_ALU_nx471), .A0 (
          L1_3_L2_1_G2_MINI_ALU_BoothOperand_10), .A1 (
          L1_3_L2_1_G2_MINI_ALU_BoothP_10)) ;
    xor2 L1_3_L2_1_G2_MINI_ALU_ix357 (.Y (L1_3_L2_1_G2_MINI_ALU_nx356), .A0 (
         L1_3_L2_1_G2_MINI_ALU_nx475), .A1 (L1_3_L2_1_G2_MINI_ALU_nx479)) ;
    inv01 L1_3_L2_1_G2_MINI_ALU_ix478 (.Y (L1_3_L2_1_G2_MINI_ALU_nx477), .A (
          L1_3_L2_1_G2_MINI_ALU_BoothP_10)) ;
    xnor2 L1_3_L2_1_G2_MINI_ALU_ix480 (.Y (L1_3_L2_1_G2_MINI_ALU_nx479), .A0 (
          L1_3_L2_1_G2_MINI_ALU_BoothOperand_11), .A1 (
          L1_3_L2_1_G2_MINI_ALU_BoothP_11)) ;
    xor2 L1_3_L2_1_G2_MINI_ALU_ix377 (.Y (L1_3_L2_1_G2_MINI_ALU_nx376), .A0 (
         L1_3_L2_1_G2_MINI_ALU_nx483), .A1 (L1_3_L2_1_G2_MINI_ALU_nx487)) ;
    inv01 L1_3_L2_1_G2_MINI_ALU_ix486 (.Y (L1_3_L2_1_G2_MINI_ALU_nx485), .A (
          L1_3_L2_1_G2_MINI_ALU_BoothP_11)) ;
    xnor2 L1_3_L2_1_G2_MINI_ALU_ix488 (.Y (L1_3_L2_1_G2_MINI_ALU_nx487), .A0 (
          L1_3_L2_1_G2_MINI_ALU_BoothOperand_12), .A1 (
          L1_3_L2_1_G2_MINI_ALU_BoothP_12)) ;
    xor2 L1_3_L2_1_G2_MINI_ALU_ix397 (.Y (L1_3_L2_1_G2_MINI_ALU_nx396), .A0 (
         L1_3_L2_1_G2_MINI_ALU_nx491), .A1 (L1_3_L2_1_G2_MINI_ALU_nx495)) ;
    inv01 L1_3_L2_1_G2_MINI_ALU_ix494 (.Y (L1_3_L2_1_G2_MINI_ALU_nx493), .A (
          L1_3_L2_1_G2_MINI_ALU_BoothP_12)) ;
    xnor2 L1_3_L2_1_G2_MINI_ALU_ix496 (.Y (L1_3_L2_1_G2_MINI_ALU_nx495), .A0 (
          L1_3_L2_1_G2_MINI_ALU_BoothOperand_13), .A1 (
          L1_3_L2_1_G2_MINI_ALU_BoothP_13)) ;
    xor2 L1_3_L2_1_G2_MINI_ALU_ix417 (.Y (L1_3_L2_1_G2_MINI_ALU_nx416), .A0 (
         L1_3_L2_1_G2_MINI_ALU_nx499), .A1 (L1_3_L2_1_G2_MINI_ALU_nx503)) ;
    inv01 L1_3_L2_1_G2_MINI_ALU_ix502 (.Y (L1_3_L2_1_G2_MINI_ALU_nx501), .A (
          L1_3_L2_1_G2_MINI_ALU_BoothP_13)) ;
    xnor2 L1_3_L2_1_G2_MINI_ALU_ix504 (.Y (L1_3_L2_1_G2_MINI_ALU_nx503), .A0 (
          L1_3_L2_1_G2_MINI_ALU_BoothOperand_14), .A1 (
          L1_3_L2_1_G2_MINI_ALU_BoothP_14)) ;
    xor2 L1_3_L2_1_G2_MINI_ALU_ix437 (.Y (L1_3_L2_1_G2_MINI_ALU_nx436), .A0 (
         L1_3_L2_1_G2_MINI_ALU_nx507), .A1 (L1_3_L2_1_G2_MINI_ALU_nx511)) ;
    inv01 L1_3_L2_1_G2_MINI_ALU_ix510 (.Y (L1_3_L2_1_G2_MINI_ALU_nx509), .A (
          L1_3_L2_1_G2_MINI_ALU_BoothP_14)) ;
    xnor2 L1_3_L2_1_G2_MINI_ALU_ix512 (.Y (L1_3_L2_1_G2_MINI_ALU_nx511), .A0 (
          L1_3_L2_1_G2_MINI_ALU_BoothOperand_15), .A1 (
          L1_3_L2_1_G2_MINI_ALU_BoothP_15)) ;
    xnor2 L1_3_L2_1_G2_MINI_ALU_ix457 (.Y (L1_3_L2_1_G2_MINI_ALU_nx456), .A0 (
          L1_3_L2_1_G2_MINI_ALU_nx515), .A1 (L1_3_L2_1_G2_MINI_ALU_nx454)) ;
    inv01 L1_3_L2_1_G2_MINI_ALU_ix518 (.Y (L1_3_L2_1_G2_MINI_ALU_nx517), .A (
          L1_3_L2_1_G2_MINI_ALU_BoothP_15)) ;
    xor2 L1_3_L2_1_G2_MINI_ALU_ix455 (.Y (L1_3_L2_1_G2_MINI_ALU_nx454), .A0 (
         L1_3_L2_1_G2_MINI_ALU_BoothOperand_16), .A1 (
         L1_3_L2_1_G2_MINI_ALU_BoothP_16)) ;
    mux21_ni L1_3_L2_1_G2_MINI_ALU_ix91 (.Y (L1FirstOperands_6__0), .A0 (
             L1_3_L2_1_G2_MINI_ALU_BoothP_1), .A1 (WindowDin_3__1__0), .S0 (
             Instr)) ;
    mux21_ni L1_3_L2_1_G2_MINI_ALU_ix99 (.Y (L1FirstOperands_6__1), .A0 (
             L1_3_L2_1_G2_MINI_ALU_BoothP_2), .A1 (WindowDin_3__1__1), .S0 (
             Instr)) ;
    mux21_ni L1_3_L2_1_G2_MINI_ALU_ix107 (.Y (L1FirstOperands_6__2), .A0 (
             L1_3_L2_1_G2_MINI_ALU_BoothP_3), .A1 (WindowDin_3__1__2), .S0 (
             Instr)) ;
    mux21_ni L1_3_L2_1_G2_MINI_ALU_ix115 (.Y (L1FirstOperands_6__3), .A0 (
             L1_3_L2_1_G2_MINI_ALU_BoothP_4), .A1 (WindowDin_3__1__3), .S0 (
             Instr)) ;
    mux21_ni L1_3_L2_1_G2_MINI_ALU_ix123 (.Y (L1FirstOperands_6__4), .A0 (
             L1_3_L2_1_G2_MINI_ALU_BoothP_5), .A1 (WindowDin_3__1__4), .S0 (
             Instr)) ;
    mux21_ni L1_3_L2_1_G2_MINI_ALU_ix131 (.Y (L1FirstOperands_6__5), .A0 (
             L1_3_L2_1_G2_MINI_ALU_BoothP_6), .A1 (WindowDin_3__1__5), .S0 (
             Instr)) ;
    mux21_ni L1_3_L2_1_G2_MINI_ALU_ix139 (.Y (L1FirstOperands_6__6), .A0 (
             L1_3_L2_1_G2_MINI_ALU_BoothP_7), .A1 (WindowDin_3__1__6), .S0 (
             Instr)) ;
    mux21_ni L1_3_L2_1_G2_MINI_ALU_ix147 (.Y (L1FirstOperands_6__7), .A0 (
             L1_3_L2_1_G2_MINI_ALU_BoothP_8), .A1 (WindowDin_3__1__7), .S0 (
             Instr)) ;
    xor2 L1_3_L2_1_G2_MINI_ALU_ix77 (.Y (L2Results_3__1), .A0 (
         L1_3_L2_1_G2_MINI_ALU_nx529), .A1 (L1_3_L2_1_G2_MINI_ALU_nx531)) ;
    nand02 L1_3_L2_1_G2_MINI_ALU_ix530 (.Y (L1_3_L2_1_G2_MINI_ALU_nx529), .A0 (
           L1Results_7__0), .A1 (L1Results_6__0)) ;
    xnor2 L1_3_L2_1_G2_MINI_ALU_ix532 (.Y (L1_3_L2_1_G2_MINI_ALU_nx531), .A0 (
          L1Results_7__1), .A1 (L1Results_6__1)) ;
    xor2 L1_3_L2_1_G2_MINI_ALU_ix75 (.Y (L2Results_3__2), .A0 (
         L1_3_L2_1_G2_MINI_ALU_nx534), .A1 (L1_3_L2_1_G2_MINI_ALU_nx537)) ;
    aoi32 L1_3_L2_1_G2_MINI_ALU_ix535 (.Y (L1_3_L2_1_G2_MINI_ALU_nx534), .A0 (
          L1Results_7__0), .A1 (L1Results_6__0), .A2 (L1_3_L2_1_G2_MINI_ALU_nx30
          ), .B0 (L1Results_6__1), .B1 (L1Results_7__1)) ;
    xnor2 L1_3_L2_1_G2_MINI_ALU_ix538 (.Y (L1_3_L2_1_G2_MINI_ALU_nx537), .A0 (
          L1Results_7__2), .A1 (L1Results_6__2)) ;
    xor2 L1_3_L2_1_G2_MINI_ALU_ix73 (.Y (L2Results_3__3), .A0 (
         L1_3_L2_1_G2_MINI_ALU_nx540), .A1 (L1_3_L2_1_G2_MINI_ALU_nx544)) ;
    aoi22 L1_3_L2_1_G2_MINI_ALU_ix541 (.Y (L1_3_L2_1_G2_MINI_ALU_nx540), .A0 (
          L1Results_6__2), .A1 (L1Results_7__2), .B0 (L1_3_L2_1_G2_MINI_ALU_nx40
          ), .B1 (L1_3_L2_1_G2_MINI_ALU_nx24)) ;
    xnor2 L1_3_L2_1_G2_MINI_ALU_ix545 (.Y (L1_3_L2_1_G2_MINI_ALU_nx544), .A0 (
          L1Results_7__3), .A1 (L1Results_6__3)) ;
    xor2 L1_3_L2_1_G2_MINI_ALU_ix71 (.Y (L2Results_3__4), .A0 (
         L1_3_L2_1_G2_MINI_ALU_nx547), .A1 (L1_3_L2_1_G2_MINI_ALU_nx551)) ;
    aoi22 L1_3_L2_1_G2_MINI_ALU_ix548 (.Y (L1_3_L2_1_G2_MINI_ALU_nx547), .A0 (
          L1Results_6__3), .A1 (L1Results_7__3), .B0 (L1_3_L2_1_G2_MINI_ALU_nx44
          ), .B1 (L1_3_L2_1_G2_MINI_ALU_nx18)) ;
    xnor2 L1_3_L2_1_G2_MINI_ALU_ix552 (.Y (L1_3_L2_1_G2_MINI_ALU_nx551), .A0 (
          L1Results_7__4), .A1 (L1Results_6__4)) ;
    xor2 L1_3_L2_1_G2_MINI_ALU_ix69 (.Y (L2Results_3__5), .A0 (
         L1_3_L2_1_G2_MINI_ALU_nx554), .A1 (L1_3_L2_1_G2_MINI_ALU_nx558)) ;
    aoi22 L1_3_L2_1_G2_MINI_ALU_ix555 (.Y (L1_3_L2_1_G2_MINI_ALU_nx554), .A0 (
          L1Results_6__4), .A1 (L1Results_7__4), .B0 (L1_3_L2_1_G2_MINI_ALU_nx48
          ), .B1 (L1_3_L2_1_G2_MINI_ALU_nx12)) ;
    xnor2 L1_3_L2_1_G2_MINI_ALU_ix559 (.Y (L1_3_L2_1_G2_MINI_ALU_nx558), .A0 (
          L1Results_7__5), .A1 (L1Results_6__5)) ;
    xor2 L1_3_L2_1_G2_MINI_ALU_ix67 (.Y (L2Results_3__6), .A0 (
         L1_3_L2_1_G2_MINI_ALU_nx561), .A1 (L1_3_L2_1_G2_MINI_ALU_nx565)) ;
    aoi22 L1_3_L2_1_G2_MINI_ALU_ix562 (.Y (L1_3_L2_1_G2_MINI_ALU_nx561), .A0 (
          L1Results_6__5), .A1 (L1Results_7__5), .B0 (L1_3_L2_1_G2_MINI_ALU_nx52
          ), .B1 (L1_3_L2_1_G2_MINI_ALU_nx6)) ;
    xnor2 L1_3_L2_1_G2_MINI_ALU_ix566 (.Y (L1_3_L2_1_G2_MINI_ALU_nx565), .A0 (
          L1Results_7__6), .A1 (L1Results_6__6)) ;
    xnor2 L1_3_L2_1_G2_MINI_ALU_ix65 (.Y (L2Results_3__7), .A0 (
          L1_3_L2_1_G2_MINI_ALU_nx568), .A1 (L1_3_L2_1_G2_MINI_ALU_nx62)) ;
    aoi22 L1_3_L2_1_G2_MINI_ALU_ix569 (.Y (L1_3_L2_1_G2_MINI_ALU_nx568), .A0 (
          L1Results_6__6), .A1 (L1Results_7__6), .B0 (L1_3_L2_1_G2_MINI_ALU_nx56
          ), .B1 (L1_3_L2_1_G2_MINI_ALU_nx0)) ;
    xor2 L1_3_L2_1_G2_MINI_ALU_ix63 (.Y (L1_3_L2_1_G2_MINI_ALU_nx62), .A0 (
         L1Results_7__7), .A1 (L1Results_6__7)) ;
    inv01 L1_3_L2_1_G2_MINI_ALU_ix155 (.Y (L1_3_L2_1_G2_MINI_ALU_nx154), .A (
          L1_3_L2_1_G2_MINI_ALU_nx383)) ;
    inv01 L1_3_L2_1_G2_MINI_ALU_ix57 (.Y (L1_3_L2_1_G2_MINI_ALU_nx56), .A (
          L1_3_L2_1_G2_MINI_ALU_nx561)) ;
    inv01 L1_3_L2_1_G2_MINI_ALU_ix53 (.Y (L1_3_L2_1_G2_MINI_ALU_nx52), .A (
          L1_3_L2_1_G2_MINI_ALU_nx554)) ;
    inv01 L1_3_L2_1_G2_MINI_ALU_ix49 (.Y (L1_3_L2_1_G2_MINI_ALU_nx48), .A (
          L1_3_L2_1_G2_MINI_ALU_nx547)) ;
    inv01 L1_3_L2_1_G2_MINI_ALU_ix45 (.Y (L1_3_L2_1_G2_MINI_ALU_nx44), .A (
          L1_3_L2_1_G2_MINI_ALU_nx540)) ;
    inv01 L1_3_L2_1_G2_MINI_ALU_ix41 (.Y (L1_3_L2_1_G2_MINI_ALU_nx40), .A (
          L1_3_L2_1_G2_MINI_ALU_nx534)) ;
    inv01 L1_3_L2_1_G2_MINI_ALU_ix31 (.Y (L1_3_L2_1_G2_MINI_ALU_nx30), .A (
          L1_3_L2_1_G2_MINI_ALU_nx531)) ;
    inv01 L1_3_L2_1_G2_MINI_ALU_ix25 (.Y (L1_3_L2_1_G2_MINI_ALU_nx24), .A (
          L1_3_L2_1_G2_MINI_ALU_nx537)) ;
    inv01 L1_3_L2_1_G2_MINI_ALU_ix19 (.Y (L1_3_L2_1_G2_MINI_ALU_nx18), .A (
          L1_3_L2_1_G2_MINI_ALU_nx544)) ;
    inv01 L1_3_L2_1_G2_MINI_ALU_ix13 (.Y (L1_3_L2_1_G2_MINI_ALU_nx12), .A (
          L1_3_L2_1_G2_MINI_ALU_nx551)) ;
    inv01 L1_3_L2_1_G2_MINI_ALU_ix7 (.Y (L1_3_L2_1_G2_MINI_ALU_nx6), .A (
          L1_3_L2_1_G2_MINI_ALU_nx558)) ;
    inv01 L1_3_L2_1_G2_MINI_ALU_ix1 (.Y (L1_3_L2_1_G2_MINI_ALU_nx0), .A (
          L1_3_L2_1_G2_MINI_ALU_nx565)) ;
    fake_gnd L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix216 (.Y (
             L1_3_L2_1_G2_MINI_ALU_WindowCellShiftedLeft_16)) ;
    nor02ii L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix81 (.Y (
            L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_nx80), .A0 (Instr), .A1 (Start)) ;
    aoi21 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix77 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_10), .A0 (
          FilterDin_3__1__1), .A1 (FilterDin_3__1__0), .B0 (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_nx4)) ;
    nor02_2x L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix5 (.Y (
             L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_nx4), .A0 (FilterDin_3__1__0), .A1 (
             FilterDin_3__1__1)) ;
    aoi21 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix67 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_11), .A0 (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_nx328), .A1 (FilterDin_3__1__2), .B0 (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_nx8)) ;
    nor03_2x L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix9 (.Y (
             L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_nx8), .A0 (FilterDin_3__1__2), .A1 (
             FilterDin_3__1__0), .A2 (FilterDin_3__1__1)) ;
    xnor2 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix59 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_12), .A0 (
          FilterDin_3__1__3), .A1 (L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_nx8)) ;
    xnor2 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix51 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_13), .A0 (
          FilterDin_3__1__4), .A1 (L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_nx12)) ;
    nor04 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix13 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_nx12), .A0 (FilterDin_3__1__3), .A1 (
          FilterDin_3__1__2), .A2 (FilterDin_3__1__0), .A3 (FilterDin_3__1__1)
          ) ;
    xnor2 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix43 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_14), .A0 (
          FilterDin_3__1__5), .A1 (L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_nx16)) ;
    nor02ii L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix17 (.Y (
            L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_nx16), .A0 (FilterDin_3__1__4), .A1 (
            L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_nx12)) ;
    xnor2 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix35 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_15), .A0 (
          FilterDin_3__1__6), .A1 (L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_nx20)) ;
    nor02ii L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix21 (.Y (
            L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_nx20), .A0 (FilterDin_3__1__5), .A1 (
            L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_nx16)) ;
    xnor2 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix27 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_16), .A0 (
          FilterDin_3__1__7), .A1 (L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_nx24)) ;
    nor02ii L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix25 (.Y (
            L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_nx24), .A0 (FilterDin_3__1__6), .A1 (
            L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_nx20)) ;
    inv01 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix329 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_nx328), .A (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_nx4)) ;
    inv02 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix383 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_nx384), .A (
          L1_3_L2_1_G2_MINI_ALU_BoothP_0)) ;
    dff L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_0 (.Q (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_0), .QB (\$dummy [820]), 
        .D (L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .CLK (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    nor02_2x L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix567 (.Y (
             L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566), .A0 (RST), .A1 (
             L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644)) ;
    dff L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_1 (.Q (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_1), .QB (\$dummy [821]), 
        .D (L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .CLK (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_2 (.Q (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_2), .QB (\$dummy [822]), 
        .D (L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .CLK (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_3 (.Q (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_3), .QB (\$dummy [823]), 
        .D (L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .CLK (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_4 (.Q (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_4), .QB (\$dummy [824]), 
        .D (L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .CLK (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_5 (.Q (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_5), .QB (\$dummy [825]), 
        .D (L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .CLK (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_6 (.Q (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_6), .QB (\$dummy [826]), 
        .D (L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .CLK (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_7 (.Q (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_7), .QB (\$dummy [827]), 
        .D (L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .CLK (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_8 (.Q (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_8), .QB (\$dummy [828]), 
        .D (L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .CLK (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_9 (.Q (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_9), .QB (\$dummy [829]), 
        .D (L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .CLK (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_10 (.Q (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_10), .QB (\$dummy [830])
        , .D (L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .CLK (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_11 (.Q (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_11), .QB (\$dummy [831])
        , .D (L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .CLK (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_12 (.Q (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_12), .QB (\$dummy [832])
        , .D (L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .CLK (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_13 (.Q (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_13), .QB (\$dummy [833])
        , .D (L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .CLK (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_14 (.Q (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_14), .QB (\$dummy [834])
        , .D (L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .CLK (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_15 (.Q (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_15), .QB (\$dummy [835])
        , .D (L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .CLK (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_16 (.Q (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_16), .QB (\$dummy [836])
        , .D (L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .CLK (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    inv02 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix623 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624), .A (CLK)) ;
    inv02 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix625 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626), .A (CLK)) ;
    inv02 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix627 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628), .A (CLK)) ;
    inv02 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix643 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644), .A (nx8258)) ;
    dff L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_0 (.Q (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_0), .QB (\$dummy [837]), 
        .D (L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .CLK (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    nor02_2x L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix567 (.Y (
             L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566), .A0 (RST), .A1 (
             L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644)) ;
    dff L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_1 (.Q (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_1), .QB (\$dummy [838]), 
        .D (L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .CLK (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_2 (.Q (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_2), .QB (\$dummy [839]), 
        .D (L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .CLK (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_3 (.Q (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_3), .QB (\$dummy [840]), 
        .D (L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .CLK (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_4 (.Q (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_4), .QB (\$dummy [841]), 
        .D (L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .CLK (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_5 (.Q (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_5), .QB (\$dummy [842]), 
        .D (L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .CLK (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_6 (.Q (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_6), .QB (\$dummy [843]), 
        .D (L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .CLK (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_7 (.Q (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_7), .QB (\$dummy [844]), 
        .D (L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .CLK (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_8 (.Q (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_8), .QB (\$dummy [845]), 
        .D (L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .CLK (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_9 (.Q (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_9), .QB (\$dummy [846]), 
        .D (L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .CLK (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_10 (.Q (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_10), .QB (\$dummy [847])
        , .D (L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .CLK (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_11 (.Q (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_11), .QB (\$dummy [848])
        , .D (L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .CLK (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_12 (.Q (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_12), .QB (\$dummy [849])
        , .D (L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .CLK (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_13 (.Q (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_13), .QB (\$dummy [850])
        , .D (L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .CLK (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_14 (.Q (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_14), .QB (\$dummy [851])
        , .D (L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .CLK (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_15 (.Q (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_15), .QB (\$dummy [852])
        , .D (L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .CLK (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_16 (.Q (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_16), .QB (\$dummy [853])
        , .D (L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .CLK (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    inv02 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix623 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624), .A (CLK)) ;
    inv02 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix625 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626), .A (CLK)) ;
    inv02 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix627 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628), .A (CLK)) ;
    inv02 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix643 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644), .A (nx8264)) ;
    dff L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_0 (.Q (
        L1_3_L2_1_G2_MINI_ALU_BoothP_0), .QB (\$dummy [854]), .D (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .CLK (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    nor02_2x L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix567 (.Y (
             L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566), .A0 (RST), .A1 (
             L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    dff L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_1 (.Q (
        L1_3_L2_1_G2_MINI_ALU_BoothP_1), .QB (\$dummy [855]), .D (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .CLK (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_2 (.Q (
        L1_3_L2_1_G2_MINI_ALU_BoothP_2), .QB (\$dummy [856]), .D (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .CLK (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_3 (.Q (
        L1_3_L2_1_G2_MINI_ALU_BoothP_3), .QB (\$dummy [857]), .D (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .CLK (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_4 (.Q (
        L1_3_L2_1_G2_MINI_ALU_BoothP_4), .QB (\$dummy [858]), .D (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .CLK (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_5 (.Q (
        L1_3_L2_1_G2_MINI_ALU_BoothP_5), .QB (\$dummy [859]), .D (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .CLK (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_6 (.Q (
        L1_3_L2_1_G2_MINI_ALU_BoothP_6), .QB (\$dummy [860]), .D (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .CLK (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_7 (.Q (
        L1_3_L2_1_G2_MINI_ALU_BoothP_7), .QB (\$dummy [861]), .D (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .CLK (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_8 (.Q (
        L1_3_L2_1_G2_MINI_ALU_BoothP_8), .QB (\$dummy [862]), .D (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .CLK (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_9 (.Q (
        L1_3_L2_1_G2_MINI_ALU_BoothP_9), .QB (\$dummy [863]), .D (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .CLK (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_10 (.Q (
        L1_3_L2_1_G2_MINI_ALU_BoothP_10), .QB (\$dummy [864]), .D (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .CLK (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_11 (.Q (
        L1_3_L2_1_G2_MINI_ALU_BoothP_11), .QB (\$dummy [865]), .D (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .CLK (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_12 (.Q (
        L1_3_L2_1_G2_MINI_ALU_BoothP_12), .QB (\$dummy [866]), .D (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .CLK (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_13 (.Q (
        L1_3_L2_1_G2_MINI_ALU_BoothP_13), .QB (\$dummy [867]), .D (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .CLK (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_14 (.Q (
        L1_3_L2_1_G2_MINI_ALU_BoothP_14), .QB (\$dummy [868]), .D (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .CLK (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_15 (.Q (
        L1_3_L2_1_G2_MINI_ALU_BoothP_15), .QB (\$dummy [869]), .D (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .CLK (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_16 (.Q (
        L1_3_L2_1_G2_MINI_ALU_BoothP_16), .QB (\$dummy [870]), .D (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .CLK (
        L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    inv02 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix623 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624), .A (CLK)) ;
    inv02 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix625 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626), .A (CLK)) ;
    inv02 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix627 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628), .A (CLK)) ;
    inv02 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix643 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644), .A (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642)) ;
    xor2 L1_3_L2_2_G2_MINI_ALU_ix83 (.Y (L2Results_4__0), .A0 (L1Results_9__0), 
         .A1 (L1Results_8__0)) ;
    xnor2 L1_3_L2_2_G2_MINI_ALU_ix380 (.Y (L1_3_L2_2_G2_MINI_ALU_nx379), .A0 (
          L1_3_L2_2_G2_MINI_ALU_nx381), .A1 (L1_3_L2_2_G2_MINI_ALU_nx383)) ;
    nand02 L1_3_L2_2_G2_MINI_ALU_ix382 (.Y (L1_3_L2_2_G2_MINI_ALU_nx381), .A0 (
           L1_3_L2_2_G2_MINI_ALU_BoothOperand_0), .A1 (nx8284)) ;
    xnor2 L1_3_L2_2_G2_MINI_ALU_ix384 (.Y (L1_3_L2_2_G2_MINI_ALU_nx383), .A0 (
          L1_3_L2_2_G2_MINI_ALU_BoothOperand_1), .A1 (
          L1_3_L2_2_G2_MINI_ALU_BoothP_1)) ;
    inv01 L1_3_L2_2_G2_MINI_ALU_ix388 (.Y (L1_3_L2_2_G2_MINI_ALU_nx387), .A (
          L1_3_L2_2_G2_MINI_ALU_BoothP_2)) ;
    xnor2 L1_3_L2_2_G2_MINI_ALU_ix390 (.Y (L1_3_L2_2_G2_MINI_ALU_nx389), .A0 (
          L1_3_L2_2_G2_MINI_ALU_nx391), .A1 (L1_3_L2_2_G2_MINI_ALU_nx395)) ;
    aoi32 L1_3_L2_2_G2_MINI_ALU_ix392 (.Y (L1_3_L2_2_G2_MINI_ALU_nx391), .A0 (
          L1_3_L2_2_G2_MINI_ALU_BoothOperand_0), .A1 (nx8284), .A2 (
          L1_3_L2_2_G2_MINI_ALU_nx154), .B0 (L1_3_L2_2_G2_MINI_ALU_BoothP_1), .B1 (
          L1_3_L2_2_G2_MINI_ALU_BoothOperand_1)) ;
    xnor2 L1_3_L2_2_G2_MINI_ALU_ix396 (.Y (L1_3_L2_2_G2_MINI_ALU_nx395), .A0 (
          L1_3_L2_2_G2_MINI_ALU_BoothOperand_2), .A1 (
          L1_3_L2_2_G2_MINI_ALU_BoothP_2)) ;
    inv01 L1_3_L2_2_G2_MINI_ALU_ix400 (.Y (L1_3_L2_2_G2_MINI_ALU_nx399), .A (
          L1_3_L2_2_G2_MINI_ALU_BoothP_3)) ;
    xnor2 L1_3_L2_2_G2_MINI_ALU_ix402 (.Y (L1_3_L2_2_G2_MINI_ALU_nx401), .A0 (
          L1_3_L2_2_G2_MINI_ALU_nx403), .A1 (L1_3_L2_2_G2_MINI_ALU_nx405)) ;
    xnor2 L1_3_L2_2_G2_MINI_ALU_ix406 (.Y (L1_3_L2_2_G2_MINI_ALU_nx405), .A0 (
          L1_3_L2_2_G2_MINI_ALU_BoothOperand_3), .A1 (
          L1_3_L2_2_G2_MINI_ALU_BoothP_3)) ;
    inv01 L1_3_L2_2_G2_MINI_ALU_ix410 (.Y (L1_3_L2_2_G2_MINI_ALU_nx409), .A (
          L1_3_L2_2_G2_MINI_ALU_BoothP_4)) ;
    xnor2 L1_3_L2_2_G2_MINI_ALU_ix412 (.Y (L1_3_L2_2_G2_MINI_ALU_nx411), .A0 (
          L1_3_L2_2_G2_MINI_ALU_nx413), .A1 (L1_3_L2_2_G2_MINI_ALU_nx415)) ;
    xnor2 L1_3_L2_2_G2_MINI_ALU_ix416 (.Y (L1_3_L2_2_G2_MINI_ALU_nx415), .A0 (
          L1_3_L2_2_G2_MINI_ALU_BoothOperand_4), .A1 (
          L1_3_L2_2_G2_MINI_ALU_BoothP_4)) ;
    inv01 L1_3_L2_2_G2_MINI_ALU_ix420 (.Y (L1_3_L2_2_G2_MINI_ALU_nx419), .A (
          L1_3_L2_2_G2_MINI_ALU_BoothP_5)) ;
    xnor2 L1_3_L2_2_G2_MINI_ALU_ix422 (.Y (L1_3_L2_2_G2_MINI_ALU_nx421), .A0 (
          L1_3_L2_2_G2_MINI_ALU_nx423), .A1 (L1_3_L2_2_G2_MINI_ALU_nx425)) ;
    xnor2 L1_3_L2_2_G2_MINI_ALU_ix426 (.Y (L1_3_L2_2_G2_MINI_ALU_nx425), .A0 (
          L1_3_L2_2_G2_MINI_ALU_BoothOperand_5), .A1 (
          L1_3_L2_2_G2_MINI_ALU_BoothP_5)) ;
    inv01 L1_3_L2_2_G2_MINI_ALU_ix430 (.Y (L1_3_L2_2_G2_MINI_ALU_nx429), .A (
          L1_3_L2_2_G2_MINI_ALU_BoothP_6)) ;
    xnor2 L1_3_L2_2_G2_MINI_ALU_ix432 (.Y (L1_3_L2_2_G2_MINI_ALU_nx431), .A0 (
          L1_3_L2_2_G2_MINI_ALU_nx433), .A1 (L1_3_L2_2_G2_MINI_ALU_nx435)) ;
    xnor2 L1_3_L2_2_G2_MINI_ALU_ix436 (.Y (L1_3_L2_2_G2_MINI_ALU_nx435), .A0 (
          L1_3_L2_2_G2_MINI_ALU_BoothOperand_6), .A1 (
          L1_3_L2_2_G2_MINI_ALU_BoothP_6)) ;
    inv01 L1_3_L2_2_G2_MINI_ALU_ix440 (.Y (L1_3_L2_2_G2_MINI_ALU_nx439), .A (
          L1_3_L2_2_G2_MINI_ALU_BoothP_7)) ;
    xnor2 L1_3_L2_2_G2_MINI_ALU_ix442 (.Y (L1_3_L2_2_G2_MINI_ALU_nx441), .A0 (
          L1_3_L2_2_G2_MINI_ALU_nx443), .A1 (L1_3_L2_2_G2_MINI_ALU_nx445)) ;
    xnor2 L1_3_L2_2_G2_MINI_ALU_ix446 (.Y (L1_3_L2_2_G2_MINI_ALU_nx445), .A0 (
          L1_3_L2_2_G2_MINI_ALU_BoothOperand_7), .A1 (
          L1_3_L2_2_G2_MINI_ALU_BoothP_7)) ;
    inv01 L1_3_L2_2_G2_MINI_ALU_ix450 (.Y (L1_3_L2_2_G2_MINI_ALU_nx449), .A (
          L1_3_L2_2_G2_MINI_ALU_BoothP_8)) ;
    xnor2 L1_3_L2_2_G2_MINI_ALU_ix452 (.Y (L1_3_L2_2_G2_MINI_ALU_nx451), .A0 (
          L1_3_L2_2_G2_MINI_ALU_nx453), .A1 (L1_3_L2_2_G2_MINI_ALU_nx455)) ;
    xnor2 L1_3_L2_2_G2_MINI_ALU_ix456 (.Y (L1_3_L2_2_G2_MINI_ALU_nx455), .A0 (
          L1_3_L2_2_G2_MINI_ALU_BoothOperand_8), .A1 (
          L1_3_L2_2_G2_MINI_ALU_BoothP_8)) ;
    xor2 L1_3_L2_2_G2_MINI_ALU_ix317 (.Y (L1_3_L2_2_G2_MINI_ALU_nx316), .A0 (
         L1_3_L2_2_G2_MINI_ALU_nx461), .A1 (L1_3_L2_2_G2_MINI_ALU_nx463)) ;
    xnor2 L1_3_L2_2_G2_MINI_ALU_ix464 (.Y (L1_3_L2_2_G2_MINI_ALU_nx463), .A0 (
          L1_3_L2_2_G2_MINI_ALU_BoothOperand_9), .A1 (
          L1_3_L2_2_G2_MINI_ALU_BoothP_9)) ;
    xor2 L1_3_L2_2_G2_MINI_ALU_ix337 (.Y (L1_3_L2_2_G2_MINI_ALU_nx336), .A0 (
         L1_3_L2_2_G2_MINI_ALU_nx467), .A1 (L1_3_L2_2_G2_MINI_ALU_nx471)) ;
    inv01 L1_3_L2_2_G2_MINI_ALU_ix470 (.Y (L1_3_L2_2_G2_MINI_ALU_nx469), .A (
          L1_3_L2_2_G2_MINI_ALU_BoothP_9)) ;
    xnor2 L1_3_L2_2_G2_MINI_ALU_ix472 (.Y (L1_3_L2_2_G2_MINI_ALU_nx471), .A0 (
          L1_3_L2_2_G2_MINI_ALU_BoothOperand_10), .A1 (
          L1_3_L2_2_G2_MINI_ALU_BoothP_10)) ;
    xor2 L1_3_L2_2_G2_MINI_ALU_ix357 (.Y (L1_3_L2_2_G2_MINI_ALU_nx356), .A0 (
         L1_3_L2_2_G2_MINI_ALU_nx475), .A1 (L1_3_L2_2_G2_MINI_ALU_nx479)) ;
    inv01 L1_3_L2_2_G2_MINI_ALU_ix478 (.Y (L1_3_L2_2_G2_MINI_ALU_nx477), .A (
          L1_3_L2_2_G2_MINI_ALU_BoothP_10)) ;
    xnor2 L1_3_L2_2_G2_MINI_ALU_ix480 (.Y (L1_3_L2_2_G2_MINI_ALU_nx479), .A0 (
          L1_3_L2_2_G2_MINI_ALU_BoothOperand_11), .A1 (
          L1_3_L2_2_G2_MINI_ALU_BoothP_11)) ;
    xor2 L1_3_L2_2_G2_MINI_ALU_ix377 (.Y (L1_3_L2_2_G2_MINI_ALU_nx376), .A0 (
         L1_3_L2_2_G2_MINI_ALU_nx483), .A1 (L1_3_L2_2_G2_MINI_ALU_nx487)) ;
    inv01 L1_3_L2_2_G2_MINI_ALU_ix486 (.Y (L1_3_L2_2_G2_MINI_ALU_nx485), .A (
          L1_3_L2_2_G2_MINI_ALU_BoothP_11)) ;
    xnor2 L1_3_L2_2_G2_MINI_ALU_ix488 (.Y (L1_3_L2_2_G2_MINI_ALU_nx487), .A0 (
          L1_3_L2_2_G2_MINI_ALU_BoothOperand_12), .A1 (
          L1_3_L2_2_G2_MINI_ALU_BoothP_12)) ;
    xor2 L1_3_L2_2_G2_MINI_ALU_ix397 (.Y (L1_3_L2_2_G2_MINI_ALU_nx396), .A0 (
         L1_3_L2_2_G2_MINI_ALU_nx491), .A1 (L1_3_L2_2_G2_MINI_ALU_nx495)) ;
    inv01 L1_3_L2_2_G2_MINI_ALU_ix494 (.Y (L1_3_L2_2_G2_MINI_ALU_nx493), .A (
          L1_3_L2_2_G2_MINI_ALU_BoothP_12)) ;
    xnor2 L1_3_L2_2_G2_MINI_ALU_ix496 (.Y (L1_3_L2_2_G2_MINI_ALU_nx495), .A0 (
          L1_3_L2_2_G2_MINI_ALU_BoothOperand_13), .A1 (
          L1_3_L2_2_G2_MINI_ALU_BoothP_13)) ;
    xor2 L1_3_L2_2_G2_MINI_ALU_ix417 (.Y (L1_3_L2_2_G2_MINI_ALU_nx416), .A0 (
         L1_3_L2_2_G2_MINI_ALU_nx499), .A1 (L1_3_L2_2_G2_MINI_ALU_nx503)) ;
    inv01 L1_3_L2_2_G2_MINI_ALU_ix502 (.Y (L1_3_L2_2_G2_MINI_ALU_nx501), .A (
          L1_3_L2_2_G2_MINI_ALU_BoothP_13)) ;
    xnor2 L1_3_L2_2_G2_MINI_ALU_ix504 (.Y (L1_3_L2_2_G2_MINI_ALU_nx503), .A0 (
          L1_3_L2_2_G2_MINI_ALU_BoothOperand_14), .A1 (
          L1_3_L2_2_G2_MINI_ALU_BoothP_14)) ;
    xor2 L1_3_L2_2_G2_MINI_ALU_ix437 (.Y (L1_3_L2_2_G2_MINI_ALU_nx436), .A0 (
         L1_3_L2_2_G2_MINI_ALU_nx507), .A1 (L1_3_L2_2_G2_MINI_ALU_nx511)) ;
    inv01 L1_3_L2_2_G2_MINI_ALU_ix510 (.Y (L1_3_L2_2_G2_MINI_ALU_nx509), .A (
          L1_3_L2_2_G2_MINI_ALU_BoothP_14)) ;
    xnor2 L1_3_L2_2_G2_MINI_ALU_ix512 (.Y (L1_3_L2_2_G2_MINI_ALU_nx511), .A0 (
          L1_3_L2_2_G2_MINI_ALU_BoothOperand_15), .A1 (
          L1_3_L2_2_G2_MINI_ALU_BoothP_15)) ;
    xnor2 L1_3_L2_2_G2_MINI_ALU_ix457 (.Y (L1_3_L2_2_G2_MINI_ALU_nx456), .A0 (
          L1_3_L2_2_G2_MINI_ALU_nx515), .A1 (L1_3_L2_2_G2_MINI_ALU_nx454)) ;
    inv01 L1_3_L2_2_G2_MINI_ALU_ix518 (.Y (L1_3_L2_2_G2_MINI_ALU_nx517), .A (
          L1_3_L2_2_G2_MINI_ALU_BoothP_15)) ;
    xor2 L1_3_L2_2_G2_MINI_ALU_ix455 (.Y (L1_3_L2_2_G2_MINI_ALU_nx454), .A0 (
         L1_3_L2_2_G2_MINI_ALU_BoothOperand_16), .A1 (
         L1_3_L2_2_G2_MINI_ALU_BoothP_16)) ;
    mux21_ni L1_3_L2_2_G2_MINI_ALU_ix91 (.Y (L1FirstOperands_8__0), .A0 (
             L1_3_L2_2_G2_MINI_ALU_BoothP_1), .A1 (WindowDin_3__2__0), .S0 (
             Instr)) ;
    mux21_ni L1_3_L2_2_G2_MINI_ALU_ix99 (.Y (L1FirstOperands_8__1), .A0 (
             L1_3_L2_2_G2_MINI_ALU_BoothP_2), .A1 (WindowDin_3__2__1), .S0 (
             Instr)) ;
    mux21_ni L1_3_L2_2_G2_MINI_ALU_ix107 (.Y (L1FirstOperands_8__2), .A0 (
             L1_3_L2_2_G2_MINI_ALU_BoothP_3), .A1 (WindowDin_3__2__2), .S0 (
             Instr)) ;
    mux21_ni L1_3_L2_2_G2_MINI_ALU_ix115 (.Y (L1FirstOperands_8__3), .A0 (
             L1_3_L2_2_G2_MINI_ALU_BoothP_4), .A1 (WindowDin_3__2__3), .S0 (
             Instr)) ;
    mux21_ni L1_3_L2_2_G2_MINI_ALU_ix123 (.Y (L1FirstOperands_8__4), .A0 (
             L1_3_L2_2_G2_MINI_ALU_BoothP_5), .A1 (WindowDin_3__2__4), .S0 (
             Instr)) ;
    mux21_ni L1_3_L2_2_G2_MINI_ALU_ix131 (.Y (L1FirstOperands_8__5), .A0 (
             L1_3_L2_2_G2_MINI_ALU_BoothP_6), .A1 (WindowDin_3__2__5), .S0 (
             Instr)) ;
    mux21_ni L1_3_L2_2_G2_MINI_ALU_ix139 (.Y (L1FirstOperands_8__6), .A0 (
             L1_3_L2_2_G2_MINI_ALU_BoothP_7), .A1 (WindowDin_3__2__6), .S0 (
             Instr)) ;
    mux21_ni L1_3_L2_2_G2_MINI_ALU_ix147 (.Y (L1FirstOperands_8__7), .A0 (
             L1_3_L2_2_G2_MINI_ALU_BoothP_8), .A1 (WindowDin_3__2__7), .S0 (
             Instr)) ;
    xor2 L1_3_L2_2_G2_MINI_ALU_ix77 (.Y (L2Results_4__1), .A0 (
         L1_3_L2_2_G2_MINI_ALU_nx529), .A1 (L1_3_L2_2_G2_MINI_ALU_nx531)) ;
    nand02 L1_3_L2_2_G2_MINI_ALU_ix530 (.Y (L1_3_L2_2_G2_MINI_ALU_nx529), .A0 (
           L1Results_9__0), .A1 (L1Results_8__0)) ;
    xnor2 L1_3_L2_2_G2_MINI_ALU_ix532 (.Y (L1_3_L2_2_G2_MINI_ALU_nx531), .A0 (
          L1Results_9__1), .A1 (L1Results_8__1)) ;
    xor2 L1_3_L2_2_G2_MINI_ALU_ix75 (.Y (L2Results_4__2), .A0 (
         L1_3_L2_2_G2_MINI_ALU_nx534), .A1 (L1_3_L2_2_G2_MINI_ALU_nx537)) ;
    aoi32 L1_3_L2_2_G2_MINI_ALU_ix535 (.Y (L1_3_L2_2_G2_MINI_ALU_nx534), .A0 (
          L1Results_9__0), .A1 (L1Results_8__0), .A2 (L1_3_L2_2_G2_MINI_ALU_nx30
          ), .B0 (L1Results_8__1), .B1 (L1Results_9__1)) ;
    xnor2 L1_3_L2_2_G2_MINI_ALU_ix538 (.Y (L1_3_L2_2_G2_MINI_ALU_nx537), .A0 (
          L1Results_9__2), .A1 (L1Results_8__2)) ;
    xor2 L1_3_L2_2_G2_MINI_ALU_ix73 (.Y (L2Results_4__3), .A0 (
         L1_3_L2_2_G2_MINI_ALU_nx540), .A1 (L1_3_L2_2_G2_MINI_ALU_nx544)) ;
    aoi22 L1_3_L2_2_G2_MINI_ALU_ix541 (.Y (L1_3_L2_2_G2_MINI_ALU_nx540), .A0 (
          L1Results_8__2), .A1 (L1Results_9__2), .B0 (L1_3_L2_2_G2_MINI_ALU_nx40
          ), .B1 (L1_3_L2_2_G2_MINI_ALU_nx24)) ;
    xnor2 L1_3_L2_2_G2_MINI_ALU_ix545 (.Y (L1_3_L2_2_G2_MINI_ALU_nx544), .A0 (
          L1Results_9__3), .A1 (L1Results_8__3)) ;
    xor2 L1_3_L2_2_G2_MINI_ALU_ix71 (.Y (L2Results_4__4), .A0 (
         L1_3_L2_2_G2_MINI_ALU_nx547), .A1 (L1_3_L2_2_G2_MINI_ALU_nx551)) ;
    aoi22 L1_3_L2_2_G2_MINI_ALU_ix548 (.Y (L1_3_L2_2_G2_MINI_ALU_nx547), .A0 (
          L1Results_8__3), .A1 (L1Results_9__3), .B0 (L1_3_L2_2_G2_MINI_ALU_nx44
          ), .B1 (L1_3_L2_2_G2_MINI_ALU_nx18)) ;
    xnor2 L1_3_L2_2_G2_MINI_ALU_ix552 (.Y (L1_3_L2_2_G2_MINI_ALU_nx551), .A0 (
          L1Results_9__4), .A1 (L1Results_8__4)) ;
    xor2 L1_3_L2_2_G2_MINI_ALU_ix69 (.Y (L2Results_4__5), .A0 (
         L1_3_L2_2_G2_MINI_ALU_nx554), .A1 (L1_3_L2_2_G2_MINI_ALU_nx558)) ;
    aoi22 L1_3_L2_2_G2_MINI_ALU_ix555 (.Y (L1_3_L2_2_G2_MINI_ALU_nx554), .A0 (
          L1Results_8__4), .A1 (L1Results_9__4), .B0 (L1_3_L2_2_G2_MINI_ALU_nx48
          ), .B1 (L1_3_L2_2_G2_MINI_ALU_nx12)) ;
    xnor2 L1_3_L2_2_G2_MINI_ALU_ix559 (.Y (L1_3_L2_2_G2_MINI_ALU_nx558), .A0 (
          L1Results_9__5), .A1 (L1Results_8__5)) ;
    xor2 L1_3_L2_2_G2_MINI_ALU_ix67 (.Y (L2Results_4__6), .A0 (
         L1_3_L2_2_G2_MINI_ALU_nx561), .A1 (L1_3_L2_2_G2_MINI_ALU_nx565)) ;
    aoi22 L1_3_L2_2_G2_MINI_ALU_ix562 (.Y (L1_3_L2_2_G2_MINI_ALU_nx561), .A0 (
          L1Results_8__5), .A1 (L1Results_9__5), .B0 (L1_3_L2_2_G2_MINI_ALU_nx52
          ), .B1 (L1_3_L2_2_G2_MINI_ALU_nx6)) ;
    xnor2 L1_3_L2_2_G2_MINI_ALU_ix566 (.Y (L1_3_L2_2_G2_MINI_ALU_nx565), .A0 (
          L1Results_9__6), .A1 (L1Results_8__6)) ;
    xnor2 L1_3_L2_2_G2_MINI_ALU_ix65 (.Y (L2Results_4__7), .A0 (
          L1_3_L2_2_G2_MINI_ALU_nx568), .A1 (L1_3_L2_2_G2_MINI_ALU_nx62)) ;
    aoi22 L1_3_L2_2_G2_MINI_ALU_ix569 (.Y (L1_3_L2_2_G2_MINI_ALU_nx568), .A0 (
          L1Results_8__6), .A1 (L1Results_9__6), .B0 (L1_3_L2_2_G2_MINI_ALU_nx56
          ), .B1 (L1_3_L2_2_G2_MINI_ALU_nx0)) ;
    xor2 L1_3_L2_2_G2_MINI_ALU_ix63 (.Y (L1_3_L2_2_G2_MINI_ALU_nx62), .A0 (
         L1Results_9__7), .A1 (L1Results_8__7)) ;
    inv01 L1_3_L2_2_G2_MINI_ALU_ix155 (.Y (L1_3_L2_2_G2_MINI_ALU_nx154), .A (
          L1_3_L2_2_G2_MINI_ALU_nx383)) ;
    inv01 L1_3_L2_2_G2_MINI_ALU_ix57 (.Y (L1_3_L2_2_G2_MINI_ALU_nx56), .A (
          L1_3_L2_2_G2_MINI_ALU_nx561)) ;
    inv01 L1_3_L2_2_G2_MINI_ALU_ix53 (.Y (L1_3_L2_2_G2_MINI_ALU_nx52), .A (
          L1_3_L2_2_G2_MINI_ALU_nx554)) ;
    inv01 L1_3_L2_2_G2_MINI_ALU_ix49 (.Y (L1_3_L2_2_G2_MINI_ALU_nx48), .A (
          L1_3_L2_2_G2_MINI_ALU_nx547)) ;
    inv01 L1_3_L2_2_G2_MINI_ALU_ix45 (.Y (L1_3_L2_2_G2_MINI_ALU_nx44), .A (
          L1_3_L2_2_G2_MINI_ALU_nx540)) ;
    inv01 L1_3_L2_2_G2_MINI_ALU_ix41 (.Y (L1_3_L2_2_G2_MINI_ALU_nx40), .A (
          L1_3_L2_2_G2_MINI_ALU_nx534)) ;
    inv01 L1_3_L2_2_G2_MINI_ALU_ix31 (.Y (L1_3_L2_2_G2_MINI_ALU_nx30), .A (
          L1_3_L2_2_G2_MINI_ALU_nx531)) ;
    inv01 L1_3_L2_2_G2_MINI_ALU_ix25 (.Y (L1_3_L2_2_G2_MINI_ALU_nx24), .A (
          L1_3_L2_2_G2_MINI_ALU_nx537)) ;
    inv01 L1_3_L2_2_G2_MINI_ALU_ix19 (.Y (L1_3_L2_2_G2_MINI_ALU_nx18), .A (
          L1_3_L2_2_G2_MINI_ALU_nx544)) ;
    inv01 L1_3_L2_2_G2_MINI_ALU_ix13 (.Y (L1_3_L2_2_G2_MINI_ALU_nx12), .A (
          L1_3_L2_2_G2_MINI_ALU_nx551)) ;
    inv01 L1_3_L2_2_G2_MINI_ALU_ix7 (.Y (L1_3_L2_2_G2_MINI_ALU_nx6), .A (
          L1_3_L2_2_G2_MINI_ALU_nx558)) ;
    inv01 L1_3_L2_2_G2_MINI_ALU_ix1 (.Y (L1_3_L2_2_G2_MINI_ALU_nx0), .A (
          L1_3_L2_2_G2_MINI_ALU_nx565)) ;
    fake_gnd L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix216 (.Y (
             L1_3_L2_2_G2_MINI_ALU_WindowCellShiftedLeft_16)) ;
    nor02ii L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix81 (.Y (
            L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_nx80), .A0 (Instr), .A1 (Start)) ;
    aoi21 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix77 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_10), .A0 (
          FilterDin_3__2__1), .A1 (FilterDin_3__2__0), .B0 (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_nx4)) ;
    nor02_2x L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix5 (.Y (
             L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_nx4), .A0 (FilterDin_3__2__0), .A1 (
             FilterDin_3__2__1)) ;
    aoi21 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix67 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_11), .A0 (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_nx328), .A1 (FilterDin_3__2__2), .B0 (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_nx8)) ;
    nor03_2x L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix9 (.Y (
             L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_nx8), .A0 (FilterDin_3__2__2), .A1 (
             FilterDin_3__2__0), .A2 (FilterDin_3__2__1)) ;
    xnor2 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix59 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_12), .A0 (
          FilterDin_3__2__3), .A1 (L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_nx8)) ;
    xnor2 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix51 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_13), .A0 (
          FilterDin_3__2__4), .A1 (L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_nx12)) ;
    nor04 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix13 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_nx12), .A0 (FilterDin_3__2__3), .A1 (
          FilterDin_3__2__2), .A2 (FilterDin_3__2__0), .A3 (FilterDin_3__2__1)
          ) ;
    xnor2 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix43 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_14), .A0 (
          FilterDin_3__2__5), .A1 (L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_nx16)) ;
    nor02ii L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix17 (.Y (
            L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_nx16), .A0 (FilterDin_3__2__4), .A1 (
            L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_nx12)) ;
    xnor2 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix35 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_15), .A0 (
          FilterDin_3__2__6), .A1 (L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_nx20)) ;
    nor02ii L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix21 (.Y (
            L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_nx20), .A0 (FilterDin_3__2__5), .A1 (
            L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_nx16)) ;
    xnor2 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix27 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_16), .A0 (
          FilterDin_3__2__7), .A1 (L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_nx24)) ;
    nor02ii L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix25 (.Y (
            L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_nx24), .A0 (FilterDin_3__2__6), .A1 (
            L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_nx20)) ;
    inv01 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix329 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_nx328), .A (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_nx4)) ;
    inv02 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix383 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_nx384), .A (
          L1_3_L2_2_G2_MINI_ALU_BoothP_0)) ;
    dff L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_0 (.Q (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_0), .QB (\$dummy [871]), 
        .D (L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .CLK (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    nor02_2x L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix567 (.Y (
             L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566), .A0 (RST), .A1 (
             L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644)) ;
    dff L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_1 (.Q (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_1), .QB (\$dummy [872]), 
        .D (L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .CLK (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_2 (.Q (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_2), .QB (\$dummy [873]), 
        .D (L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .CLK (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_3 (.Q (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_3), .QB (\$dummy [874]), 
        .D (L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .CLK (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_4 (.Q (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_4), .QB (\$dummy [875]), 
        .D (L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .CLK (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_5 (.Q (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_5), .QB (\$dummy [876]), 
        .D (L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .CLK (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_6 (.Q (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_6), .QB (\$dummy [877]), 
        .D (L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .CLK (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_7 (.Q (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_7), .QB (\$dummy [878]), 
        .D (L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .CLK (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_8 (.Q (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_8), .QB (\$dummy [879]), 
        .D (L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .CLK (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_9 (.Q (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_9), .QB (\$dummy [880]), 
        .D (L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .CLK (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_10 (.Q (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_10), .QB (\$dummy [881])
        , .D (L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .CLK (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_11 (.Q (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_11), .QB (\$dummy [882])
        , .D (L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .CLK (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_12 (.Q (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_12), .QB (\$dummy [883])
        , .D (L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .CLK (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_13 (.Q (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_13), .QB (\$dummy [884])
        , .D (L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .CLK (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_14 (.Q (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_14), .QB (\$dummy [885])
        , .D (L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .CLK (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_15 (.Q (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_15), .QB (\$dummy [886])
        , .D (L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .CLK (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_16 (.Q (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_16), .QB (\$dummy [887])
        , .D (L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .CLK (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    inv02 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix623 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624), .A (CLK)) ;
    inv02 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix625 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626), .A (CLK)) ;
    inv02 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix627 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628), .A (CLK)) ;
    inv02 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix643 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644), .A (nx8298)) ;
    dff L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_0 (.Q (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_0), .QB (\$dummy [888]), 
        .D (L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .CLK (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    nor02_2x L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix567 (.Y (
             L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566), .A0 (RST), .A1 (
             L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644)) ;
    dff L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_1 (.Q (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_1), .QB (\$dummy [889]), 
        .D (L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .CLK (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_2 (.Q (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_2), .QB (\$dummy [890]), 
        .D (L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .CLK (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_3 (.Q (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_3), .QB (\$dummy [891]), 
        .D (L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .CLK (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_4 (.Q (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_4), .QB (\$dummy [892]), 
        .D (L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .CLK (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_5 (.Q (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_5), .QB (\$dummy [893]), 
        .D (L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .CLK (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_6 (.Q (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_6), .QB (\$dummy [894]), 
        .D (L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .CLK (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_7 (.Q (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_7), .QB (\$dummy [895]), 
        .D (L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .CLK (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_8 (.Q (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_8), .QB (\$dummy [896]), 
        .D (L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .CLK (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_9 (.Q (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_9), .QB (\$dummy [897]), 
        .D (L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .CLK (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_10 (.Q (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_10), .QB (\$dummy [898])
        , .D (L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .CLK (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_11 (.Q (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_11), .QB (\$dummy [899])
        , .D (L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .CLK (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_12 (.Q (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_12), .QB (\$dummy [900])
        , .D (L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .CLK (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_13 (.Q (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_13), .QB (\$dummy [901])
        , .D (L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .CLK (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_14 (.Q (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_14), .QB (\$dummy [902])
        , .D (L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .CLK (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_15 (.Q (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_15), .QB (\$dummy [903])
        , .D (L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .CLK (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_16 (.Q (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_16), .QB (\$dummy [904])
        , .D (L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .CLK (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    inv02 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix623 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624), .A (CLK)) ;
    inv02 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix625 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626), .A (CLK)) ;
    inv02 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix627 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628), .A (CLK)) ;
    inv02 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix643 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644), .A (nx8304)) ;
    dff L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_0 (.Q (
        L1_3_L2_2_G2_MINI_ALU_BoothP_0), .QB (\$dummy [905]), .D (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .CLK (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    nor02_2x L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix567 (.Y (
             L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566), .A0 (RST), .A1 (
             L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    dff L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_1 (.Q (
        L1_3_L2_2_G2_MINI_ALU_BoothP_1), .QB (\$dummy [906]), .D (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .CLK (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_2 (.Q (
        L1_3_L2_2_G2_MINI_ALU_BoothP_2), .QB (\$dummy [907]), .D (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .CLK (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_3 (.Q (
        L1_3_L2_2_G2_MINI_ALU_BoothP_3), .QB (\$dummy [908]), .D (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .CLK (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_4 (.Q (
        L1_3_L2_2_G2_MINI_ALU_BoothP_4), .QB (\$dummy [909]), .D (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .CLK (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_5 (.Q (
        L1_3_L2_2_G2_MINI_ALU_BoothP_5), .QB (\$dummy [910]), .D (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .CLK (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_6 (.Q (
        L1_3_L2_2_G2_MINI_ALU_BoothP_6), .QB (\$dummy [911]), .D (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .CLK (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_7 (.Q (
        L1_3_L2_2_G2_MINI_ALU_BoothP_7), .QB (\$dummy [912]), .D (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .CLK (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_8 (.Q (
        L1_3_L2_2_G2_MINI_ALU_BoothP_8), .QB (\$dummy [913]), .D (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .CLK (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_9 (.Q (
        L1_3_L2_2_G2_MINI_ALU_BoothP_9), .QB (\$dummy [914]), .D (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .CLK (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_10 (.Q (
        L1_3_L2_2_G2_MINI_ALU_BoothP_10), .QB (\$dummy [915]), .D (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .CLK (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_11 (.Q (
        L1_3_L2_2_G2_MINI_ALU_BoothP_11), .QB (\$dummy [916]), .D (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .CLK (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_12 (.Q (
        L1_3_L2_2_G2_MINI_ALU_BoothP_12), .QB (\$dummy [917]), .D (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .CLK (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_13 (.Q (
        L1_3_L2_2_G2_MINI_ALU_BoothP_13), .QB (\$dummy [918]), .D (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .CLK (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_14 (.Q (
        L1_3_L2_2_G2_MINI_ALU_BoothP_14), .QB (\$dummy [919]), .D (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .CLK (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_15 (.Q (
        L1_3_L2_2_G2_MINI_ALU_BoothP_15), .QB (\$dummy [920]), .D (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .CLK (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_16 (.Q (
        L1_3_L2_2_G2_MINI_ALU_BoothP_16), .QB (\$dummy [921]), .D (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .CLK (
        L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    inv02 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix623 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624), .A (CLK)) ;
    inv02 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix625 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626), .A (CLK)) ;
    inv02 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix627 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628), .A (CLK)) ;
    inv02 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix643 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644), .A (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642)) ;
    xor2 L1_3_L2_3_G2_MINI_ALU_ix83 (.Y (L2Results_5__0), .A0 (L1Results_11__0)
         , .A1 (L1Results_10__0)) ;
    xnor2 L1_3_L2_3_G2_MINI_ALU_ix380 (.Y (L1_3_L2_3_G2_MINI_ALU_nx379), .A0 (
          L1_3_L2_3_G2_MINI_ALU_nx381), .A1 (L1_3_L2_3_G2_MINI_ALU_nx383)) ;
    nand02 L1_3_L2_3_G2_MINI_ALU_ix382 (.Y (L1_3_L2_3_G2_MINI_ALU_nx381), .A0 (
           L1_3_L2_3_G2_MINI_ALU_BoothOperand_0), .A1 (nx8324)) ;
    xnor2 L1_3_L2_3_G2_MINI_ALU_ix384 (.Y (L1_3_L2_3_G2_MINI_ALU_nx383), .A0 (
          L1_3_L2_3_G2_MINI_ALU_BoothOperand_1), .A1 (
          L1_3_L2_3_G2_MINI_ALU_BoothP_1)) ;
    inv01 L1_3_L2_3_G2_MINI_ALU_ix388 (.Y (L1_3_L2_3_G2_MINI_ALU_nx387), .A (
          L1_3_L2_3_G2_MINI_ALU_BoothP_2)) ;
    xnor2 L1_3_L2_3_G2_MINI_ALU_ix390 (.Y (L1_3_L2_3_G2_MINI_ALU_nx389), .A0 (
          L1_3_L2_3_G2_MINI_ALU_nx391), .A1 (L1_3_L2_3_G2_MINI_ALU_nx395)) ;
    aoi32 L1_3_L2_3_G2_MINI_ALU_ix392 (.Y (L1_3_L2_3_G2_MINI_ALU_nx391), .A0 (
          L1_3_L2_3_G2_MINI_ALU_BoothOperand_0), .A1 (nx8324), .A2 (
          L1_3_L2_3_G2_MINI_ALU_nx154), .B0 (L1_3_L2_3_G2_MINI_ALU_BoothP_1), .B1 (
          L1_3_L2_3_G2_MINI_ALU_BoothOperand_1)) ;
    xnor2 L1_3_L2_3_G2_MINI_ALU_ix396 (.Y (L1_3_L2_3_G2_MINI_ALU_nx395), .A0 (
          L1_3_L2_3_G2_MINI_ALU_BoothOperand_2), .A1 (
          L1_3_L2_3_G2_MINI_ALU_BoothP_2)) ;
    inv01 L1_3_L2_3_G2_MINI_ALU_ix400 (.Y (L1_3_L2_3_G2_MINI_ALU_nx399), .A (
          L1_3_L2_3_G2_MINI_ALU_BoothP_3)) ;
    xnor2 L1_3_L2_3_G2_MINI_ALU_ix402 (.Y (L1_3_L2_3_G2_MINI_ALU_nx401), .A0 (
          L1_3_L2_3_G2_MINI_ALU_nx403), .A1 (L1_3_L2_3_G2_MINI_ALU_nx405)) ;
    xnor2 L1_3_L2_3_G2_MINI_ALU_ix406 (.Y (L1_3_L2_3_G2_MINI_ALU_nx405), .A0 (
          L1_3_L2_3_G2_MINI_ALU_BoothOperand_3), .A1 (
          L1_3_L2_3_G2_MINI_ALU_BoothP_3)) ;
    inv01 L1_3_L2_3_G2_MINI_ALU_ix410 (.Y (L1_3_L2_3_G2_MINI_ALU_nx409), .A (
          L1_3_L2_3_G2_MINI_ALU_BoothP_4)) ;
    xnor2 L1_3_L2_3_G2_MINI_ALU_ix412 (.Y (L1_3_L2_3_G2_MINI_ALU_nx411), .A0 (
          L1_3_L2_3_G2_MINI_ALU_nx413), .A1 (L1_3_L2_3_G2_MINI_ALU_nx415)) ;
    xnor2 L1_3_L2_3_G2_MINI_ALU_ix416 (.Y (L1_3_L2_3_G2_MINI_ALU_nx415), .A0 (
          L1_3_L2_3_G2_MINI_ALU_BoothOperand_4), .A1 (
          L1_3_L2_3_G2_MINI_ALU_BoothP_4)) ;
    inv01 L1_3_L2_3_G2_MINI_ALU_ix420 (.Y (L1_3_L2_3_G2_MINI_ALU_nx419), .A (
          L1_3_L2_3_G2_MINI_ALU_BoothP_5)) ;
    xnor2 L1_3_L2_3_G2_MINI_ALU_ix422 (.Y (L1_3_L2_3_G2_MINI_ALU_nx421), .A0 (
          L1_3_L2_3_G2_MINI_ALU_nx423), .A1 (L1_3_L2_3_G2_MINI_ALU_nx425)) ;
    xnor2 L1_3_L2_3_G2_MINI_ALU_ix426 (.Y (L1_3_L2_3_G2_MINI_ALU_nx425), .A0 (
          L1_3_L2_3_G2_MINI_ALU_BoothOperand_5), .A1 (
          L1_3_L2_3_G2_MINI_ALU_BoothP_5)) ;
    inv01 L1_3_L2_3_G2_MINI_ALU_ix430 (.Y (L1_3_L2_3_G2_MINI_ALU_nx429), .A (
          L1_3_L2_3_G2_MINI_ALU_BoothP_6)) ;
    xnor2 L1_3_L2_3_G2_MINI_ALU_ix432 (.Y (L1_3_L2_3_G2_MINI_ALU_nx431), .A0 (
          L1_3_L2_3_G2_MINI_ALU_nx433), .A1 (L1_3_L2_3_G2_MINI_ALU_nx435)) ;
    xnor2 L1_3_L2_3_G2_MINI_ALU_ix436 (.Y (L1_3_L2_3_G2_MINI_ALU_nx435), .A0 (
          L1_3_L2_3_G2_MINI_ALU_BoothOperand_6), .A1 (
          L1_3_L2_3_G2_MINI_ALU_BoothP_6)) ;
    inv01 L1_3_L2_3_G2_MINI_ALU_ix440 (.Y (L1_3_L2_3_G2_MINI_ALU_nx439), .A (
          L1_3_L2_3_G2_MINI_ALU_BoothP_7)) ;
    xnor2 L1_3_L2_3_G2_MINI_ALU_ix442 (.Y (L1_3_L2_3_G2_MINI_ALU_nx441), .A0 (
          L1_3_L2_3_G2_MINI_ALU_nx443), .A1 (L1_3_L2_3_G2_MINI_ALU_nx445)) ;
    xnor2 L1_3_L2_3_G2_MINI_ALU_ix446 (.Y (L1_3_L2_3_G2_MINI_ALU_nx445), .A0 (
          L1_3_L2_3_G2_MINI_ALU_BoothOperand_7), .A1 (
          L1_3_L2_3_G2_MINI_ALU_BoothP_7)) ;
    inv01 L1_3_L2_3_G2_MINI_ALU_ix450 (.Y (L1_3_L2_3_G2_MINI_ALU_nx449), .A (
          L1_3_L2_3_G2_MINI_ALU_BoothP_8)) ;
    xnor2 L1_3_L2_3_G2_MINI_ALU_ix452 (.Y (L1_3_L2_3_G2_MINI_ALU_nx451), .A0 (
          L1_3_L2_3_G2_MINI_ALU_nx453), .A1 (L1_3_L2_3_G2_MINI_ALU_nx455)) ;
    xnor2 L1_3_L2_3_G2_MINI_ALU_ix456 (.Y (L1_3_L2_3_G2_MINI_ALU_nx455), .A0 (
          L1_3_L2_3_G2_MINI_ALU_BoothOperand_8), .A1 (
          L1_3_L2_3_G2_MINI_ALU_BoothP_8)) ;
    xor2 L1_3_L2_3_G2_MINI_ALU_ix317 (.Y (L1_3_L2_3_G2_MINI_ALU_nx316), .A0 (
         L1_3_L2_3_G2_MINI_ALU_nx461), .A1 (L1_3_L2_3_G2_MINI_ALU_nx463)) ;
    xnor2 L1_3_L2_3_G2_MINI_ALU_ix464 (.Y (L1_3_L2_3_G2_MINI_ALU_nx463), .A0 (
          L1_3_L2_3_G2_MINI_ALU_BoothOperand_9), .A1 (
          L1_3_L2_3_G2_MINI_ALU_BoothP_9)) ;
    xor2 L1_3_L2_3_G2_MINI_ALU_ix337 (.Y (L1_3_L2_3_G2_MINI_ALU_nx336), .A0 (
         L1_3_L2_3_G2_MINI_ALU_nx467), .A1 (L1_3_L2_3_G2_MINI_ALU_nx471)) ;
    inv01 L1_3_L2_3_G2_MINI_ALU_ix470 (.Y (L1_3_L2_3_G2_MINI_ALU_nx469), .A (
          L1_3_L2_3_G2_MINI_ALU_BoothP_9)) ;
    xnor2 L1_3_L2_3_G2_MINI_ALU_ix472 (.Y (L1_3_L2_3_G2_MINI_ALU_nx471), .A0 (
          L1_3_L2_3_G2_MINI_ALU_BoothOperand_10), .A1 (
          L1_3_L2_3_G2_MINI_ALU_BoothP_10)) ;
    xor2 L1_3_L2_3_G2_MINI_ALU_ix357 (.Y (L1_3_L2_3_G2_MINI_ALU_nx356), .A0 (
         L1_3_L2_3_G2_MINI_ALU_nx475), .A1 (L1_3_L2_3_G2_MINI_ALU_nx479)) ;
    inv01 L1_3_L2_3_G2_MINI_ALU_ix478 (.Y (L1_3_L2_3_G2_MINI_ALU_nx477), .A (
          L1_3_L2_3_G2_MINI_ALU_BoothP_10)) ;
    xnor2 L1_3_L2_3_G2_MINI_ALU_ix480 (.Y (L1_3_L2_3_G2_MINI_ALU_nx479), .A0 (
          L1_3_L2_3_G2_MINI_ALU_BoothOperand_11), .A1 (
          L1_3_L2_3_G2_MINI_ALU_BoothP_11)) ;
    xor2 L1_3_L2_3_G2_MINI_ALU_ix377 (.Y (L1_3_L2_3_G2_MINI_ALU_nx376), .A0 (
         L1_3_L2_3_G2_MINI_ALU_nx483), .A1 (L1_3_L2_3_G2_MINI_ALU_nx487)) ;
    inv01 L1_3_L2_3_G2_MINI_ALU_ix486 (.Y (L1_3_L2_3_G2_MINI_ALU_nx485), .A (
          L1_3_L2_3_G2_MINI_ALU_BoothP_11)) ;
    xnor2 L1_3_L2_3_G2_MINI_ALU_ix488 (.Y (L1_3_L2_3_G2_MINI_ALU_nx487), .A0 (
          L1_3_L2_3_G2_MINI_ALU_BoothOperand_12), .A1 (
          L1_3_L2_3_G2_MINI_ALU_BoothP_12)) ;
    xor2 L1_3_L2_3_G2_MINI_ALU_ix397 (.Y (L1_3_L2_3_G2_MINI_ALU_nx396), .A0 (
         L1_3_L2_3_G2_MINI_ALU_nx491), .A1 (L1_3_L2_3_G2_MINI_ALU_nx495)) ;
    inv01 L1_3_L2_3_G2_MINI_ALU_ix494 (.Y (L1_3_L2_3_G2_MINI_ALU_nx493), .A (
          L1_3_L2_3_G2_MINI_ALU_BoothP_12)) ;
    xnor2 L1_3_L2_3_G2_MINI_ALU_ix496 (.Y (L1_3_L2_3_G2_MINI_ALU_nx495), .A0 (
          L1_3_L2_3_G2_MINI_ALU_BoothOperand_13), .A1 (
          L1_3_L2_3_G2_MINI_ALU_BoothP_13)) ;
    xor2 L1_3_L2_3_G2_MINI_ALU_ix417 (.Y (L1_3_L2_3_G2_MINI_ALU_nx416), .A0 (
         L1_3_L2_3_G2_MINI_ALU_nx499), .A1 (L1_3_L2_3_G2_MINI_ALU_nx503)) ;
    inv01 L1_3_L2_3_G2_MINI_ALU_ix502 (.Y (L1_3_L2_3_G2_MINI_ALU_nx501), .A (
          L1_3_L2_3_G2_MINI_ALU_BoothP_13)) ;
    xnor2 L1_3_L2_3_G2_MINI_ALU_ix504 (.Y (L1_3_L2_3_G2_MINI_ALU_nx503), .A0 (
          L1_3_L2_3_G2_MINI_ALU_BoothOperand_14), .A1 (
          L1_3_L2_3_G2_MINI_ALU_BoothP_14)) ;
    xor2 L1_3_L2_3_G2_MINI_ALU_ix437 (.Y (L1_3_L2_3_G2_MINI_ALU_nx436), .A0 (
         L1_3_L2_3_G2_MINI_ALU_nx507), .A1 (L1_3_L2_3_G2_MINI_ALU_nx511)) ;
    inv01 L1_3_L2_3_G2_MINI_ALU_ix510 (.Y (L1_3_L2_3_G2_MINI_ALU_nx509), .A (
          L1_3_L2_3_G2_MINI_ALU_BoothP_14)) ;
    xnor2 L1_3_L2_3_G2_MINI_ALU_ix512 (.Y (L1_3_L2_3_G2_MINI_ALU_nx511), .A0 (
          L1_3_L2_3_G2_MINI_ALU_BoothOperand_15), .A1 (
          L1_3_L2_3_G2_MINI_ALU_BoothP_15)) ;
    xnor2 L1_3_L2_3_G2_MINI_ALU_ix457 (.Y (L1_3_L2_3_G2_MINI_ALU_nx456), .A0 (
          L1_3_L2_3_G2_MINI_ALU_nx515), .A1 (L1_3_L2_3_G2_MINI_ALU_nx454)) ;
    inv01 L1_3_L2_3_G2_MINI_ALU_ix518 (.Y (L1_3_L2_3_G2_MINI_ALU_nx517), .A (
          L1_3_L2_3_G2_MINI_ALU_BoothP_15)) ;
    xor2 L1_3_L2_3_G2_MINI_ALU_ix455 (.Y (L1_3_L2_3_G2_MINI_ALU_nx454), .A0 (
         L1_3_L2_3_G2_MINI_ALU_BoothOperand_16), .A1 (
         L1_3_L2_3_G2_MINI_ALU_BoothP_16)) ;
    mux21_ni L1_3_L2_3_G2_MINI_ALU_ix91 (.Y (L1FirstOperands_10__0), .A0 (
             L1_3_L2_3_G2_MINI_ALU_BoothP_1), .A1 (WindowDin_3__3__0), .S0 (
             Instr)) ;
    mux21_ni L1_3_L2_3_G2_MINI_ALU_ix99 (.Y (L1FirstOperands_10__1), .A0 (
             L1_3_L2_3_G2_MINI_ALU_BoothP_2), .A1 (WindowDin_3__3__1), .S0 (
             Instr)) ;
    mux21_ni L1_3_L2_3_G2_MINI_ALU_ix107 (.Y (L1FirstOperands_10__2), .A0 (
             L1_3_L2_3_G2_MINI_ALU_BoothP_3), .A1 (WindowDin_3__3__2), .S0 (
             Instr)) ;
    mux21_ni L1_3_L2_3_G2_MINI_ALU_ix115 (.Y (L1FirstOperands_10__3), .A0 (
             L1_3_L2_3_G2_MINI_ALU_BoothP_4), .A1 (WindowDin_3__3__3), .S0 (
             Instr)) ;
    mux21_ni L1_3_L2_3_G2_MINI_ALU_ix123 (.Y (L1FirstOperands_10__4), .A0 (
             L1_3_L2_3_G2_MINI_ALU_BoothP_5), .A1 (WindowDin_3__3__4), .S0 (
             Instr)) ;
    mux21_ni L1_3_L2_3_G2_MINI_ALU_ix131 (.Y (L1FirstOperands_10__5), .A0 (
             L1_3_L2_3_G2_MINI_ALU_BoothP_6), .A1 (WindowDin_3__3__5), .S0 (
             Instr)) ;
    mux21_ni L1_3_L2_3_G2_MINI_ALU_ix139 (.Y (L1FirstOperands_10__6), .A0 (
             L1_3_L2_3_G2_MINI_ALU_BoothP_7), .A1 (WindowDin_3__3__6), .S0 (
             Instr)) ;
    mux21_ni L1_3_L2_3_G2_MINI_ALU_ix147 (.Y (L1FirstOperands_10__7), .A0 (
             L1_3_L2_3_G2_MINI_ALU_BoothP_8), .A1 (WindowDin_3__3__7), .S0 (
             Instr)) ;
    xor2 L1_3_L2_3_G2_MINI_ALU_ix77 (.Y (L2Results_5__1), .A0 (
         L1_3_L2_3_G2_MINI_ALU_nx529), .A1 (L1_3_L2_3_G2_MINI_ALU_nx531)) ;
    nand02 L1_3_L2_3_G2_MINI_ALU_ix530 (.Y (L1_3_L2_3_G2_MINI_ALU_nx529), .A0 (
           L1Results_11__0), .A1 (L1Results_10__0)) ;
    xnor2 L1_3_L2_3_G2_MINI_ALU_ix532 (.Y (L1_3_L2_3_G2_MINI_ALU_nx531), .A0 (
          L1Results_11__1), .A1 (L1Results_10__1)) ;
    xor2 L1_3_L2_3_G2_MINI_ALU_ix75 (.Y (L2Results_5__2), .A0 (
         L1_3_L2_3_G2_MINI_ALU_nx534), .A1 (L1_3_L2_3_G2_MINI_ALU_nx537)) ;
    aoi32 L1_3_L2_3_G2_MINI_ALU_ix535 (.Y (L1_3_L2_3_G2_MINI_ALU_nx534), .A0 (
          L1Results_11__0), .A1 (L1Results_10__0), .A2 (
          L1_3_L2_3_G2_MINI_ALU_nx30), .B0 (L1Results_10__1), .B1 (
          L1Results_11__1)) ;
    xnor2 L1_3_L2_3_G2_MINI_ALU_ix538 (.Y (L1_3_L2_3_G2_MINI_ALU_nx537), .A0 (
          L1Results_11__2), .A1 (L1Results_10__2)) ;
    xor2 L1_3_L2_3_G2_MINI_ALU_ix73 (.Y (L2Results_5__3), .A0 (
         L1_3_L2_3_G2_MINI_ALU_nx540), .A1 (L1_3_L2_3_G2_MINI_ALU_nx544)) ;
    aoi22 L1_3_L2_3_G2_MINI_ALU_ix541 (.Y (L1_3_L2_3_G2_MINI_ALU_nx540), .A0 (
          L1Results_10__2), .A1 (L1Results_11__2), .B0 (
          L1_3_L2_3_G2_MINI_ALU_nx40), .B1 (L1_3_L2_3_G2_MINI_ALU_nx24)) ;
    xnor2 L1_3_L2_3_G2_MINI_ALU_ix545 (.Y (L1_3_L2_3_G2_MINI_ALU_nx544), .A0 (
          L1Results_11__3), .A1 (L1Results_10__3)) ;
    xor2 L1_3_L2_3_G2_MINI_ALU_ix71 (.Y (L2Results_5__4), .A0 (
         L1_3_L2_3_G2_MINI_ALU_nx547), .A1 (L1_3_L2_3_G2_MINI_ALU_nx551)) ;
    aoi22 L1_3_L2_3_G2_MINI_ALU_ix548 (.Y (L1_3_L2_3_G2_MINI_ALU_nx547), .A0 (
          L1Results_10__3), .A1 (L1Results_11__3), .B0 (
          L1_3_L2_3_G2_MINI_ALU_nx44), .B1 (L1_3_L2_3_G2_MINI_ALU_nx18)) ;
    xnor2 L1_3_L2_3_G2_MINI_ALU_ix552 (.Y (L1_3_L2_3_G2_MINI_ALU_nx551), .A0 (
          L1Results_11__4), .A1 (L1Results_10__4)) ;
    xor2 L1_3_L2_3_G2_MINI_ALU_ix69 (.Y (L2Results_5__5), .A0 (
         L1_3_L2_3_G2_MINI_ALU_nx554), .A1 (L1_3_L2_3_G2_MINI_ALU_nx558)) ;
    aoi22 L1_3_L2_3_G2_MINI_ALU_ix555 (.Y (L1_3_L2_3_G2_MINI_ALU_nx554), .A0 (
          L1Results_10__4), .A1 (L1Results_11__4), .B0 (
          L1_3_L2_3_G2_MINI_ALU_nx48), .B1 (L1_3_L2_3_G2_MINI_ALU_nx12)) ;
    xnor2 L1_3_L2_3_G2_MINI_ALU_ix559 (.Y (L1_3_L2_3_G2_MINI_ALU_nx558), .A0 (
          L1Results_11__5), .A1 (L1Results_10__5)) ;
    xor2 L1_3_L2_3_G2_MINI_ALU_ix67 (.Y (L2Results_5__6), .A0 (
         L1_3_L2_3_G2_MINI_ALU_nx561), .A1 (L1_3_L2_3_G2_MINI_ALU_nx565)) ;
    aoi22 L1_3_L2_3_G2_MINI_ALU_ix562 (.Y (L1_3_L2_3_G2_MINI_ALU_nx561), .A0 (
          L1Results_10__5), .A1 (L1Results_11__5), .B0 (
          L1_3_L2_3_G2_MINI_ALU_nx52), .B1 (L1_3_L2_3_G2_MINI_ALU_nx6)) ;
    xnor2 L1_3_L2_3_G2_MINI_ALU_ix566 (.Y (L1_3_L2_3_G2_MINI_ALU_nx565), .A0 (
          L1Results_11__6), .A1 (L1Results_10__6)) ;
    xnor2 L1_3_L2_3_G2_MINI_ALU_ix65 (.Y (L2Results_5__7), .A0 (
          L1_3_L2_3_G2_MINI_ALU_nx568), .A1 (L1_3_L2_3_G2_MINI_ALU_nx62)) ;
    aoi22 L1_3_L2_3_G2_MINI_ALU_ix569 (.Y (L1_3_L2_3_G2_MINI_ALU_nx568), .A0 (
          L1Results_10__6), .A1 (L1Results_11__6), .B0 (
          L1_3_L2_3_G2_MINI_ALU_nx56), .B1 (L1_3_L2_3_G2_MINI_ALU_nx0)) ;
    xor2 L1_3_L2_3_G2_MINI_ALU_ix63 (.Y (L1_3_L2_3_G2_MINI_ALU_nx62), .A0 (
         L1Results_11__7), .A1 (L1Results_10__7)) ;
    inv01 L1_3_L2_3_G2_MINI_ALU_ix155 (.Y (L1_3_L2_3_G2_MINI_ALU_nx154), .A (
          L1_3_L2_3_G2_MINI_ALU_nx383)) ;
    inv01 L1_3_L2_3_G2_MINI_ALU_ix57 (.Y (L1_3_L2_3_G2_MINI_ALU_nx56), .A (
          L1_3_L2_3_G2_MINI_ALU_nx561)) ;
    inv01 L1_3_L2_3_G2_MINI_ALU_ix53 (.Y (L1_3_L2_3_G2_MINI_ALU_nx52), .A (
          L1_3_L2_3_G2_MINI_ALU_nx554)) ;
    inv01 L1_3_L2_3_G2_MINI_ALU_ix49 (.Y (L1_3_L2_3_G2_MINI_ALU_nx48), .A (
          L1_3_L2_3_G2_MINI_ALU_nx547)) ;
    inv01 L1_3_L2_3_G2_MINI_ALU_ix45 (.Y (L1_3_L2_3_G2_MINI_ALU_nx44), .A (
          L1_3_L2_3_G2_MINI_ALU_nx540)) ;
    inv01 L1_3_L2_3_G2_MINI_ALU_ix41 (.Y (L1_3_L2_3_G2_MINI_ALU_nx40), .A (
          L1_3_L2_3_G2_MINI_ALU_nx534)) ;
    inv01 L1_3_L2_3_G2_MINI_ALU_ix31 (.Y (L1_3_L2_3_G2_MINI_ALU_nx30), .A (
          L1_3_L2_3_G2_MINI_ALU_nx531)) ;
    inv01 L1_3_L2_3_G2_MINI_ALU_ix25 (.Y (L1_3_L2_3_G2_MINI_ALU_nx24), .A (
          L1_3_L2_3_G2_MINI_ALU_nx537)) ;
    inv01 L1_3_L2_3_G2_MINI_ALU_ix19 (.Y (L1_3_L2_3_G2_MINI_ALU_nx18), .A (
          L1_3_L2_3_G2_MINI_ALU_nx544)) ;
    inv01 L1_3_L2_3_G2_MINI_ALU_ix13 (.Y (L1_3_L2_3_G2_MINI_ALU_nx12), .A (
          L1_3_L2_3_G2_MINI_ALU_nx551)) ;
    inv01 L1_3_L2_3_G2_MINI_ALU_ix7 (.Y (L1_3_L2_3_G2_MINI_ALU_nx6), .A (
          L1_3_L2_3_G2_MINI_ALU_nx558)) ;
    inv01 L1_3_L2_3_G2_MINI_ALU_ix1 (.Y (L1_3_L2_3_G2_MINI_ALU_nx0), .A (
          L1_3_L2_3_G2_MINI_ALU_nx565)) ;
    fake_gnd L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix216 (.Y (
             L1_3_L2_3_G2_MINI_ALU_WindowCellShiftedLeft_16)) ;
    nor02ii L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix81 (.Y (
            L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx80), .A0 (Instr), .A1 (Start)) ;
    aoi21 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix77 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_10), .A0 (
          FilterDin_3__3__1), .A1 (FilterDin_3__3__0), .B0 (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx4)) ;
    nor02_2x L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix5 (.Y (
             L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx4), .A0 (FilterDin_3__3__0), .A1 (
             FilterDin_3__3__1)) ;
    aoi21 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix67 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_11), .A0 (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx328), .A1 (FilterDin_3__3__2), .B0 (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx8)) ;
    nor03_2x L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix9 (.Y (
             L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx8), .A0 (FilterDin_3__3__2), .A1 (
             FilterDin_3__3__0), .A2 (FilterDin_3__3__1)) ;
    xnor2 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix59 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_12), .A0 (
          FilterDin_3__3__3), .A1 (L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx8)) ;
    xnor2 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix51 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_13), .A0 (
          FilterDin_3__3__4), .A1 (L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx12)) ;
    nor04 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix13 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx12), .A0 (FilterDin_3__3__3), .A1 (
          FilterDin_3__3__2), .A2 (FilterDin_3__3__0), .A3 (FilterDin_3__3__1)
          ) ;
    xnor2 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix43 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_14), .A0 (
          FilterDin_3__3__5), .A1 (L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx16)) ;
    nor02ii L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix17 (.Y (
            L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx16), .A0 (FilterDin_3__3__4), .A1 (
            L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx12)) ;
    xnor2 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix35 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_15), .A0 (
          FilterDin_3__3__6), .A1 (L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx20)) ;
    nor02ii L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix21 (.Y (
            L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx20), .A0 (FilterDin_3__3__5), .A1 (
            L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx16)) ;
    xnor2 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix27 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_16), .A0 (
          FilterDin_3__3__7), .A1 (L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx24)) ;
    nor02ii L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix25 (.Y (
            L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx24), .A0 (FilterDin_3__3__6), .A1 (
            L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx20)) ;
    inv01 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix329 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx328), .A (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx4)) ;
    inv02 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix383 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx384), .A (
          L1_3_L2_3_G2_MINI_ALU_BoothP_0)) ;
    dff L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_0 (.Q (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_0), .QB (\$dummy [922]), 
        .D (L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .CLK (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    nor02_2x L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix567 (.Y (
             L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566), .A0 (RST), .A1 (
             L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644)) ;
    dff L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_1 (.Q (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_1), .QB (\$dummy [923]), 
        .D (L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .CLK (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_2 (.Q (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_2), .QB (\$dummy [924]), 
        .D (L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .CLK (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_3 (.Q (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_3), .QB (\$dummy [925]), 
        .D (L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .CLK (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_4 (.Q (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_4), .QB (\$dummy [926]), 
        .D (L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .CLK (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_5 (.Q (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_5), .QB (\$dummy [927]), 
        .D (L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .CLK (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_6 (.Q (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_6), .QB (\$dummy [928]), 
        .D (L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .CLK (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_7 (.Q (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_7), .QB (\$dummy [929]), 
        .D (L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .CLK (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_8 (.Q (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_8), .QB (\$dummy [930]), 
        .D (L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .CLK (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_9 (.Q (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_9), .QB (\$dummy [931]), 
        .D (L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .CLK (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_10 (.Q (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_10), .QB (\$dummy [932])
        , .D (L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .CLK (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_11 (.Q (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_11), .QB (\$dummy [933])
        , .D (L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .CLK (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_12 (.Q (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_12), .QB (\$dummy [934])
        , .D (L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .CLK (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_13 (.Q (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_13), .QB (\$dummy [935])
        , .D (L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .CLK (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_14 (.Q (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_14), .QB (\$dummy [936])
        , .D (L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .CLK (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_15 (.Q (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_15), .QB (\$dummy [937])
        , .D (L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .CLK (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_16 (.Q (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_16), .QB (\$dummy [938])
        , .D (L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .CLK (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    inv02 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix623 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624), .A (CLK)) ;
    inv02 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix625 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626), .A (CLK)) ;
    inv02 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix627 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628), .A (CLK)) ;
    inv02 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix643 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644), .A (nx8338)) ;
    dff L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_0 (.Q (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_0), .QB (\$dummy [939]), 
        .D (L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .CLK (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    nor02_2x L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix567 (.Y (
             L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566), .A0 (RST), .A1 (
             L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644)) ;
    dff L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_1 (.Q (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_1), .QB (\$dummy [940]), 
        .D (L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .CLK (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_2 (.Q (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_2), .QB (\$dummy [941]), 
        .D (L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .CLK (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_3 (.Q (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_3), .QB (\$dummy [942]), 
        .D (L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .CLK (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_4 (.Q (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_4), .QB (\$dummy [943]), 
        .D (L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .CLK (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_5 (.Q (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_5), .QB (\$dummy [944]), 
        .D (L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .CLK (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_6 (.Q (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_6), .QB (\$dummy [945]), 
        .D (L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .CLK (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_7 (.Q (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_7), .QB (\$dummy [946]), 
        .D (L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .CLK (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_8 (.Q (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_8), .QB (\$dummy [947]), 
        .D (L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .CLK (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_9 (.Q (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_9), .QB (\$dummy [948]), 
        .D (L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .CLK (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_10 (.Q (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_10), .QB (\$dummy [949])
        , .D (L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .CLK (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_11 (.Q (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_11), .QB (\$dummy [950])
        , .D (L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .CLK (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_12 (.Q (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_12), .QB (\$dummy [951])
        , .D (L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .CLK (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_13 (.Q (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_13), .QB (\$dummy [952])
        , .D (L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .CLK (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_14 (.Q (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_14), .QB (\$dummy [953])
        , .D (L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .CLK (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_15 (.Q (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_15), .QB (\$dummy [954])
        , .D (L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .CLK (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_16 (.Q (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_16), .QB (\$dummy [955])
        , .D (L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .CLK (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    inv02 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix623 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624), .A (CLK)) ;
    inv02 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix625 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626), .A (CLK)) ;
    inv02 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix627 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628), .A (CLK)) ;
    inv02 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix643 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644), .A (nx8344)) ;
    dff L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_0 (.Q (
        L1_3_L2_3_G2_MINI_ALU_BoothP_0), .QB (\$dummy [956]), .D (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .CLK (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    nor02_2x L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix567 (.Y (
             L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566), .A0 (RST), .A1 (
             L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    dff L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_1 (.Q (
        L1_3_L2_3_G2_MINI_ALU_BoothP_1), .QB (\$dummy [957]), .D (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .CLK (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_2 (.Q (
        L1_3_L2_3_G2_MINI_ALU_BoothP_2), .QB (\$dummy [958]), .D (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .CLK (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_3 (.Q (
        L1_3_L2_3_G2_MINI_ALU_BoothP_3), .QB (\$dummy [959]), .D (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .CLK (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_4 (.Q (
        L1_3_L2_3_G2_MINI_ALU_BoothP_4), .QB (\$dummy [960]), .D (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .CLK (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_5 (.Q (
        L1_3_L2_3_G2_MINI_ALU_BoothP_5), .QB (\$dummy [961]), .D (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .CLK (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_6 (.Q (
        L1_3_L2_3_G2_MINI_ALU_BoothP_6), .QB (\$dummy [962]), .D (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .CLK (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_7 (.Q (
        L1_3_L2_3_G2_MINI_ALU_BoothP_7), .QB (\$dummy [963]), .D (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .CLK (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_8 (.Q (
        L1_3_L2_3_G2_MINI_ALU_BoothP_8), .QB (\$dummy [964]), .D (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .CLK (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_9 (.Q (
        L1_3_L2_3_G2_MINI_ALU_BoothP_9), .QB (\$dummy [965]), .D (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .CLK (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_10 (.Q (
        L1_3_L2_3_G2_MINI_ALU_BoothP_10), .QB (\$dummy [966]), .D (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .CLK (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_11 (.Q (
        L1_3_L2_3_G2_MINI_ALU_BoothP_11), .QB (\$dummy [967]), .D (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .CLK (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_12 (.Q (
        L1_3_L2_3_G2_MINI_ALU_BoothP_12), .QB (\$dummy [968]), .D (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .CLK (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_13 (.Q (
        L1_3_L2_3_G2_MINI_ALU_BoothP_13), .QB (\$dummy [969]), .D (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .CLK (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_14 (.Q (
        L1_3_L2_3_G2_MINI_ALU_BoothP_14), .QB (\$dummy [970]), .D (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .CLK (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_15 (.Q (
        L1_3_L2_3_G2_MINI_ALU_BoothP_15), .QB (\$dummy [971]), .D (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .CLK (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_16 (.Q (
        L1_3_L2_3_G2_MINI_ALU_BoothP_16), .QB (\$dummy [972]), .D (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .CLK (
        L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    inv02 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix623 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624), .A (CLK)) ;
    inv02 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix625 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626), .A (CLK)) ;
    inv02 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix627 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628), .A (CLK)) ;
    inv02 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix643 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644), .A (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642)) ;
    xor2 L1_3_L2_4_G3_MINI_ALU_ix83 (.Y (L3Results_0__0), .A0 (L2Results_1__0), 
         .A1 (L2Results_0__0)) ;
    xnor2 L1_3_L2_4_G3_MINI_ALU_ix380 (.Y (L1_3_L2_4_G3_MINI_ALU_nx379), .A0 (
          L1_3_L2_4_G3_MINI_ALU_nx381), .A1 (L1_3_L2_4_G3_MINI_ALU_nx383)) ;
    nand02 L1_3_L2_4_G3_MINI_ALU_ix382 (.Y (L1_3_L2_4_G3_MINI_ALU_nx381), .A0 (
           L1_3_L2_4_G3_MINI_ALU_BoothOperand_0), .A1 (nx8364)) ;
    xnor2 L1_3_L2_4_G3_MINI_ALU_ix384 (.Y (L1_3_L2_4_G3_MINI_ALU_nx383), .A0 (
          L1_3_L2_4_G3_MINI_ALU_BoothOperand_1), .A1 (
          L1_3_L2_4_G3_MINI_ALU_BoothP_1)) ;
    inv01 L1_3_L2_4_G3_MINI_ALU_ix388 (.Y (L1_3_L2_4_G3_MINI_ALU_nx387), .A (
          L1_3_L2_4_G3_MINI_ALU_BoothP_2)) ;
    xnor2 L1_3_L2_4_G3_MINI_ALU_ix390 (.Y (L1_3_L2_4_G3_MINI_ALU_nx389), .A0 (
          L1_3_L2_4_G3_MINI_ALU_nx391), .A1 (L1_3_L2_4_G3_MINI_ALU_nx395)) ;
    aoi32 L1_3_L2_4_G3_MINI_ALU_ix392 (.Y (L1_3_L2_4_G3_MINI_ALU_nx391), .A0 (
          L1_3_L2_4_G3_MINI_ALU_BoothOperand_0), .A1 (nx8364), .A2 (
          L1_3_L2_4_G3_MINI_ALU_nx154), .B0 (L1_3_L2_4_G3_MINI_ALU_BoothP_1), .B1 (
          L1_3_L2_4_G3_MINI_ALU_BoothOperand_1)) ;
    xnor2 L1_3_L2_4_G3_MINI_ALU_ix396 (.Y (L1_3_L2_4_G3_MINI_ALU_nx395), .A0 (
          L1_3_L2_4_G3_MINI_ALU_BoothOperand_2), .A1 (
          L1_3_L2_4_G3_MINI_ALU_BoothP_2)) ;
    inv01 L1_3_L2_4_G3_MINI_ALU_ix400 (.Y (L1_3_L2_4_G3_MINI_ALU_nx399), .A (
          L1_3_L2_4_G3_MINI_ALU_BoothP_3)) ;
    xnor2 L1_3_L2_4_G3_MINI_ALU_ix402 (.Y (L1_3_L2_4_G3_MINI_ALU_nx401), .A0 (
          L1_3_L2_4_G3_MINI_ALU_nx403), .A1 (L1_3_L2_4_G3_MINI_ALU_nx405)) ;
    xnor2 L1_3_L2_4_G3_MINI_ALU_ix406 (.Y (L1_3_L2_4_G3_MINI_ALU_nx405), .A0 (
          L1_3_L2_4_G3_MINI_ALU_BoothOperand_3), .A1 (
          L1_3_L2_4_G3_MINI_ALU_BoothP_3)) ;
    inv01 L1_3_L2_4_G3_MINI_ALU_ix410 (.Y (L1_3_L2_4_G3_MINI_ALU_nx409), .A (
          L1_3_L2_4_G3_MINI_ALU_BoothP_4)) ;
    xnor2 L1_3_L2_4_G3_MINI_ALU_ix412 (.Y (L1_3_L2_4_G3_MINI_ALU_nx411), .A0 (
          L1_3_L2_4_G3_MINI_ALU_nx413), .A1 (L1_3_L2_4_G3_MINI_ALU_nx415)) ;
    xnor2 L1_3_L2_4_G3_MINI_ALU_ix416 (.Y (L1_3_L2_4_G3_MINI_ALU_nx415), .A0 (
          L1_3_L2_4_G3_MINI_ALU_BoothOperand_4), .A1 (
          L1_3_L2_4_G3_MINI_ALU_BoothP_4)) ;
    inv01 L1_3_L2_4_G3_MINI_ALU_ix420 (.Y (L1_3_L2_4_G3_MINI_ALU_nx419), .A (
          L1_3_L2_4_G3_MINI_ALU_BoothP_5)) ;
    xnor2 L1_3_L2_4_G3_MINI_ALU_ix422 (.Y (L1_3_L2_4_G3_MINI_ALU_nx421), .A0 (
          L1_3_L2_4_G3_MINI_ALU_nx423), .A1 (L1_3_L2_4_G3_MINI_ALU_nx425)) ;
    xnor2 L1_3_L2_4_G3_MINI_ALU_ix426 (.Y (L1_3_L2_4_G3_MINI_ALU_nx425), .A0 (
          L1_3_L2_4_G3_MINI_ALU_BoothOperand_5), .A1 (
          L1_3_L2_4_G3_MINI_ALU_BoothP_5)) ;
    inv01 L1_3_L2_4_G3_MINI_ALU_ix430 (.Y (L1_3_L2_4_G3_MINI_ALU_nx429), .A (
          L1_3_L2_4_G3_MINI_ALU_BoothP_6)) ;
    xnor2 L1_3_L2_4_G3_MINI_ALU_ix432 (.Y (L1_3_L2_4_G3_MINI_ALU_nx431), .A0 (
          L1_3_L2_4_G3_MINI_ALU_nx433), .A1 (L1_3_L2_4_G3_MINI_ALU_nx435)) ;
    xnor2 L1_3_L2_4_G3_MINI_ALU_ix436 (.Y (L1_3_L2_4_G3_MINI_ALU_nx435), .A0 (
          L1_3_L2_4_G3_MINI_ALU_BoothOperand_6), .A1 (
          L1_3_L2_4_G3_MINI_ALU_BoothP_6)) ;
    inv01 L1_3_L2_4_G3_MINI_ALU_ix440 (.Y (L1_3_L2_4_G3_MINI_ALU_nx439), .A (
          L1_3_L2_4_G3_MINI_ALU_BoothP_7)) ;
    xnor2 L1_3_L2_4_G3_MINI_ALU_ix442 (.Y (L1_3_L2_4_G3_MINI_ALU_nx441), .A0 (
          L1_3_L2_4_G3_MINI_ALU_nx443), .A1 (L1_3_L2_4_G3_MINI_ALU_nx445)) ;
    xnor2 L1_3_L2_4_G3_MINI_ALU_ix446 (.Y (L1_3_L2_4_G3_MINI_ALU_nx445), .A0 (
          L1_3_L2_4_G3_MINI_ALU_BoothOperand_7), .A1 (
          L1_3_L2_4_G3_MINI_ALU_BoothP_7)) ;
    inv01 L1_3_L2_4_G3_MINI_ALU_ix450 (.Y (L1_3_L2_4_G3_MINI_ALU_nx449), .A (
          L1_3_L2_4_G3_MINI_ALU_BoothP_8)) ;
    xnor2 L1_3_L2_4_G3_MINI_ALU_ix452 (.Y (L1_3_L2_4_G3_MINI_ALU_nx451), .A0 (
          L1_3_L2_4_G3_MINI_ALU_nx453), .A1 (L1_3_L2_4_G3_MINI_ALU_nx455)) ;
    xnor2 L1_3_L2_4_G3_MINI_ALU_ix456 (.Y (L1_3_L2_4_G3_MINI_ALU_nx455), .A0 (
          L1_3_L2_4_G3_MINI_ALU_BoothOperand_8), .A1 (
          L1_3_L2_4_G3_MINI_ALU_BoothP_8)) ;
    xor2 L1_3_L2_4_G3_MINI_ALU_ix317 (.Y (L1_3_L2_4_G3_MINI_ALU_nx316), .A0 (
         L1_3_L2_4_G3_MINI_ALU_nx461), .A1 (L1_3_L2_4_G3_MINI_ALU_nx463)) ;
    xnor2 L1_3_L2_4_G3_MINI_ALU_ix464 (.Y (L1_3_L2_4_G3_MINI_ALU_nx463), .A0 (
          L1_3_L2_4_G3_MINI_ALU_BoothOperand_9), .A1 (
          L1_3_L2_4_G3_MINI_ALU_BoothP_9)) ;
    xor2 L1_3_L2_4_G3_MINI_ALU_ix337 (.Y (L1_3_L2_4_G3_MINI_ALU_nx336), .A0 (
         L1_3_L2_4_G3_MINI_ALU_nx467), .A1 (L1_3_L2_4_G3_MINI_ALU_nx471)) ;
    inv01 L1_3_L2_4_G3_MINI_ALU_ix470 (.Y (L1_3_L2_4_G3_MINI_ALU_nx469), .A (
          L1_3_L2_4_G3_MINI_ALU_BoothP_9)) ;
    xnor2 L1_3_L2_4_G3_MINI_ALU_ix472 (.Y (L1_3_L2_4_G3_MINI_ALU_nx471), .A0 (
          L1_3_L2_4_G3_MINI_ALU_BoothOperand_10), .A1 (
          L1_3_L2_4_G3_MINI_ALU_BoothP_10)) ;
    xor2 L1_3_L2_4_G3_MINI_ALU_ix357 (.Y (L1_3_L2_4_G3_MINI_ALU_nx356), .A0 (
         L1_3_L2_4_G3_MINI_ALU_nx475), .A1 (L1_3_L2_4_G3_MINI_ALU_nx479)) ;
    inv01 L1_3_L2_4_G3_MINI_ALU_ix478 (.Y (L1_3_L2_4_G3_MINI_ALU_nx477), .A (
          L1_3_L2_4_G3_MINI_ALU_BoothP_10)) ;
    xnor2 L1_3_L2_4_G3_MINI_ALU_ix480 (.Y (L1_3_L2_4_G3_MINI_ALU_nx479), .A0 (
          L1_3_L2_4_G3_MINI_ALU_BoothOperand_11), .A1 (
          L1_3_L2_4_G3_MINI_ALU_BoothP_11)) ;
    xor2 L1_3_L2_4_G3_MINI_ALU_ix377 (.Y (L1_3_L2_4_G3_MINI_ALU_nx376), .A0 (
         L1_3_L2_4_G3_MINI_ALU_nx483), .A1 (L1_3_L2_4_G3_MINI_ALU_nx487)) ;
    inv01 L1_3_L2_4_G3_MINI_ALU_ix486 (.Y (L1_3_L2_4_G3_MINI_ALU_nx485), .A (
          L1_3_L2_4_G3_MINI_ALU_BoothP_11)) ;
    xnor2 L1_3_L2_4_G3_MINI_ALU_ix488 (.Y (L1_3_L2_4_G3_MINI_ALU_nx487), .A0 (
          L1_3_L2_4_G3_MINI_ALU_BoothOperand_12), .A1 (
          L1_3_L2_4_G3_MINI_ALU_BoothP_12)) ;
    xor2 L1_3_L2_4_G3_MINI_ALU_ix397 (.Y (L1_3_L2_4_G3_MINI_ALU_nx396), .A0 (
         L1_3_L2_4_G3_MINI_ALU_nx491), .A1 (L1_3_L2_4_G3_MINI_ALU_nx495)) ;
    inv01 L1_3_L2_4_G3_MINI_ALU_ix494 (.Y (L1_3_L2_4_G3_MINI_ALU_nx493), .A (
          L1_3_L2_4_G3_MINI_ALU_BoothP_12)) ;
    xnor2 L1_3_L2_4_G3_MINI_ALU_ix496 (.Y (L1_3_L2_4_G3_MINI_ALU_nx495), .A0 (
          L1_3_L2_4_G3_MINI_ALU_BoothOperand_13), .A1 (
          L1_3_L2_4_G3_MINI_ALU_BoothP_13)) ;
    xor2 L1_3_L2_4_G3_MINI_ALU_ix417 (.Y (L1_3_L2_4_G3_MINI_ALU_nx416), .A0 (
         L1_3_L2_4_G3_MINI_ALU_nx499), .A1 (L1_3_L2_4_G3_MINI_ALU_nx503)) ;
    inv01 L1_3_L2_4_G3_MINI_ALU_ix502 (.Y (L1_3_L2_4_G3_MINI_ALU_nx501), .A (
          L1_3_L2_4_G3_MINI_ALU_BoothP_13)) ;
    xnor2 L1_3_L2_4_G3_MINI_ALU_ix504 (.Y (L1_3_L2_4_G3_MINI_ALU_nx503), .A0 (
          L1_3_L2_4_G3_MINI_ALU_BoothOperand_14), .A1 (
          L1_3_L2_4_G3_MINI_ALU_BoothP_14)) ;
    xor2 L1_3_L2_4_G3_MINI_ALU_ix437 (.Y (L1_3_L2_4_G3_MINI_ALU_nx436), .A0 (
         L1_3_L2_4_G3_MINI_ALU_nx507), .A1 (L1_3_L2_4_G3_MINI_ALU_nx511)) ;
    inv01 L1_3_L2_4_G3_MINI_ALU_ix510 (.Y (L1_3_L2_4_G3_MINI_ALU_nx509), .A (
          L1_3_L2_4_G3_MINI_ALU_BoothP_14)) ;
    xnor2 L1_3_L2_4_G3_MINI_ALU_ix512 (.Y (L1_3_L2_4_G3_MINI_ALU_nx511), .A0 (
          L1_3_L2_4_G3_MINI_ALU_BoothOperand_15), .A1 (
          L1_3_L2_4_G3_MINI_ALU_BoothP_15)) ;
    xnor2 L1_3_L2_4_G3_MINI_ALU_ix457 (.Y (L1_3_L2_4_G3_MINI_ALU_nx456), .A0 (
          L1_3_L2_4_G3_MINI_ALU_nx515), .A1 (L1_3_L2_4_G3_MINI_ALU_nx454)) ;
    inv01 L1_3_L2_4_G3_MINI_ALU_ix518 (.Y (L1_3_L2_4_G3_MINI_ALU_nx517), .A (
          L1_3_L2_4_G3_MINI_ALU_BoothP_15)) ;
    xor2 L1_3_L2_4_G3_MINI_ALU_ix455 (.Y (L1_3_L2_4_G3_MINI_ALU_nx454), .A0 (
         L1_3_L2_4_G3_MINI_ALU_BoothOperand_16), .A1 (
         L1_3_L2_4_G3_MINI_ALU_BoothP_16)) ;
    mux21_ni L1_3_L2_4_G3_MINI_ALU_ix91 (.Y (L1FirstOperands_1__0), .A0 (
             L1_3_L2_4_G3_MINI_ALU_BoothP_1), .A1 (WindowDin_3__4__0), .S0 (
             Instr)) ;
    mux21_ni L1_3_L2_4_G3_MINI_ALU_ix99 (.Y (L1FirstOperands_1__1), .A0 (
             L1_3_L2_4_G3_MINI_ALU_BoothP_2), .A1 (WindowDin_3__4__1), .S0 (
             Instr)) ;
    mux21_ni L1_3_L2_4_G3_MINI_ALU_ix107 (.Y (L1FirstOperands_1__2), .A0 (
             L1_3_L2_4_G3_MINI_ALU_BoothP_3), .A1 (WindowDin_3__4__2), .S0 (
             Instr)) ;
    mux21_ni L1_3_L2_4_G3_MINI_ALU_ix115 (.Y (L1FirstOperands_1__3), .A0 (
             L1_3_L2_4_G3_MINI_ALU_BoothP_4), .A1 (WindowDin_3__4__3), .S0 (
             Instr)) ;
    mux21_ni L1_3_L2_4_G3_MINI_ALU_ix123 (.Y (L1FirstOperands_1__4), .A0 (
             L1_3_L2_4_G3_MINI_ALU_BoothP_5), .A1 (WindowDin_3__4__4), .S0 (
             Instr)) ;
    mux21_ni L1_3_L2_4_G3_MINI_ALU_ix131 (.Y (L1FirstOperands_1__5), .A0 (
             L1_3_L2_4_G3_MINI_ALU_BoothP_6), .A1 (WindowDin_3__4__5), .S0 (
             Instr)) ;
    mux21_ni L1_3_L2_4_G3_MINI_ALU_ix139 (.Y (L1FirstOperands_1__6), .A0 (
             L1_3_L2_4_G3_MINI_ALU_BoothP_7), .A1 (WindowDin_3__4__6), .S0 (
             Instr)) ;
    mux21_ni L1_3_L2_4_G3_MINI_ALU_ix147 (.Y (L1FirstOperands_1__7), .A0 (
             L1_3_L2_4_G3_MINI_ALU_BoothP_8), .A1 (WindowDin_3__4__7), .S0 (
             Instr)) ;
    xor2 L1_3_L2_4_G3_MINI_ALU_ix77 (.Y (L3Results_0__1), .A0 (
         L1_3_L2_4_G3_MINI_ALU_nx529), .A1 (L1_3_L2_4_G3_MINI_ALU_nx531)) ;
    nand02 L1_3_L2_4_G3_MINI_ALU_ix530 (.Y (L1_3_L2_4_G3_MINI_ALU_nx529), .A0 (
           L2Results_1__0), .A1 (L2Results_0__0)) ;
    xnor2 L1_3_L2_4_G3_MINI_ALU_ix532 (.Y (L1_3_L2_4_G3_MINI_ALU_nx531), .A0 (
          L2Results_1__1), .A1 (L2Results_0__1)) ;
    xor2 L1_3_L2_4_G3_MINI_ALU_ix75 (.Y (L3Results_0__2), .A0 (
         L1_3_L2_4_G3_MINI_ALU_nx534), .A1 (L1_3_L2_4_G3_MINI_ALU_nx537)) ;
    aoi32 L1_3_L2_4_G3_MINI_ALU_ix535 (.Y (L1_3_L2_4_G3_MINI_ALU_nx534), .A0 (
          L2Results_1__0), .A1 (L2Results_0__0), .A2 (L1_3_L2_4_G3_MINI_ALU_nx30
          ), .B0 (L2Results_0__1), .B1 (L2Results_1__1)) ;
    xnor2 L1_3_L2_4_G3_MINI_ALU_ix538 (.Y (L1_3_L2_4_G3_MINI_ALU_nx537), .A0 (
          L2Results_1__2), .A1 (L2Results_0__2)) ;
    xor2 L1_3_L2_4_G3_MINI_ALU_ix73 (.Y (L3Results_0__3), .A0 (
         L1_3_L2_4_G3_MINI_ALU_nx540), .A1 (L1_3_L2_4_G3_MINI_ALU_nx544)) ;
    aoi22 L1_3_L2_4_G3_MINI_ALU_ix541 (.Y (L1_3_L2_4_G3_MINI_ALU_nx540), .A0 (
          L2Results_0__2), .A1 (L2Results_1__2), .B0 (L1_3_L2_4_G3_MINI_ALU_nx40
          ), .B1 (L1_3_L2_4_G3_MINI_ALU_nx24)) ;
    xnor2 L1_3_L2_4_G3_MINI_ALU_ix545 (.Y (L1_3_L2_4_G3_MINI_ALU_nx544), .A0 (
          L2Results_1__3), .A1 (L2Results_0__3)) ;
    xor2 L1_3_L2_4_G3_MINI_ALU_ix71 (.Y (L3Results_0__4), .A0 (
         L1_3_L2_4_G3_MINI_ALU_nx547), .A1 (L1_3_L2_4_G3_MINI_ALU_nx551)) ;
    aoi22 L1_3_L2_4_G3_MINI_ALU_ix548 (.Y (L1_3_L2_4_G3_MINI_ALU_nx547), .A0 (
          L2Results_0__3), .A1 (L2Results_1__3), .B0 (L1_3_L2_4_G3_MINI_ALU_nx44
          ), .B1 (L1_3_L2_4_G3_MINI_ALU_nx18)) ;
    xnor2 L1_3_L2_4_G3_MINI_ALU_ix552 (.Y (L1_3_L2_4_G3_MINI_ALU_nx551), .A0 (
          L2Results_1__4), .A1 (L2Results_0__4)) ;
    xor2 L1_3_L2_4_G3_MINI_ALU_ix69 (.Y (L3Results_0__5), .A0 (
         L1_3_L2_4_G3_MINI_ALU_nx554), .A1 (L1_3_L2_4_G3_MINI_ALU_nx558)) ;
    aoi22 L1_3_L2_4_G3_MINI_ALU_ix555 (.Y (L1_3_L2_4_G3_MINI_ALU_nx554), .A0 (
          L2Results_0__4), .A1 (L2Results_1__4), .B0 (L1_3_L2_4_G3_MINI_ALU_nx48
          ), .B1 (L1_3_L2_4_G3_MINI_ALU_nx12)) ;
    xnor2 L1_3_L2_4_G3_MINI_ALU_ix559 (.Y (L1_3_L2_4_G3_MINI_ALU_nx558), .A0 (
          L2Results_1__5), .A1 (L2Results_0__5)) ;
    xor2 L1_3_L2_4_G3_MINI_ALU_ix67 (.Y (L3Results_0__6), .A0 (
         L1_3_L2_4_G3_MINI_ALU_nx561), .A1 (L1_3_L2_4_G3_MINI_ALU_nx565)) ;
    aoi22 L1_3_L2_4_G3_MINI_ALU_ix562 (.Y (L1_3_L2_4_G3_MINI_ALU_nx561), .A0 (
          L2Results_0__5), .A1 (L2Results_1__5), .B0 (L1_3_L2_4_G3_MINI_ALU_nx52
          ), .B1 (L1_3_L2_4_G3_MINI_ALU_nx6)) ;
    xnor2 L1_3_L2_4_G3_MINI_ALU_ix566 (.Y (L1_3_L2_4_G3_MINI_ALU_nx565), .A0 (
          L2Results_1__6), .A1 (L2Results_0__6)) ;
    xnor2 L1_3_L2_4_G3_MINI_ALU_ix65 (.Y (L3Results_0__7), .A0 (
          L1_3_L2_4_G3_MINI_ALU_nx568), .A1 (L1_3_L2_4_G3_MINI_ALU_nx62)) ;
    aoi22 L1_3_L2_4_G3_MINI_ALU_ix569 (.Y (L1_3_L2_4_G3_MINI_ALU_nx568), .A0 (
          L2Results_0__6), .A1 (L2Results_1__6), .B0 (L1_3_L2_4_G3_MINI_ALU_nx56
          ), .B1 (L1_3_L2_4_G3_MINI_ALU_nx0)) ;
    xor2 L1_3_L2_4_G3_MINI_ALU_ix63 (.Y (L1_3_L2_4_G3_MINI_ALU_nx62), .A0 (
         L2Results_1__7), .A1 (L2Results_0__7)) ;
    inv01 L1_3_L2_4_G3_MINI_ALU_ix155 (.Y (L1_3_L2_4_G3_MINI_ALU_nx154), .A (
          L1_3_L2_4_G3_MINI_ALU_nx383)) ;
    inv01 L1_3_L2_4_G3_MINI_ALU_ix57 (.Y (L1_3_L2_4_G3_MINI_ALU_nx56), .A (
          L1_3_L2_4_G3_MINI_ALU_nx561)) ;
    inv01 L1_3_L2_4_G3_MINI_ALU_ix53 (.Y (L1_3_L2_4_G3_MINI_ALU_nx52), .A (
          L1_3_L2_4_G3_MINI_ALU_nx554)) ;
    inv01 L1_3_L2_4_G3_MINI_ALU_ix49 (.Y (L1_3_L2_4_G3_MINI_ALU_nx48), .A (
          L1_3_L2_4_G3_MINI_ALU_nx547)) ;
    inv01 L1_3_L2_4_G3_MINI_ALU_ix45 (.Y (L1_3_L2_4_G3_MINI_ALU_nx44), .A (
          L1_3_L2_4_G3_MINI_ALU_nx540)) ;
    inv01 L1_3_L2_4_G3_MINI_ALU_ix41 (.Y (L1_3_L2_4_G3_MINI_ALU_nx40), .A (
          L1_3_L2_4_G3_MINI_ALU_nx534)) ;
    inv01 L1_3_L2_4_G3_MINI_ALU_ix31 (.Y (L1_3_L2_4_G3_MINI_ALU_nx30), .A (
          L1_3_L2_4_G3_MINI_ALU_nx531)) ;
    inv01 L1_3_L2_4_G3_MINI_ALU_ix25 (.Y (L1_3_L2_4_G3_MINI_ALU_nx24), .A (
          L1_3_L2_4_G3_MINI_ALU_nx537)) ;
    inv01 L1_3_L2_4_G3_MINI_ALU_ix19 (.Y (L1_3_L2_4_G3_MINI_ALU_nx18), .A (
          L1_3_L2_4_G3_MINI_ALU_nx544)) ;
    inv01 L1_3_L2_4_G3_MINI_ALU_ix13 (.Y (L1_3_L2_4_G3_MINI_ALU_nx12), .A (
          L1_3_L2_4_G3_MINI_ALU_nx551)) ;
    inv01 L1_3_L2_4_G3_MINI_ALU_ix7 (.Y (L1_3_L2_4_G3_MINI_ALU_nx6), .A (
          L1_3_L2_4_G3_MINI_ALU_nx558)) ;
    inv01 L1_3_L2_4_G3_MINI_ALU_ix1 (.Y (L1_3_L2_4_G3_MINI_ALU_nx0), .A (
          L1_3_L2_4_G3_MINI_ALU_nx565)) ;
    fake_gnd L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix216 (.Y (
             L1_3_L2_4_G3_MINI_ALU_WindowCellShiftedLeft_16)) ;
    nor02ii L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix81 (.Y (
            L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_nx80), .A0 (Instr), .A1 (Start)) ;
    aoi21 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix77 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_10), .A0 (
          FilterDin_3__4__1), .A1 (FilterDin_3__4__0), .B0 (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_nx4)) ;
    nor02_2x L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix5 (.Y (
             L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_nx4), .A0 (FilterDin_3__4__0), .A1 (
             FilterDin_3__4__1)) ;
    aoi21 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix67 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_11), .A0 (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_nx328), .A1 (FilterDin_3__4__2), .B0 (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_nx8)) ;
    nor03_2x L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix9 (.Y (
             L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_nx8), .A0 (FilterDin_3__4__2), .A1 (
             FilterDin_3__4__0), .A2 (FilterDin_3__4__1)) ;
    xnor2 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix59 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_12), .A0 (
          FilterDin_3__4__3), .A1 (L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_nx8)) ;
    xnor2 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix51 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_13), .A0 (
          FilterDin_3__4__4), .A1 (L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_nx12)) ;
    nor04 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix13 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_nx12), .A0 (FilterDin_3__4__3), .A1 (
          FilterDin_3__4__2), .A2 (FilterDin_3__4__0), .A3 (FilterDin_3__4__1)
          ) ;
    xnor2 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix43 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_14), .A0 (
          FilterDin_3__4__5), .A1 (L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_nx16)) ;
    nor02ii L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix17 (.Y (
            L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_nx16), .A0 (FilterDin_3__4__4), .A1 (
            L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_nx12)) ;
    xnor2 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix35 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_15), .A0 (
          FilterDin_3__4__6), .A1 (L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_nx20)) ;
    nor02ii L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix21 (.Y (
            L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_nx20), .A0 (FilterDin_3__4__5), .A1 (
            L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_nx16)) ;
    xnor2 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix27 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_16), .A0 (
          FilterDin_3__4__7), .A1 (L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_nx24)) ;
    nor02ii L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix25 (.Y (
            L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_nx24), .A0 (FilterDin_3__4__6), .A1 (
            L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_nx20)) ;
    inv01 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix329 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_nx328), .A (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_nx4)) ;
    inv02 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix383 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_nx384), .A (
          L1_3_L2_4_G3_MINI_ALU_BoothP_0)) ;
    dff L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_0 (.Q (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_0), .QB (\$dummy [973]), 
        .D (L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .CLK (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    nor02_2x L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix567 (.Y (
             L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566), .A0 (RST), .A1 (
             L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644)) ;
    dff L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_1 (.Q (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_1), .QB (\$dummy [974]), 
        .D (L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .CLK (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_2 (.Q (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_2), .QB (\$dummy [975]), 
        .D (L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .CLK (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_3 (.Q (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_3), .QB (\$dummy [976]), 
        .D (L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .CLK (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_4 (.Q (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_4), .QB (\$dummy [977]), 
        .D (L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .CLK (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_5 (.Q (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_5), .QB (\$dummy [978]), 
        .D (L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .CLK (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_6 (.Q (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_6), .QB (\$dummy [979]), 
        .D (L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .CLK (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_7 (.Q (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_7), .QB (\$dummy [980]), 
        .D (L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .CLK (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_8 (.Q (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_8), .QB (\$dummy [981]), 
        .D (L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .CLK (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_9 (.Q (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_9), .QB (\$dummy [982]), 
        .D (L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .CLK (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_10 (.Q (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_10), .QB (\$dummy [983])
        , .D (L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .CLK (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_11 (.Q (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_11), .QB (\$dummy [984])
        , .D (L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .CLK (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_12 (.Q (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_12), .QB (\$dummy [985])
        , .D (L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .CLK (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_13 (.Q (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_13), .QB (\$dummy [986])
        , .D (L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .CLK (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_14 (.Q (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_14), .QB (\$dummy [987])
        , .D (L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .CLK (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_15 (.Q (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_15), .QB (\$dummy [988])
        , .D (L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .CLK (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_16 (.Q (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_16), .QB (\$dummy [989])
        , .D (L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .CLK (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    inv02 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix623 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624), .A (CLK)) ;
    inv02 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix625 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626), .A (CLK)) ;
    inv02 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix627 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628), .A (CLK)) ;
    inv02 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix643 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644), .A (nx8378)) ;
    dff L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_0 (.Q (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_0), .QB (\$dummy [990]), 
        .D (L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .CLK (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    nor02_2x L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix567 (.Y (
             L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566), .A0 (RST), .A1 (
             L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644)) ;
    dff L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_1 (.Q (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_1), .QB (\$dummy [991]), 
        .D (L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .CLK (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_2 (.Q (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_2), .QB (\$dummy [992]), 
        .D (L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .CLK (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_3 (.Q (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_3), .QB (\$dummy [993]), 
        .D (L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .CLK (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_4 (.Q (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_4), .QB (\$dummy [994]), 
        .D (L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .CLK (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_5 (.Q (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_5), .QB (\$dummy [995]), 
        .D (L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .CLK (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_6 (.Q (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_6), .QB (\$dummy [996]), 
        .D (L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .CLK (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_7 (.Q (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_7), .QB (\$dummy [997]), 
        .D (L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .CLK (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_8 (.Q (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_8), .QB (\$dummy [998]), 
        .D (L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .CLK (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_9 (.Q (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_9), .QB (\$dummy [999]), 
        .D (L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .CLK (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_10 (.Q (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_10), .QB (\$dummy [1000])
        , .D (L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .CLK (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_11 (.Q (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_11), .QB (\$dummy [1001])
        , .D (L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .CLK (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_12 (.Q (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_12), .QB (\$dummy [1002])
        , .D (L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .CLK (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_13 (.Q (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_13), .QB (\$dummy [1003])
        , .D (L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .CLK (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_14 (.Q (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_14), .QB (\$dummy [1004])
        , .D (L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .CLK (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_15 (.Q (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_15), .QB (\$dummy [1005])
        , .D (L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .CLK (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_16 (.Q (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_16), .QB (\$dummy [1006])
        , .D (L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .CLK (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    inv02 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix623 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624), .A (CLK)) ;
    inv02 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix625 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626), .A (CLK)) ;
    inv02 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix627 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628), .A (CLK)) ;
    inv02 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix643 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644), .A (nx8384)) ;
    dff L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_0 (.Q (
        L1_3_L2_4_G3_MINI_ALU_BoothP_0), .QB (\$dummy [1007]), .D (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .CLK (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    nor02_2x L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix567 (.Y (
             L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566), .A0 (RST), .A1 (
             L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    dff L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_1 (.Q (
        L1_3_L2_4_G3_MINI_ALU_BoothP_1), .QB (\$dummy [1008]), .D (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .CLK (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_2 (.Q (
        L1_3_L2_4_G3_MINI_ALU_BoothP_2), .QB (\$dummy [1009]), .D (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .CLK (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_3 (.Q (
        L1_3_L2_4_G3_MINI_ALU_BoothP_3), .QB (\$dummy [1010]), .D (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .CLK (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_4 (.Q (
        L1_3_L2_4_G3_MINI_ALU_BoothP_4), .QB (\$dummy [1011]), .D (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .CLK (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_5 (.Q (
        L1_3_L2_4_G3_MINI_ALU_BoothP_5), .QB (\$dummy [1012]), .D (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .CLK (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_6 (.Q (
        L1_3_L2_4_G3_MINI_ALU_BoothP_6), .QB (\$dummy [1013]), .D (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .CLK (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_7 (.Q (
        L1_3_L2_4_G3_MINI_ALU_BoothP_7), .QB (\$dummy [1014]), .D (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .CLK (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_8 (.Q (
        L1_3_L2_4_G3_MINI_ALU_BoothP_8), .QB (\$dummy [1015]), .D (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .CLK (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_9 (.Q (
        L1_3_L2_4_G3_MINI_ALU_BoothP_9), .QB (\$dummy [1016]), .D (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .CLK (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_10 (.Q (
        L1_3_L2_4_G3_MINI_ALU_BoothP_10), .QB (\$dummy [1017]), .D (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .CLK (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_11 (.Q (
        L1_3_L2_4_G3_MINI_ALU_BoothP_11), .QB (\$dummy [1018]), .D (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .CLK (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_12 (.Q (
        L1_3_L2_4_G3_MINI_ALU_BoothP_12), .QB (\$dummy [1019]), .D (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .CLK (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_13 (.Q (
        L1_3_L2_4_G3_MINI_ALU_BoothP_13), .QB (\$dummy [1020]), .D (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .CLK (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_14 (.Q (
        L1_3_L2_4_G3_MINI_ALU_BoothP_14), .QB (\$dummy [1021]), .D (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .CLK (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_15 (.Q (
        L1_3_L2_4_G3_MINI_ALU_BoothP_15), .QB (\$dummy [1022]), .D (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .CLK (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_16 (.Q (
        L1_3_L2_4_G3_MINI_ALU_BoothP_16), .QB (\$dummy [1023]), .D (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .CLK (
        L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    inv02 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix623 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624), .A (CLK)) ;
    inv02 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix625 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626), .A (CLK)) ;
    inv02 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix627 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628), .A (CLK)) ;
    inv02 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix643 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644), .A (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642)) ;
    xor2 L1_4_L2_0_G3_MINI_ALU_ix83 (.Y (L3Results_1__0), .A0 (L2Results_3__0), 
         .A1 (L2Results_2__0)) ;
    xnor2 L1_4_L2_0_G3_MINI_ALU_ix380 (.Y (L1_4_L2_0_G3_MINI_ALU_nx379), .A0 (
          L1_4_L2_0_G3_MINI_ALU_nx381), .A1 (L1_4_L2_0_G3_MINI_ALU_nx383)) ;
    nand02 L1_4_L2_0_G3_MINI_ALU_ix382 (.Y (L1_4_L2_0_G3_MINI_ALU_nx381), .A0 (
           L1_4_L2_0_G3_MINI_ALU_BoothOperand_0), .A1 (nx8404)) ;
    xnor2 L1_4_L2_0_G3_MINI_ALU_ix384 (.Y (L1_4_L2_0_G3_MINI_ALU_nx383), .A0 (
          L1_4_L2_0_G3_MINI_ALU_BoothOperand_1), .A1 (
          L1_4_L2_0_G3_MINI_ALU_BoothP_1)) ;
    inv01 L1_4_L2_0_G3_MINI_ALU_ix388 (.Y (L1_4_L2_0_G3_MINI_ALU_nx387), .A (
          L1_4_L2_0_G3_MINI_ALU_BoothP_2)) ;
    xnor2 L1_4_L2_0_G3_MINI_ALU_ix390 (.Y (L1_4_L2_0_G3_MINI_ALU_nx389), .A0 (
          L1_4_L2_0_G3_MINI_ALU_nx391), .A1 (L1_4_L2_0_G3_MINI_ALU_nx395)) ;
    aoi32 L1_4_L2_0_G3_MINI_ALU_ix392 (.Y (L1_4_L2_0_G3_MINI_ALU_nx391), .A0 (
          L1_4_L2_0_G3_MINI_ALU_BoothOperand_0), .A1 (nx8404), .A2 (
          L1_4_L2_0_G3_MINI_ALU_nx154), .B0 (L1_4_L2_0_G3_MINI_ALU_BoothP_1), .B1 (
          L1_4_L2_0_G3_MINI_ALU_BoothOperand_1)) ;
    xnor2 L1_4_L2_0_G3_MINI_ALU_ix396 (.Y (L1_4_L2_0_G3_MINI_ALU_nx395), .A0 (
          L1_4_L2_0_G3_MINI_ALU_BoothOperand_2), .A1 (
          L1_4_L2_0_G3_MINI_ALU_BoothP_2)) ;
    inv01 L1_4_L2_0_G3_MINI_ALU_ix400 (.Y (L1_4_L2_0_G3_MINI_ALU_nx399), .A (
          L1_4_L2_0_G3_MINI_ALU_BoothP_3)) ;
    xnor2 L1_4_L2_0_G3_MINI_ALU_ix402 (.Y (L1_4_L2_0_G3_MINI_ALU_nx401), .A0 (
          L1_4_L2_0_G3_MINI_ALU_nx403), .A1 (L1_4_L2_0_G3_MINI_ALU_nx405)) ;
    xnor2 L1_4_L2_0_G3_MINI_ALU_ix406 (.Y (L1_4_L2_0_G3_MINI_ALU_nx405), .A0 (
          L1_4_L2_0_G3_MINI_ALU_BoothOperand_3), .A1 (
          L1_4_L2_0_G3_MINI_ALU_BoothP_3)) ;
    inv01 L1_4_L2_0_G3_MINI_ALU_ix410 (.Y (L1_4_L2_0_G3_MINI_ALU_nx409), .A (
          L1_4_L2_0_G3_MINI_ALU_BoothP_4)) ;
    xnor2 L1_4_L2_0_G3_MINI_ALU_ix412 (.Y (L1_4_L2_0_G3_MINI_ALU_nx411), .A0 (
          L1_4_L2_0_G3_MINI_ALU_nx413), .A1 (L1_4_L2_0_G3_MINI_ALU_nx415)) ;
    xnor2 L1_4_L2_0_G3_MINI_ALU_ix416 (.Y (L1_4_L2_0_G3_MINI_ALU_nx415), .A0 (
          L1_4_L2_0_G3_MINI_ALU_BoothOperand_4), .A1 (
          L1_4_L2_0_G3_MINI_ALU_BoothP_4)) ;
    inv01 L1_4_L2_0_G3_MINI_ALU_ix420 (.Y (L1_4_L2_0_G3_MINI_ALU_nx419), .A (
          L1_4_L2_0_G3_MINI_ALU_BoothP_5)) ;
    xnor2 L1_4_L2_0_G3_MINI_ALU_ix422 (.Y (L1_4_L2_0_G3_MINI_ALU_nx421), .A0 (
          L1_4_L2_0_G3_MINI_ALU_nx423), .A1 (L1_4_L2_0_G3_MINI_ALU_nx425)) ;
    xnor2 L1_4_L2_0_G3_MINI_ALU_ix426 (.Y (L1_4_L2_0_G3_MINI_ALU_nx425), .A0 (
          L1_4_L2_0_G3_MINI_ALU_BoothOperand_5), .A1 (
          L1_4_L2_0_G3_MINI_ALU_BoothP_5)) ;
    inv01 L1_4_L2_0_G3_MINI_ALU_ix430 (.Y (L1_4_L2_0_G3_MINI_ALU_nx429), .A (
          L1_4_L2_0_G3_MINI_ALU_BoothP_6)) ;
    xnor2 L1_4_L2_0_G3_MINI_ALU_ix432 (.Y (L1_4_L2_0_G3_MINI_ALU_nx431), .A0 (
          L1_4_L2_0_G3_MINI_ALU_nx433), .A1 (L1_4_L2_0_G3_MINI_ALU_nx435)) ;
    xnor2 L1_4_L2_0_G3_MINI_ALU_ix436 (.Y (L1_4_L2_0_G3_MINI_ALU_nx435), .A0 (
          L1_4_L2_0_G3_MINI_ALU_BoothOperand_6), .A1 (
          L1_4_L2_0_G3_MINI_ALU_BoothP_6)) ;
    inv01 L1_4_L2_0_G3_MINI_ALU_ix440 (.Y (L1_4_L2_0_G3_MINI_ALU_nx439), .A (
          L1_4_L2_0_G3_MINI_ALU_BoothP_7)) ;
    xnor2 L1_4_L2_0_G3_MINI_ALU_ix442 (.Y (L1_4_L2_0_G3_MINI_ALU_nx441), .A0 (
          L1_4_L2_0_G3_MINI_ALU_nx443), .A1 (L1_4_L2_0_G3_MINI_ALU_nx445)) ;
    xnor2 L1_4_L2_0_G3_MINI_ALU_ix446 (.Y (L1_4_L2_0_G3_MINI_ALU_nx445), .A0 (
          L1_4_L2_0_G3_MINI_ALU_BoothOperand_7), .A1 (
          L1_4_L2_0_G3_MINI_ALU_BoothP_7)) ;
    inv01 L1_4_L2_0_G3_MINI_ALU_ix450 (.Y (L1_4_L2_0_G3_MINI_ALU_nx449), .A (
          L1_4_L2_0_G3_MINI_ALU_BoothP_8)) ;
    xnor2 L1_4_L2_0_G3_MINI_ALU_ix452 (.Y (L1_4_L2_0_G3_MINI_ALU_nx451), .A0 (
          L1_4_L2_0_G3_MINI_ALU_nx453), .A1 (L1_4_L2_0_G3_MINI_ALU_nx455)) ;
    xnor2 L1_4_L2_0_G3_MINI_ALU_ix456 (.Y (L1_4_L2_0_G3_MINI_ALU_nx455), .A0 (
          L1_4_L2_0_G3_MINI_ALU_BoothOperand_8), .A1 (
          L1_4_L2_0_G3_MINI_ALU_BoothP_8)) ;
    xor2 L1_4_L2_0_G3_MINI_ALU_ix317 (.Y (L1_4_L2_0_G3_MINI_ALU_nx316), .A0 (
         L1_4_L2_0_G3_MINI_ALU_nx461), .A1 (L1_4_L2_0_G3_MINI_ALU_nx463)) ;
    xnor2 L1_4_L2_0_G3_MINI_ALU_ix464 (.Y (L1_4_L2_0_G3_MINI_ALU_nx463), .A0 (
          L1_4_L2_0_G3_MINI_ALU_BoothOperand_9), .A1 (
          L1_4_L2_0_G3_MINI_ALU_BoothP_9)) ;
    xor2 L1_4_L2_0_G3_MINI_ALU_ix337 (.Y (L1_4_L2_0_G3_MINI_ALU_nx336), .A0 (
         L1_4_L2_0_G3_MINI_ALU_nx467), .A1 (L1_4_L2_0_G3_MINI_ALU_nx471)) ;
    inv01 L1_4_L2_0_G3_MINI_ALU_ix470 (.Y (L1_4_L2_0_G3_MINI_ALU_nx469), .A (
          L1_4_L2_0_G3_MINI_ALU_BoothP_9)) ;
    xnor2 L1_4_L2_0_G3_MINI_ALU_ix472 (.Y (L1_4_L2_0_G3_MINI_ALU_nx471), .A0 (
          L1_4_L2_0_G3_MINI_ALU_BoothOperand_10), .A1 (
          L1_4_L2_0_G3_MINI_ALU_BoothP_10)) ;
    xor2 L1_4_L2_0_G3_MINI_ALU_ix357 (.Y (L1_4_L2_0_G3_MINI_ALU_nx356), .A0 (
         L1_4_L2_0_G3_MINI_ALU_nx475), .A1 (L1_4_L2_0_G3_MINI_ALU_nx479)) ;
    inv01 L1_4_L2_0_G3_MINI_ALU_ix478 (.Y (L1_4_L2_0_G3_MINI_ALU_nx477), .A (
          L1_4_L2_0_G3_MINI_ALU_BoothP_10)) ;
    xnor2 L1_4_L2_0_G3_MINI_ALU_ix480 (.Y (L1_4_L2_0_G3_MINI_ALU_nx479), .A0 (
          L1_4_L2_0_G3_MINI_ALU_BoothOperand_11), .A1 (
          L1_4_L2_0_G3_MINI_ALU_BoothP_11)) ;
    xor2 L1_4_L2_0_G3_MINI_ALU_ix377 (.Y (L1_4_L2_0_G3_MINI_ALU_nx376), .A0 (
         L1_4_L2_0_G3_MINI_ALU_nx483), .A1 (L1_4_L2_0_G3_MINI_ALU_nx487)) ;
    inv01 L1_4_L2_0_G3_MINI_ALU_ix486 (.Y (L1_4_L2_0_G3_MINI_ALU_nx485), .A (
          L1_4_L2_0_G3_MINI_ALU_BoothP_11)) ;
    xnor2 L1_4_L2_0_G3_MINI_ALU_ix488 (.Y (L1_4_L2_0_G3_MINI_ALU_nx487), .A0 (
          L1_4_L2_0_G3_MINI_ALU_BoothOperand_12), .A1 (
          L1_4_L2_0_G3_MINI_ALU_BoothP_12)) ;
    xor2 L1_4_L2_0_G3_MINI_ALU_ix397 (.Y (L1_4_L2_0_G3_MINI_ALU_nx396), .A0 (
         L1_4_L2_0_G3_MINI_ALU_nx491), .A1 (L1_4_L2_0_G3_MINI_ALU_nx495)) ;
    inv01 L1_4_L2_0_G3_MINI_ALU_ix494 (.Y (L1_4_L2_0_G3_MINI_ALU_nx493), .A (
          L1_4_L2_0_G3_MINI_ALU_BoothP_12)) ;
    xnor2 L1_4_L2_0_G3_MINI_ALU_ix496 (.Y (L1_4_L2_0_G3_MINI_ALU_nx495), .A0 (
          L1_4_L2_0_G3_MINI_ALU_BoothOperand_13), .A1 (
          L1_4_L2_0_G3_MINI_ALU_BoothP_13)) ;
    xor2 L1_4_L2_0_G3_MINI_ALU_ix417 (.Y (L1_4_L2_0_G3_MINI_ALU_nx416), .A0 (
         L1_4_L2_0_G3_MINI_ALU_nx499), .A1 (L1_4_L2_0_G3_MINI_ALU_nx503)) ;
    inv01 L1_4_L2_0_G3_MINI_ALU_ix502 (.Y (L1_4_L2_0_G3_MINI_ALU_nx501), .A (
          L1_4_L2_0_G3_MINI_ALU_BoothP_13)) ;
    xnor2 L1_4_L2_0_G3_MINI_ALU_ix504 (.Y (L1_4_L2_0_G3_MINI_ALU_nx503), .A0 (
          L1_4_L2_0_G3_MINI_ALU_BoothOperand_14), .A1 (
          L1_4_L2_0_G3_MINI_ALU_BoothP_14)) ;
    xor2 L1_4_L2_0_G3_MINI_ALU_ix437 (.Y (L1_4_L2_0_G3_MINI_ALU_nx436), .A0 (
         L1_4_L2_0_G3_MINI_ALU_nx507), .A1 (L1_4_L2_0_G3_MINI_ALU_nx511)) ;
    inv01 L1_4_L2_0_G3_MINI_ALU_ix510 (.Y (L1_4_L2_0_G3_MINI_ALU_nx509), .A (
          L1_4_L2_0_G3_MINI_ALU_BoothP_14)) ;
    xnor2 L1_4_L2_0_G3_MINI_ALU_ix512 (.Y (L1_4_L2_0_G3_MINI_ALU_nx511), .A0 (
          L1_4_L2_0_G3_MINI_ALU_BoothOperand_15), .A1 (
          L1_4_L2_0_G3_MINI_ALU_BoothP_15)) ;
    xnor2 L1_4_L2_0_G3_MINI_ALU_ix457 (.Y (L1_4_L2_0_G3_MINI_ALU_nx456), .A0 (
          L1_4_L2_0_G3_MINI_ALU_nx515), .A1 (L1_4_L2_0_G3_MINI_ALU_nx454)) ;
    inv01 L1_4_L2_0_G3_MINI_ALU_ix518 (.Y (L1_4_L2_0_G3_MINI_ALU_nx517), .A (
          L1_4_L2_0_G3_MINI_ALU_BoothP_15)) ;
    xor2 L1_4_L2_0_G3_MINI_ALU_ix455 (.Y (L1_4_L2_0_G3_MINI_ALU_nx454), .A0 (
         L1_4_L2_0_G3_MINI_ALU_BoothOperand_16), .A1 (
         L1_4_L2_0_G3_MINI_ALU_BoothP_16)) ;
    mux21_ni L1_4_L2_0_G3_MINI_ALU_ix91 (.Y (L1FirstOperands_5__0), .A0 (
             L1_4_L2_0_G3_MINI_ALU_BoothP_1), .A1 (WindowDin_4__0__0), .S0 (
             Instr)) ;
    mux21_ni L1_4_L2_0_G3_MINI_ALU_ix99 (.Y (L1FirstOperands_5__1), .A0 (
             L1_4_L2_0_G3_MINI_ALU_BoothP_2), .A1 (WindowDin_4__0__1), .S0 (
             Instr)) ;
    mux21_ni L1_4_L2_0_G3_MINI_ALU_ix107 (.Y (L1FirstOperands_5__2), .A0 (
             L1_4_L2_0_G3_MINI_ALU_BoothP_3), .A1 (WindowDin_4__0__2), .S0 (
             Instr)) ;
    mux21_ni L1_4_L2_0_G3_MINI_ALU_ix115 (.Y (L1FirstOperands_5__3), .A0 (
             L1_4_L2_0_G3_MINI_ALU_BoothP_4), .A1 (WindowDin_4__0__3), .S0 (
             Instr)) ;
    mux21_ni L1_4_L2_0_G3_MINI_ALU_ix123 (.Y (L1FirstOperands_5__4), .A0 (
             L1_4_L2_0_G3_MINI_ALU_BoothP_5), .A1 (WindowDin_4__0__4), .S0 (
             Instr)) ;
    mux21_ni L1_4_L2_0_G3_MINI_ALU_ix131 (.Y (L1FirstOperands_5__5), .A0 (
             L1_4_L2_0_G3_MINI_ALU_BoothP_6), .A1 (WindowDin_4__0__5), .S0 (
             Instr)) ;
    mux21_ni L1_4_L2_0_G3_MINI_ALU_ix139 (.Y (L1FirstOperands_5__6), .A0 (
             L1_4_L2_0_G3_MINI_ALU_BoothP_7), .A1 (WindowDin_4__0__6), .S0 (
             Instr)) ;
    mux21_ni L1_4_L2_0_G3_MINI_ALU_ix147 (.Y (L1FirstOperands_5__7), .A0 (
             L1_4_L2_0_G3_MINI_ALU_BoothP_8), .A1 (WindowDin_4__0__7), .S0 (
             Instr)) ;
    xor2 L1_4_L2_0_G3_MINI_ALU_ix77 (.Y (L3Results_1__1), .A0 (
         L1_4_L2_0_G3_MINI_ALU_nx529), .A1 (L1_4_L2_0_G3_MINI_ALU_nx531)) ;
    nand02 L1_4_L2_0_G3_MINI_ALU_ix530 (.Y (L1_4_L2_0_G3_MINI_ALU_nx529), .A0 (
           L2Results_3__0), .A1 (L2Results_2__0)) ;
    xnor2 L1_4_L2_0_G3_MINI_ALU_ix532 (.Y (L1_4_L2_0_G3_MINI_ALU_nx531), .A0 (
          L2Results_3__1), .A1 (L2Results_2__1)) ;
    xor2 L1_4_L2_0_G3_MINI_ALU_ix75 (.Y (L3Results_1__2), .A0 (
         L1_4_L2_0_G3_MINI_ALU_nx534), .A1 (L1_4_L2_0_G3_MINI_ALU_nx537)) ;
    aoi32 L1_4_L2_0_G3_MINI_ALU_ix535 (.Y (L1_4_L2_0_G3_MINI_ALU_nx534), .A0 (
          L2Results_3__0), .A1 (L2Results_2__0), .A2 (L1_4_L2_0_G3_MINI_ALU_nx30
          ), .B0 (L2Results_2__1), .B1 (L2Results_3__1)) ;
    xnor2 L1_4_L2_0_G3_MINI_ALU_ix538 (.Y (L1_4_L2_0_G3_MINI_ALU_nx537), .A0 (
          L2Results_3__2), .A1 (L2Results_2__2)) ;
    xor2 L1_4_L2_0_G3_MINI_ALU_ix73 (.Y (L3Results_1__3), .A0 (
         L1_4_L2_0_G3_MINI_ALU_nx540), .A1 (L1_4_L2_0_G3_MINI_ALU_nx544)) ;
    aoi22 L1_4_L2_0_G3_MINI_ALU_ix541 (.Y (L1_4_L2_0_G3_MINI_ALU_nx540), .A0 (
          L2Results_2__2), .A1 (L2Results_3__2), .B0 (L1_4_L2_0_G3_MINI_ALU_nx40
          ), .B1 (L1_4_L2_0_G3_MINI_ALU_nx24)) ;
    xnor2 L1_4_L2_0_G3_MINI_ALU_ix545 (.Y (L1_4_L2_0_G3_MINI_ALU_nx544), .A0 (
          L2Results_3__3), .A1 (L2Results_2__3)) ;
    xor2 L1_4_L2_0_G3_MINI_ALU_ix71 (.Y (L3Results_1__4), .A0 (
         L1_4_L2_0_G3_MINI_ALU_nx547), .A1 (L1_4_L2_0_G3_MINI_ALU_nx551)) ;
    aoi22 L1_4_L2_0_G3_MINI_ALU_ix548 (.Y (L1_4_L2_0_G3_MINI_ALU_nx547), .A0 (
          L2Results_2__3), .A1 (L2Results_3__3), .B0 (L1_4_L2_0_G3_MINI_ALU_nx44
          ), .B1 (L1_4_L2_0_G3_MINI_ALU_nx18)) ;
    xnor2 L1_4_L2_0_G3_MINI_ALU_ix552 (.Y (L1_4_L2_0_G3_MINI_ALU_nx551), .A0 (
          L2Results_3__4), .A1 (L2Results_2__4)) ;
    xor2 L1_4_L2_0_G3_MINI_ALU_ix69 (.Y (L3Results_1__5), .A0 (
         L1_4_L2_0_G3_MINI_ALU_nx554), .A1 (L1_4_L2_0_G3_MINI_ALU_nx558)) ;
    aoi22 L1_4_L2_0_G3_MINI_ALU_ix555 (.Y (L1_4_L2_0_G3_MINI_ALU_nx554), .A0 (
          L2Results_2__4), .A1 (L2Results_3__4), .B0 (L1_4_L2_0_G3_MINI_ALU_nx48
          ), .B1 (L1_4_L2_0_G3_MINI_ALU_nx12)) ;
    xnor2 L1_4_L2_0_G3_MINI_ALU_ix559 (.Y (L1_4_L2_0_G3_MINI_ALU_nx558), .A0 (
          L2Results_3__5), .A1 (L2Results_2__5)) ;
    xor2 L1_4_L2_0_G3_MINI_ALU_ix67 (.Y (L3Results_1__6), .A0 (
         L1_4_L2_0_G3_MINI_ALU_nx561), .A1 (L1_4_L2_0_G3_MINI_ALU_nx565)) ;
    aoi22 L1_4_L2_0_G3_MINI_ALU_ix562 (.Y (L1_4_L2_0_G3_MINI_ALU_nx561), .A0 (
          L2Results_2__5), .A1 (L2Results_3__5), .B0 (L1_4_L2_0_G3_MINI_ALU_nx52
          ), .B1 (L1_4_L2_0_G3_MINI_ALU_nx6)) ;
    xnor2 L1_4_L2_0_G3_MINI_ALU_ix566 (.Y (L1_4_L2_0_G3_MINI_ALU_nx565), .A0 (
          L2Results_3__6), .A1 (L2Results_2__6)) ;
    xnor2 L1_4_L2_0_G3_MINI_ALU_ix65 (.Y (L3Results_1__7), .A0 (
          L1_4_L2_0_G3_MINI_ALU_nx568), .A1 (L1_4_L2_0_G3_MINI_ALU_nx62)) ;
    aoi22 L1_4_L2_0_G3_MINI_ALU_ix569 (.Y (L1_4_L2_0_G3_MINI_ALU_nx568), .A0 (
          L2Results_2__6), .A1 (L2Results_3__6), .B0 (L1_4_L2_0_G3_MINI_ALU_nx56
          ), .B1 (L1_4_L2_0_G3_MINI_ALU_nx0)) ;
    xor2 L1_4_L2_0_G3_MINI_ALU_ix63 (.Y (L1_4_L2_0_G3_MINI_ALU_nx62), .A0 (
         L2Results_3__7), .A1 (L2Results_2__7)) ;
    inv01 L1_4_L2_0_G3_MINI_ALU_ix155 (.Y (L1_4_L2_0_G3_MINI_ALU_nx154), .A (
          L1_4_L2_0_G3_MINI_ALU_nx383)) ;
    inv01 L1_4_L2_0_G3_MINI_ALU_ix57 (.Y (L1_4_L2_0_G3_MINI_ALU_nx56), .A (
          L1_4_L2_0_G3_MINI_ALU_nx561)) ;
    inv01 L1_4_L2_0_G3_MINI_ALU_ix53 (.Y (L1_4_L2_0_G3_MINI_ALU_nx52), .A (
          L1_4_L2_0_G3_MINI_ALU_nx554)) ;
    inv01 L1_4_L2_0_G3_MINI_ALU_ix49 (.Y (L1_4_L2_0_G3_MINI_ALU_nx48), .A (
          L1_4_L2_0_G3_MINI_ALU_nx547)) ;
    inv01 L1_4_L2_0_G3_MINI_ALU_ix45 (.Y (L1_4_L2_0_G3_MINI_ALU_nx44), .A (
          L1_4_L2_0_G3_MINI_ALU_nx540)) ;
    inv01 L1_4_L2_0_G3_MINI_ALU_ix41 (.Y (L1_4_L2_0_G3_MINI_ALU_nx40), .A (
          L1_4_L2_0_G3_MINI_ALU_nx534)) ;
    inv01 L1_4_L2_0_G3_MINI_ALU_ix31 (.Y (L1_4_L2_0_G3_MINI_ALU_nx30), .A (
          L1_4_L2_0_G3_MINI_ALU_nx531)) ;
    inv01 L1_4_L2_0_G3_MINI_ALU_ix25 (.Y (L1_4_L2_0_G3_MINI_ALU_nx24), .A (
          L1_4_L2_0_G3_MINI_ALU_nx537)) ;
    inv01 L1_4_L2_0_G3_MINI_ALU_ix19 (.Y (L1_4_L2_0_G3_MINI_ALU_nx18), .A (
          L1_4_L2_0_G3_MINI_ALU_nx544)) ;
    inv01 L1_4_L2_0_G3_MINI_ALU_ix13 (.Y (L1_4_L2_0_G3_MINI_ALU_nx12), .A (
          L1_4_L2_0_G3_MINI_ALU_nx551)) ;
    inv01 L1_4_L2_0_G3_MINI_ALU_ix7 (.Y (L1_4_L2_0_G3_MINI_ALU_nx6), .A (
          L1_4_L2_0_G3_MINI_ALU_nx558)) ;
    inv01 L1_4_L2_0_G3_MINI_ALU_ix1 (.Y (L1_4_L2_0_G3_MINI_ALU_nx0), .A (
          L1_4_L2_0_G3_MINI_ALU_nx565)) ;
    fake_gnd L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix216 (.Y (
             L1_4_L2_0_G3_MINI_ALU_WindowCellShiftedLeft_16)) ;
    nor02ii L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix81 (.Y (
            L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_nx80), .A0 (Instr), .A1 (Start)) ;
    aoi21 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix77 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_10), .A0 (
          FilterDin_4__0__1), .A1 (FilterDin_4__0__0), .B0 (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_nx4)) ;
    nor02_2x L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix5 (.Y (
             L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_nx4), .A0 (FilterDin_4__0__0), .A1 (
             FilterDin_4__0__1)) ;
    aoi21 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix67 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_11), .A0 (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_nx328), .A1 (FilterDin_4__0__2), .B0 (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_nx8)) ;
    nor03_2x L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix9 (.Y (
             L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_nx8), .A0 (FilterDin_4__0__2), .A1 (
             FilterDin_4__0__0), .A2 (FilterDin_4__0__1)) ;
    xnor2 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix59 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_12), .A0 (
          FilterDin_4__0__3), .A1 (L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_nx8)) ;
    xnor2 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix51 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_13), .A0 (
          FilterDin_4__0__4), .A1 (L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_nx12)) ;
    nor04 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix13 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_nx12), .A0 (FilterDin_4__0__3), .A1 (
          FilterDin_4__0__2), .A2 (FilterDin_4__0__0), .A3 (FilterDin_4__0__1)
          ) ;
    xnor2 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix43 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_14), .A0 (
          FilterDin_4__0__5), .A1 (L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_nx16)) ;
    nor02ii L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix17 (.Y (
            L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_nx16), .A0 (FilterDin_4__0__4), .A1 (
            L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_nx12)) ;
    xnor2 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix35 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_15), .A0 (
          FilterDin_4__0__6), .A1 (L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_nx20)) ;
    nor02ii L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix21 (.Y (
            L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_nx20), .A0 (FilterDin_4__0__5), .A1 (
            L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_nx16)) ;
    xnor2 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix27 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_16), .A0 (
          FilterDin_4__0__7), .A1 (L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_nx24)) ;
    nor02ii L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix25 (.Y (
            L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_nx24), .A0 (FilterDin_4__0__6), .A1 (
            L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_nx20)) ;
    inv01 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix329 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_nx328), .A (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_nx4)) ;
    inv02 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix383 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_nx384), .A (
          L1_4_L2_0_G3_MINI_ALU_BoothP_0)) ;
    dff L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_0 (.Q (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_0), .QB (\$dummy [1024])
        , .D (L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .CLK (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    nor02_2x L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix567 (.Y (
             L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566), .A0 (RST), .A1 (
             L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644)) ;
    dff L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_1 (.Q (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_1), .QB (\$dummy [1025])
        , .D (L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .CLK (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_2 (.Q (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_2), .QB (\$dummy [1026])
        , .D (L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .CLK (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_3 (.Q (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_3), .QB (\$dummy [1027])
        , .D (L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .CLK (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_4 (.Q (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_4), .QB (\$dummy [1028])
        , .D (L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .CLK (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_5 (.Q (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_5), .QB (\$dummy [1029])
        , .D (L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .CLK (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_6 (.Q (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_6), .QB (\$dummy [1030])
        , .D (L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .CLK (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_7 (.Q (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_7), .QB (\$dummy [1031])
        , .D (L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .CLK (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_8 (.Q (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_8), .QB (\$dummy [1032])
        , .D (L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .CLK (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_9 (.Q (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_9), .QB (\$dummy [1033])
        , .D (L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .CLK (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_10 (.Q (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_10), .QB (\$dummy [1034])
        , .D (L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .CLK (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_11 (.Q (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_11), .QB (\$dummy [1035])
        , .D (L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .CLK (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_12 (.Q (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_12), .QB (\$dummy [1036])
        , .D (L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .CLK (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_13 (.Q (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_13), .QB (\$dummy [1037])
        , .D (L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .CLK (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_14 (.Q (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_14), .QB (\$dummy [1038])
        , .D (L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .CLK (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_15 (.Q (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_15), .QB (\$dummy [1039])
        , .D (L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .CLK (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_16 (.Q (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_16), .QB (\$dummy [1040])
        , .D (L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .CLK (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    inv02 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix623 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624), .A (CLK)) ;
    inv02 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix625 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626), .A (CLK)) ;
    inv02 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix627 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628), .A (CLK)) ;
    inv02 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix643 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644), .A (nx8418)) ;
    dff L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_0 (.Q (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_0), .QB (\$dummy [1041])
        , .D (L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .CLK (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    nor02_2x L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix567 (.Y (
             L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566), .A0 (RST), .A1 (
             L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644)) ;
    dff L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_1 (.Q (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_1), .QB (\$dummy [1042])
        , .D (L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .CLK (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_2 (.Q (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_2), .QB (\$dummy [1043])
        , .D (L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .CLK (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_3 (.Q (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_3), .QB (\$dummy [1044])
        , .D (L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .CLK (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_4 (.Q (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_4), .QB (\$dummy [1045])
        , .D (L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .CLK (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_5 (.Q (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_5), .QB (\$dummy [1046])
        , .D (L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .CLK (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_6 (.Q (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_6), .QB (\$dummy [1047])
        , .D (L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .CLK (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_7 (.Q (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_7), .QB (\$dummy [1048])
        , .D (L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .CLK (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_8 (.Q (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_8), .QB (\$dummy [1049])
        , .D (L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .CLK (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_9 (.Q (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_9), .QB (\$dummy [1050])
        , .D (L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .CLK (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_10 (.Q (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_10), .QB (\$dummy [1051])
        , .D (L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .CLK (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_11 (.Q (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_11), .QB (\$dummy [1052])
        , .D (L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .CLK (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_12 (.Q (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_12), .QB (\$dummy [1053])
        , .D (L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .CLK (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_13 (.Q (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_13), .QB (\$dummy [1054])
        , .D (L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .CLK (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_14 (.Q (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_14), .QB (\$dummy [1055])
        , .D (L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .CLK (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_15 (.Q (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_15), .QB (\$dummy [1056])
        , .D (L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .CLK (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_16 (.Q (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_16), .QB (\$dummy [1057])
        , .D (L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .CLK (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    inv02 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix623 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624), .A (CLK)) ;
    inv02 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix625 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626), .A (CLK)) ;
    inv02 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix627 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628), .A (CLK)) ;
    inv02 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix643 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644), .A (nx8424)) ;
    dff L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_0 (.Q (
        L1_4_L2_0_G3_MINI_ALU_BoothP_0), .QB (\$dummy [1058]), .D (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .CLK (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    nor02_2x L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix567 (.Y (
             L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566), .A0 (RST), .A1 (
             L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    dff L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_1 (.Q (
        L1_4_L2_0_G3_MINI_ALU_BoothP_1), .QB (\$dummy [1059]), .D (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .CLK (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_2 (.Q (
        L1_4_L2_0_G3_MINI_ALU_BoothP_2), .QB (\$dummy [1060]), .D (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .CLK (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_3 (.Q (
        L1_4_L2_0_G3_MINI_ALU_BoothP_3), .QB (\$dummy [1061]), .D (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .CLK (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_4 (.Q (
        L1_4_L2_0_G3_MINI_ALU_BoothP_4), .QB (\$dummy [1062]), .D (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .CLK (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_5 (.Q (
        L1_4_L2_0_G3_MINI_ALU_BoothP_5), .QB (\$dummy [1063]), .D (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .CLK (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_6 (.Q (
        L1_4_L2_0_G3_MINI_ALU_BoothP_6), .QB (\$dummy [1064]), .D (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .CLK (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_7 (.Q (
        L1_4_L2_0_G3_MINI_ALU_BoothP_7), .QB (\$dummy [1065]), .D (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .CLK (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_8 (.Q (
        L1_4_L2_0_G3_MINI_ALU_BoothP_8), .QB (\$dummy [1066]), .D (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .CLK (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_9 (.Q (
        L1_4_L2_0_G3_MINI_ALU_BoothP_9), .QB (\$dummy [1067]), .D (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .CLK (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_10 (.Q (
        L1_4_L2_0_G3_MINI_ALU_BoothP_10), .QB (\$dummy [1068]), .D (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .CLK (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_11 (.Q (
        L1_4_L2_0_G3_MINI_ALU_BoothP_11), .QB (\$dummy [1069]), .D (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .CLK (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_12 (.Q (
        L1_4_L2_0_G3_MINI_ALU_BoothP_12), .QB (\$dummy [1070]), .D (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .CLK (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_13 (.Q (
        L1_4_L2_0_G3_MINI_ALU_BoothP_13), .QB (\$dummy [1071]), .D (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .CLK (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_14 (.Q (
        L1_4_L2_0_G3_MINI_ALU_BoothP_14), .QB (\$dummy [1072]), .D (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .CLK (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_15 (.Q (
        L1_4_L2_0_G3_MINI_ALU_BoothP_15), .QB (\$dummy [1073]), .D (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .CLK (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_16 (.Q (
        L1_4_L2_0_G3_MINI_ALU_BoothP_16), .QB (\$dummy [1074]), .D (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .CLK (
        L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    inv02 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix623 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624), .A (CLK)) ;
    inv02 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix625 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626), .A (CLK)) ;
    inv02 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix627 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628), .A (CLK)) ;
    inv02 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix643 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644), .A (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642)) ;
    xor2 L1_4_L2_1_G3_MINI_ALU_ix83 (.Y (L3Results_2__0), .A0 (L2Results_5__0), 
         .A1 (L2Results_4__0)) ;
    xnor2 L1_4_L2_1_G3_MINI_ALU_ix380 (.Y (L1_4_L2_1_G3_MINI_ALU_nx379), .A0 (
          L1_4_L2_1_G3_MINI_ALU_nx381), .A1 (L1_4_L2_1_G3_MINI_ALU_nx383)) ;
    nand02 L1_4_L2_1_G3_MINI_ALU_ix382 (.Y (L1_4_L2_1_G3_MINI_ALU_nx381), .A0 (
           L1_4_L2_1_G3_MINI_ALU_BoothOperand_0), .A1 (nx8444)) ;
    xnor2 L1_4_L2_1_G3_MINI_ALU_ix384 (.Y (L1_4_L2_1_G3_MINI_ALU_nx383), .A0 (
          L1_4_L2_1_G3_MINI_ALU_BoothOperand_1), .A1 (
          L1_4_L2_1_G3_MINI_ALU_BoothP_1)) ;
    inv01 L1_4_L2_1_G3_MINI_ALU_ix388 (.Y (L1_4_L2_1_G3_MINI_ALU_nx387), .A (
          L1_4_L2_1_G3_MINI_ALU_BoothP_2)) ;
    xnor2 L1_4_L2_1_G3_MINI_ALU_ix390 (.Y (L1_4_L2_1_G3_MINI_ALU_nx389), .A0 (
          L1_4_L2_1_G3_MINI_ALU_nx391), .A1 (L1_4_L2_1_G3_MINI_ALU_nx395)) ;
    aoi32 L1_4_L2_1_G3_MINI_ALU_ix392 (.Y (L1_4_L2_1_G3_MINI_ALU_nx391), .A0 (
          L1_4_L2_1_G3_MINI_ALU_BoothOperand_0), .A1 (nx8444), .A2 (
          L1_4_L2_1_G3_MINI_ALU_nx154), .B0 (L1_4_L2_1_G3_MINI_ALU_BoothP_1), .B1 (
          L1_4_L2_1_G3_MINI_ALU_BoothOperand_1)) ;
    xnor2 L1_4_L2_1_G3_MINI_ALU_ix396 (.Y (L1_4_L2_1_G3_MINI_ALU_nx395), .A0 (
          L1_4_L2_1_G3_MINI_ALU_BoothOperand_2), .A1 (
          L1_4_L2_1_G3_MINI_ALU_BoothP_2)) ;
    inv01 L1_4_L2_1_G3_MINI_ALU_ix400 (.Y (L1_4_L2_1_G3_MINI_ALU_nx399), .A (
          L1_4_L2_1_G3_MINI_ALU_BoothP_3)) ;
    xnor2 L1_4_L2_1_G3_MINI_ALU_ix402 (.Y (L1_4_L2_1_G3_MINI_ALU_nx401), .A0 (
          L1_4_L2_1_G3_MINI_ALU_nx403), .A1 (L1_4_L2_1_G3_MINI_ALU_nx405)) ;
    xnor2 L1_4_L2_1_G3_MINI_ALU_ix406 (.Y (L1_4_L2_1_G3_MINI_ALU_nx405), .A0 (
          L1_4_L2_1_G3_MINI_ALU_BoothOperand_3), .A1 (
          L1_4_L2_1_G3_MINI_ALU_BoothP_3)) ;
    inv01 L1_4_L2_1_G3_MINI_ALU_ix410 (.Y (L1_4_L2_1_G3_MINI_ALU_nx409), .A (
          L1_4_L2_1_G3_MINI_ALU_BoothP_4)) ;
    xnor2 L1_4_L2_1_G3_MINI_ALU_ix412 (.Y (L1_4_L2_1_G3_MINI_ALU_nx411), .A0 (
          L1_4_L2_1_G3_MINI_ALU_nx413), .A1 (L1_4_L2_1_G3_MINI_ALU_nx415)) ;
    xnor2 L1_4_L2_1_G3_MINI_ALU_ix416 (.Y (L1_4_L2_1_G3_MINI_ALU_nx415), .A0 (
          L1_4_L2_1_G3_MINI_ALU_BoothOperand_4), .A1 (
          L1_4_L2_1_G3_MINI_ALU_BoothP_4)) ;
    inv01 L1_4_L2_1_G3_MINI_ALU_ix420 (.Y (L1_4_L2_1_G3_MINI_ALU_nx419), .A (
          L1_4_L2_1_G3_MINI_ALU_BoothP_5)) ;
    xnor2 L1_4_L2_1_G3_MINI_ALU_ix422 (.Y (L1_4_L2_1_G3_MINI_ALU_nx421), .A0 (
          L1_4_L2_1_G3_MINI_ALU_nx423), .A1 (L1_4_L2_1_G3_MINI_ALU_nx425)) ;
    xnor2 L1_4_L2_1_G3_MINI_ALU_ix426 (.Y (L1_4_L2_1_G3_MINI_ALU_nx425), .A0 (
          L1_4_L2_1_G3_MINI_ALU_BoothOperand_5), .A1 (
          L1_4_L2_1_G3_MINI_ALU_BoothP_5)) ;
    inv01 L1_4_L2_1_G3_MINI_ALU_ix430 (.Y (L1_4_L2_1_G3_MINI_ALU_nx429), .A (
          L1_4_L2_1_G3_MINI_ALU_BoothP_6)) ;
    xnor2 L1_4_L2_1_G3_MINI_ALU_ix432 (.Y (L1_4_L2_1_G3_MINI_ALU_nx431), .A0 (
          L1_4_L2_1_G3_MINI_ALU_nx433), .A1 (L1_4_L2_1_G3_MINI_ALU_nx435)) ;
    xnor2 L1_4_L2_1_G3_MINI_ALU_ix436 (.Y (L1_4_L2_1_G3_MINI_ALU_nx435), .A0 (
          L1_4_L2_1_G3_MINI_ALU_BoothOperand_6), .A1 (
          L1_4_L2_1_G3_MINI_ALU_BoothP_6)) ;
    inv01 L1_4_L2_1_G3_MINI_ALU_ix440 (.Y (L1_4_L2_1_G3_MINI_ALU_nx439), .A (
          L1_4_L2_1_G3_MINI_ALU_BoothP_7)) ;
    xnor2 L1_4_L2_1_G3_MINI_ALU_ix442 (.Y (L1_4_L2_1_G3_MINI_ALU_nx441), .A0 (
          L1_4_L2_1_G3_MINI_ALU_nx443), .A1 (L1_4_L2_1_G3_MINI_ALU_nx445)) ;
    xnor2 L1_4_L2_1_G3_MINI_ALU_ix446 (.Y (L1_4_L2_1_G3_MINI_ALU_nx445), .A0 (
          L1_4_L2_1_G3_MINI_ALU_BoothOperand_7), .A1 (
          L1_4_L2_1_G3_MINI_ALU_BoothP_7)) ;
    inv01 L1_4_L2_1_G3_MINI_ALU_ix450 (.Y (L1_4_L2_1_G3_MINI_ALU_nx449), .A (
          L1_4_L2_1_G3_MINI_ALU_BoothP_8)) ;
    xnor2 L1_4_L2_1_G3_MINI_ALU_ix452 (.Y (L1_4_L2_1_G3_MINI_ALU_nx451), .A0 (
          L1_4_L2_1_G3_MINI_ALU_nx453), .A1 (L1_4_L2_1_G3_MINI_ALU_nx455)) ;
    xnor2 L1_4_L2_1_G3_MINI_ALU_ix456 (.Y (L1_4_L2_1_G3_MINI_ALU_nx455), .A0 (
          L1_4_L2_1_G3_MINI_ALU_BoothOperand_8), .A1 (
          L1_4_L2_1_G3_MINI_ALU_BoothP_8)) ;
    xor2 L1_4_L2_1_G3_MINI_ALU_ix317 (.Y (L1_4_L2_1_G3_MINI_ALU_nx316), .A0 (
         L1_4_L2_1_G3_MINI_ALU_nx461), .A1 (L1_4_L2_1_G3_MINI_ALU_nx463)) ;
    xnor2 L1_4_L2_1_G3_MINI_ALU_ix464 (.Y (L1_4_L2_1_G3_MINI_ALU_nx463), .A0 (
          L1_4_L2_1_G3_MINI_ALU_BoothOperand_9), .A1 (
          L1_4_L2_1_G3_MINI_ALU_BoothP_9)) ;
    xor2 L1_4_L2_1_G3_MINI_ALU_ix337 (.Y (L1_4_L2_1_G3_MINI_ALU_nx336), .A0 (
         L1_4_L2_1_G3_MINI_ALU_nx467), .A1 (L1_4_L2_1_G3_MINI_ALU_nx471)) ;
    inv01 L1_4_L2_1_G3_MINI_ALU_ix470 (.Y (L1_4_L2_1_G3_MINI_ALU_nx469), .A (
          L1_4_L2_1_G3_MINI_ALU_BoothP_9)) ;
    xnor2 L1_4_L2_1_G3_MINI_ALU_ix472 (.Y (L1_4_L2_1_G3_MINI_ALU_nx471), .A0 (
          L1_4_L2_1_G3_MINI_ALU_BoothOperand_10), .A1 (
          L1_4_L2_1_G3_MINI_ALU_BoothP_10)) ;
    xor2 L1_4_L2_1_G3_MINI_ALU_ix357 (.Y (L1_4_L2_1_G3_MINI_ALU_nx356), .A0 (
         L1_4_L2_1_G3_MINI_ALU_nx475), .A1 (L1_4_L2_1_G3_MINI_ALU_nx479)) ;
    inv01 L1_4_L2_1_G3_MINI_ALU_ix478 (.Y (L1_4_L2_1_G3_MINI_ALU_nx477), .A (
          L1_4_L2_1_G3_MINI_ALU_BoothP_10)) ;
    xnor2 L1_4_L2_1_G3_MINI_ALU_ix480 (.Y (L1_4_L2_1_G3_MINI_ALU_nx479), .A0 (
          L1_4_L2_1_G3_MINI_ALU_BoothOperand_11), .A1 (
          L1_4_L2_1_G3_MINI_ALU_BoothP_11)) ;
    xor2 L1_4_L2_1_G3_MINI_ALU_ix377 (.Y (L1_4_L2_1_G3_MINI_ALU_nx376), .A0 (
         L1_4_L2_1_G3_MINI_ALU_nx483), .A1 (L1_4_L2_1_G3_MINI_ALU_nx487)) ;
    inv01 L1_4_L2_1_G3_MINI_ALU_ix486 (.Y (L1_4_L2_1_G3_MINI_ALU_nx485), .A (
          L1_4_L2_1_G3_MINI_ALU_BoothP_11)) ;
    xnor2 L1_4_L2_1_G3_MINI_ALU_ix488 (.Y (L1_4_L2_1_G3_MINI_ALU_nx487), .A0 (
          L1_4_L2_1_G3_MINI_ALU_BoothOperand_12), .A1 (
          L1_4_L2_1_G3_MINI_ALU_BoothP_12)) ;
    xor2 L1_4_L2_1_G3_MINI_ALU_ix397 (.Y (L1_4_L2_1_G3_MINI_ALU_nx396), .A0 (
         L1_4_L2_1_G3_MINI_ALU_nx491), .A1 (L1_4_L2_1_G3_MINI_ALU_nx495)) ;
    inv01 L1_4_L2_1_G3_MINI_ALU_ix494 (.Y (L1_4_L2_1_G3_MINI_ALU_nx493), .A (
          L1_4_L2_1_G3_MINI_ALU_BoothP_12)) ;
    xnor2 L1_4_L2_1_G3_MINI_ALU_ix496 (.Y (L1_4_L2_1_G3_MINI_ALU_nx495), .A0 (
          L1_4_L2_1_G3_MINI_ALU_BoothOperand_13), .A1 (
          L1_4_L2_1_G3_MINI_ALU_BoothP_13)) ;
    xor2 L1_4_L2_1_G3_MINI_ALU_ix417 (.Y (L1_4_L2_1_G3_MINI_ALU_nx416), .A0 (
         L1_4_L2_1_G3_MINI_ALU_nx499), .A1 (L1_4_L2_1_G3_MINI_ALU_nx503)) ;
    inv01 L1_4_L2_1_G3_MINI_ALU_ix502 (.Y (L1_4_L2_1_G3_MINI_ALU_nx501), .A (
          L1_4_L2_1_G3_MINI_ALU_BoothP_13)) ;
    xnor2 L1_4_L2_1_G3_MINI_ALU_ix504 (.Y (L1_4_L2_1_G3_MINI_ALU_nx503), .A0 (
          L1_4_L2_1_G3_MINI_ALU_BoothOperand_14), .A1 (
          L1_4_L2_1_G3_MINI_ALU_BoothP_14)) ;
    xor2 L1_4_L2_1_G3_MINI_ALU_ix437 (.Y (L1_4_L2_1_G3_MINI_ALU_nx436), .A0 (
         L1_4_L2_1_G3_MINI_ALU_nx507), .A1 (L1_4_L2_1_G3_MINI_ALU_nx511)) ;
    inv01 L1_4_L2_1_G3_MINI_ALU_ix510 (.Y (L1_4_L2_1_G3_MINI_ALU_nx509), .A (
          L1_4_L2_1_G3_MINI_ALU_BoothP_14)) ;
    xnor2 L1_4_L2_1_G3_MINI_ALU_ix512 (.Y (L1_4_L2_1_G3_MINI_ALU_nx511), .A0 (
          L1_4_L2_1_G3_MINI_ALU_BoothOperand_15), .A1 (
          L1_4_L2_1_G3_MINI_ALU_BoothP_15)) ;
    xnor2 L1_4_L2_1_G3_MINI_ALU_ix457 (.Y (L1_4_L2_1_G3_MINI_ALU_nx456), .A0 (
          L1_4_L2_1_G3_MINI_ALU_nx515), .A1 (L1_4_L2_1_G3_MINI_ALU_nx454)) ;
    inv01 L1_4_L2_1_G3_MINI_ALU_ix518 (.Y (L1_4_L2_1_G3_MINI_ALU_nx517), .A (
          L1_4_L2_1_G3_MINI_ALU_BoothP_15)) ;
    xor2 L1_4_L2_1_G3_MINI_ALU_ix455 (.Y (L1_4_L2_1_G3_MINI_ALU_nx454), .A0 (
         L1_4_L2_1_G3_MINI_ALU_BoothOperand_16), .A1 (
         L1_4_L2_1_G3_MINI_ALU_BoothP_16)) ;
    mux21_ni L1_4_L2_1_G3_MINI_ALU_ix91 (.Y (L1FirstOperands_9__0), .A0 (
             L1_4_L2_1_G3_MINI_ALU_BoothP_1), .A1 (WindowDin_4__1__0), .S0 (
             Instr)) ;
    mux21_ni L1_4_L2_1_G3_MINI_ALU_ix99 (.Y (L1FirstOperands_9__1), .A0 (
             L1_4_L2_1_G3_MINI_ALU_BoothP_2), .A1 (WindowDin_4__1__1), .S0 (
             Instr)) ;
    mux21_ni L1_4_L2_1_G3_MINI_ALU_ix107 (.Y (L1FirstOperands_9__2), .A0 (
             L1_4_L2_1_G3_MINI_ALU_BoothP_3), .A1 (WindowDin_4__1__2), .S0 (
             Instr)) ;
    mux21_ni L1_4_L2_1_G3_MINI_ALU_ix115 (.Y (L1FirstOperands_9__3), .A0 (
             L1_4_L2_1_G3_MINI_ALU_BoothP_4), .A1 (WindowDin_4__1__3), .S0 (
             Instr)) ;
    mux21_ni L1_4_L2_1_G3_MINI_ALU_ix123 (.Y (L1FirstOperands_9__4), .A0 (
             L1_4_L2_1_G3_MINI_ALU_BoothP_5), .A1 (WindowDin_4__1__4), .S0 (
             Instr)) ;
    mux21_ni L1_4_L2_1_G3_MINI_ALU_ix131 (.Y (L1FirstOperands_9__5), .A0 (
             L1_4_L2_1_G3_MINI_ALU_BoothP_6), .A1 (WindowDin_4__1__5), .S0 (
             Instr)) ;
    mux21_ni L1_4_L2_1_G3_MINI_ALU_ix139 (.Y (L1FirstOperands_9__6), .A0 (
             L1_4_L2_1_G3_MINI_ALU_BoothP_7), .A1 (WindowDin_4__1__6), .S0 (
             Instr)) ;
    mux21_ni L1_4_L2_1_G3_MINI_ALU_ix147 (.Y (L1FirstOperands_9__7), .A0 (
             L1_4_L2_1_G3_MINI_ALU_BoothP_8), .A1 (WindowDin_4__1__7), .S0 (
             Instr)) ;
    xor2 L1_4_L2_1_G3_MINI_ALU_ix77 (.Y (L3Results_2__1), .A0 (
         L1_4_L2_1_G3_MINI_ALU_nx529), .A1 (L1_4_L2_1_G3_MINI_ALU_nx531)) ;
    nand02 L1_4_L2_1_G3_MINI_ALU_ix530 (.Y (L1_4_L2_1_G3_MINI_ALU_nx529), .A0 (
           L2Results_5__0), .A1 (L2Results_4__0)) ;
    xnor2 L1_4_L2_1_G3_MINI_ALU_ix532 (.Y (L1_4_L2_1_G3_MINI_ALU_nx531), .A0 (
          L2Results_5__1), .A1 (L2Results_4__1)) ;
    xor2 L1_4_L2_1_G3_MINI_ALU_ix75 (.Y (L3Results_2__2), .A0 (
         L1_4_L2_1_G3_MINI_ALU_nx534), .A1 (L1_4_L2_1_G3_MINI_ALU_nx537)) ;
    aoi32 L1_4_L2_1_G3_MINI_ALU_ix535 (.Y (L1_4_L2_1_G3_MINI_ALU_nx534), .A0 (
          L2Results_5__0), .A1 (L2Results_4__0), .A2 (L1_4_L2_1_G3_MINI_ALU_nx30
          ), .B0 (L2Results_4__1), .B1 (L2Results_5__1)) ;
    xnor2 L1_4_L2_1_G3_MINI_ALU_ix538 (.Y (L1_4_L2_1_G3_MINI_ALU_nx537), .A0 (
          L2Results_5__2), .A1 (L2Results_4__2)) ;
    xor2 L1_4_L2_1_G3_MINI_ALU_ix73 (.Y (L3Results_2__3), .A0 (
         L1_4_L2_1_G3_MINI_ALU_nx540), .A1 (L1_4_L2_1_G3_MINI_ALU_nx544)) ;
    aoi22 L1_4_L2_1_G3_MINI_ALU_ix541 (.Y (L1_4_L2_1_G3_MINI_ALU_nx540), .A0 (
          L2Results_4__2), .A1 (L2Results_5__2), .B0 (L1_4_L2_1_G3_MINI_ALU_nx40
          ), .B1 (L1_4_L2_1_G3_MINI_ALU_nx24)) ;
    xnor2 L1_4_L2_1_G3_MINI_ALU_ix545 (.Y (L1_4_L2_1_G3_MINI_ALU_nx544), .A0 (
          L2Results_5__3), .A1 (L2Results_4__3)) ;
    xor2 L1_4_L2_1_G3_MINI_ALU_ix71 (.Y (L3Results_2__4), .A0 (
         L1_4_L2_1_G3_MINI_ALU_nx547), .A1 (L1_4_L2_1_G3_MINI_ALU_nx551)) ;
    aoi22 L1_4_L2_1_G3_MINI_ALU_ix548 (.Y (L1_4_L2_1_G3_MINI_ALU_nx547), .A0 (
          L2Results_4__3), .A1 (L2Results_5__3), .B0 (L1_4_L2_1_G3_MINI_ALU_nx44
          ), .B1 (L1_4_L2_1_G3_MINI_ALU_nx18)) ;
    xnor2 L1_4_L2_1_G3_MINI_ALU_ix552 (.Y (L1_4_L2_1_G3_MINI_ALU_nx551), .A0 (
          L2Results_5__4), .A1 (L2Results_4__4)) ;
    xor2 L1_4_L2_1_G3_MINI_ALU_ix69 (.Y (L3Results_2__5), .A0 (
         L1_4_L2_1_G3_MINI_ALU_nx554), .A1 (L1_4_L2_1_G3_MINI_ALU_nx558)) ;
    aoi22 L1_4_L2_1_G3_MINI_ALU_ix555 (.Y (L1_4_L2_1_G3_MINI_ALU_nx554), .A0 (
          L2Results_4__4), .A1 (L2Results_5__4), .B0 (L1_4_L2_1_G3_MINI_ALU_nx48
          ), .B1 (L1_4_L2_1_G3_MINI_ALU_nx12)) ;
    xnor2 L1_4_L2_1_G3_MINI_ALU_ix559 (.Y (L1_4_L2_1_G3_MINI_ALU_nx558), .A0 (
          L2Results_5__5), .A1 (L2Results_4__5)) ;
    xor2 L1_4_L2_1_G3_MINI_ALU_ix67 (.Y (L3Results_2__6), .A0 (
         L1_4_L2_1_G3_MINI_ALU_nx561), .A1 (L1_4_L2_1_G3_MINI_ALU_nx565)) ;
    aoi22 L1_4_L2_1_G3_MINI_ALU_ix562 (.Y (L1_4_L2_1_G3_MINI_ALU_nx561), .A0 (
          L2Results_4__5), .A1 (L2Results_5__5), .B0 (L1_4_L2_1_G3_MINI_ALU_nx52
          ), .B1 (L1_4_L2_1_G3_MINI_ALU_nx6)) ;
    xnor2 L1_4_L2_1_G3_MINI_ALU_ix566 (.Y (L1_4_L2_1_G3_MINI_ALU_nx565), .A0 (
          L2Results_5__6), .A1 (L2Results_4__6)) ;
    xnor2 L1_4_L2_1_G3_MINI_ALU_ix65 (.Y (L3Results_2__7), .A0 (
          L1_4_L2_1_G3_MINI_ALU_nx568), .A1 (L1_4_L2_1_G3_MINI_ALU_nx62)) ;
    aoi22 L1_4_L2_1_G3_MINI_ALU_ix569 (.Y (L1_4_L2_1_G3_MINI_ALU_nx568), .A0 (
          L2Results_4__6), .A1 (L2Results_5__6), .B0 (L1_4_L2_1_G3_MINI_ALU_nx56
          ), .B1 (L1_4_L2_1_G3_MINI_ALU_nx0)) ;
    xor2 L1_4_L2_1_G3_MINI_ALU_ix63 (.Y (L1_4_L2_1_G3_MINI_ALU_nx62), .A0 (
         L2Results_5__7), .A1 (L2Results_4__7)) ;
    inv01 L1_4_L2_1_G3_MINI_ALU_ix155 (.Y (L1_4_L2_1_G3_MINI_ALU_nx154), .A (
          L1_4_L2_1_G3_MINI_ALU_nx383)) ;
    inv01 L1_4_L2_1_G3_MINI_ALU_ix57 (.Y (L1_4_L2_1_G3_MINI_ALU_nx56), .A (
          L1_4_L2_1_G3_MINI_ALU_nx561)) ;
    inv01 L1_4_L2_1_G3_MINI_ALU_ix53 (.Y (L1_4_L2_1_G3_MINI_ALU_nx52), .A (
          L1_4_L2_1_G3_MINI_ALU_nx554)) ;
    inv01 L1_4_L2_1_G3_MINI_ALU_ix49 (.Y (L1_4_L2_1_G3_MINI_ALU_nx48), .A (
          L1_4_L2_1_G3_MINI_ALU_nx547)) ;
    inv01 L1_4_L2_1_G3_MINI_ALU_ix45 (.Y (L1_4_L2_1_G3_MINI_ALU_nx44), .A (
          L1_4_L2_1_G3_MINI_ALU_nx540)) ;
    inv01 L1_4_L2_1_G3_MINI_ALU_ix41 (.Y (L1_4_L2_1_G3_MINI_ALU_nx40), .A (
          L1_4_L2_1_G3_MINI_ALU_nx534)) ;
    inv01 L1_4_L2_1_G3_MINI_ALU_ix31 (.Y (L1_4_L2_1_G3_MINI_ALU_nx30), .A (
          L1_4_L2_1_G3_MINI_ALU_nx531)) ;
    inv01 L1_4_L2_1_G3_MINI_ALU_ix25 (.Y (L1_4_L2_1_G3_MINI_ALU_nx24), .A (
          L1_4_L2_1_G3_MINI_ALU_nx537)) ;
    inv01 L1_4_L2_1_G3_MINI_ALU_ix19 (.Y (L1_4_L2_1_G3_MINI_ALU_nx18), .A (
          L1_4_L2_1_G3_MINI_ALU_nx544)) ;
    inv01 L1_4_L2_1_G3_MINI_ALU_ix13 (.Y (L1_4_L2_1_G3_MINI_ALU_nx12), .A (
          L1_4_L2_1_G3_MINI_ALU_nx551)) ;
    inv01 L1_4_L2_1_G3_MINI_ALU_ix7 (.Y (L1_4_L2_1_G3_MINI_ALU_nx6), .A (
          L1_4_L2_1_G3_MINI_ALU_nx558)) ;
    inv01 L1_4_L2_1_G3_MINI_ALU_ix1 (.Y (L1_4_L2_1_G3_MINI_ALU_nx0), .A (
          L1_4_L2_1_G3_MINI_ALU_nx565)) ;
    fake_gnd L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix216 (.Y (
             L1_4_L2_1_G3_MINI_ALU_WindowCellShiftedLeft_16)) ;
    nor02ii L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix81 (.Y (
            L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_nx80), .A0 (Instr), .A1 (Start)) ;
    aoi21 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix77 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_10), .A0 (
          FilterDin_4__1__1), .A1 (FilterDin_4__1__0), .B0 (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_nx4)) ;
    nor02_2x L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix5 (.Y (
             L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_nx4), .A0 (FilterDin_4__1__0), .A1 (
             FilterDin_4__1__1)) ;
    aoi21 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix67 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_11), .A0 (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_nx328), .A1 (FilterDin_4__1__2), .B0 (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_nx8)) ;
    nor03_2x L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix9 (.Y (
             L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_nx8), .A0 (FilterDin_4__1__2), .A1 (
             FilterDin_4__1__0), .A2 (FilterDin_4__1__1)) ;
    xnor2 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix59 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_12), .A0 (
          FilterDin_4__1__3), .A1 (L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_nx8)) ;
    xnor2 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix51 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_13), .A0 (
          FilterDin_4__1__4), .A1 (L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_nx12)) ;
    nor04 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix13 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_nx12), .A0 (FilterDin_4__1__3), .A1 (
          FilterDin_4__1__2), .A2 (FilterDin_4__1__0), .A3 (FilterDin_4__1__1)
          ) ;
    xnor2 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix43 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_14), .A0 (
          FilterDin_4__1__5), .A1 (L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_nx16)) ;
    nor02ii L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix17 (.Y (
            L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_nx16), .A0 (FilterDin_4__1__4), .A1 (
            L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_nx12)) ;
    xnor2 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix35 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_15), .A0 (
          FilterDin_4__1__6), .A1 (L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_nx20)) ;
    nor02ii L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix21 (.Y (
            L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_nx20), .A0 (FilterDin_4__1__5), .A1 (
            L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_nx16)) ;
    xnor2 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix27 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_16), .A0 (
          FilterDin_4__1__7), .A1 (L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_nx24)) ;
    nor02ii L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix25 (.Y (
            L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_nx24), .A0 (FilterDin_4__1__6), .A1 (
            L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_nx20)) ;
    inv01 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix329 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_nx328), .A (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_nx4)) ;
    inv02 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix383 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_nx384), .A (
          L1_4_L2_1_G3_MINI_ALU_BoothP_0)) ;
    dff L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_0 (.Q (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_0), .QB (\$dummy [1075])
        , .D (L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .CLK (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    nor02_2x L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix567 (.Y (
             L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566), .A0 (RST), .A1 (
             L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644)) ;
    dff L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_1 (.Q (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_1), .QB (\$dummy [1076])
        , .D (L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .CLK (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_2 (.Q (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_2), .QB (\$dummy [1077])
        , .D (L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .CLK (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_3 (.Q (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_3), .QB (\$dummy [1078])
        , .D (L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .CLK (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_4 (.Q (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_4), .QB (\$dummy [1079])
        , .D (L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .CLK (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_5 (.Q (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_5), .QB (\$dummy [1080])
        , .D (L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .CLK (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_6 (.Q (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_6), .QB (\$dummy [1081])
        , .D (L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .CLK (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_7 (.Q (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_7), .QB (\$dummy [1082])
        , .D (L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .CLK (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_8 (.Q (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_8), .QB (\$dummy [1083])
        , .D (L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .CLK (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_9 (.Q (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_9), .QB (\$dummy [1084])
        , .D (L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .CLK (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_10 (.Q (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_10), .QB (\$dummy [1085])
        , .D (L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .CLK (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_11 (.Q (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_11), .QB (\$dummy [1086])
        , .D (L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .CLK (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_12 (.Q (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_12), .QB (\$dummy [1087])
        , .D (L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .CLK (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_13 (.Q (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_13), .QB (\$dummy [1088])
        , .D (L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .CLK (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_14 (.Q (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_14), .QB (\$dummy [1089])
        , .D (L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .CLK (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_15 (.Q (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_15), .QB (\$dummy [1090])
        , .D (L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .CLK (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_16 (.Q (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_16), .QB (\$dummy [1091])
        , .D (L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .CLK (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    inv02 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix623 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624), .A (CLK)) ;
    inv02 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix625 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626), .A (CLK)) ;
    inv02 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix627 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628), .A (CLK)) ;
    inv02 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix643 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644), .A (nx8458)) ;
    dff L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_0 (.Q (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_0), .QB (\$dummy [1092])
        , .D (L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .CLK (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    nor02_2x L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix567 (.Y (
             L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566), .A0 (RST), .A1 (
             L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644)) ;
    dff L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_1 (.Q (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_1), .QB (\$dummy [1093])
        , .D (L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .CLK (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_2 (.Q (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_2), .QB (\$dummy [1094])
        , .D (L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .CLK (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_3 (.Q (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_3), .QB (\$dummy [1095])
        , .D (L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .CLK (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_4 (.Q (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_4), .QB (\$dummy [1096])
        , .D (L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .CLK (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_5 (.Q (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_5), .QB (\$dummy [1097])
        , .D (L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .CLK (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_6 (.Q (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_6), .QB (\$dummy [1098])
        , .D (L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .CLK (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_7 (.Q (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_7), .QB (\$dummy [1099])
        , .D (L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .CLK (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_8 (.Q (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_8), .QB (\$dummy [1100])
        , .D (L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .CLK (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_9 (.Q (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_9), .QB (\$dummy [1101])
        , .D (L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .CLK (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_10 (.Q (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_10), .QB (\$dummy [1102])
        , .D (L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .CLK (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_11 (.Q (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_11), .QB (\$dummy [1103])
        , .D (L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .CLK (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_12 (.Q (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_12), .QB (\$dummy [1104])
        , .D (L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .CLK (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_13 (.Q (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_13), .QB (\$dummy [1105])
        , .D (L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .CLK (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_14 (.Q (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_14), .QB (\$dummy [1106])
        , .D (L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .CLK (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_15 (.Q (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_15), .QB (\$dummy [1107])
        , .D (L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .CLK (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_16 (.Q (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_16), .QB (\$dummy [1108])
        , .D (L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .CLK (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    inv02 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix623 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624), .A (CLK)) ;
    inv02 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix625 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626), .A (CLK)) ;
    inv02 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix627 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628), .A (CLK)) ;
    inv02 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix643 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644), .A (nx8464)) ;
    dff L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_0 (.Q (
        L1_4_L2_1_G3_MINI_ALU_BoothP_0), .QB (\$dummy [1109]), .D (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .CLK (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    nor02_2x L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix567 (.Y (
             L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566), .A0 (RST), .A1 (
             L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    dff L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_1 (.Q (
        L1_4_L2_1_G3_MINI_ALU_BoothP_1), .QB (\$dummy [1110]), .D (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .CLK (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_2 (.Q (
        L1_4_L2_1_G3_MINI_ALU_BoothP_2), .QB (\$dummy [1111]), .D (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .CLK (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_3 (.Q (
        L1_4_L2_1_G3_MINI_ALU_BoothP_3), .QB (\$dummy [1112]), .D (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .CLK (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_4 (.Q (
        L1_4_L2_1_G3_MINI_ALU_BoothP_4), .QB (\$dummy [1113]), .D (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .CLK (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_5 (.Q (
        L1_4_L2_1_G3_MINI_ALU_BoothP_5), .QB (\$dummy [1114]), .D (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .CLK (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_6 (.Q (
        L1_4_L2_1_G3_MINI_ALU_BoothP_6), .QB (\$dummy [1115]), .D (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .CLK (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_7 (.Q (
        L1_4_L2_1_G3_MINI_ALU_BoothP_7), .QB (\$dummy [1116]), .D (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .CLK (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_8 (.Q (
        L1_4_L2_1_G3_MINI_ALU_BoothP_8), .QB (\$dummy [1117]), .D (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .CLK (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_9 (.Q (
        L1_4_L2_1_G3_MINI_ALU_BoothP_9), .QB (\$dummy [1118]), .D (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .CLK (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_10 (.Q (
        L1_4_L2_1_G3_MINI_ALU_BoothP_10), .QB (\$dummy [1119]), .D (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .CLK (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_11 (.Q (
        L1_4_L2_1_G3_MINI_ALU_BoothP_11), .QB (\$dummy [1120]), .D (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .CLK (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_12 (.Q (
        L1_4_L2_1_G3_MINI_ALU_BoothP_12), .QB (\$dummy [1121]), .D (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .CLK (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_13 (.Q (
        L1_4_L2_1_G3_MINI_ALU_BoothP_13), .QB (\$dummy [1122]), .D (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .CLK (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_14 (.Q (
        L1_4_L2_1_G3_MINI_ALU_BoothP_14), .QB (\$dummy [1123]), .D (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .CLK (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_15 (.Q (
        L1_4_L2_1_G3_MINI_ALU_BoothP_15), .QB (\$dummy [1124]), .D (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .CLK (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_16 (.Q (
        L1_4_L2_1_G3_MINI_ALU_BoothP_16), .QB (\$dummy [1125]), .D (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .CLK (
        L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    inv02 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix623 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624), .A (CLK)) ;
    inv02 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix625 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626), .A (CLK)) ;
    inv02 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix627 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628), .A (CLK)) ;
    inv02 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix643 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644), .A (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642)) ;
    xor2 L1_4_L2_2_G4_MINI_ALU_ix83 (.Y (L4Results_0__0), .A0 (L3Results_1__0), 
         .A1 (L3Results_0__0)) ;
    xnor2 L1_4_L2_2_G4_MINI_ALU_ix380 (.Y (L1_4_L2_2_G4_MINI_ALU_nx379), .A0 (
          L1_4_L2_2_G4_MINI_ALU_nx381), .A1 (L1_4_L2_2_G4_MINI_ALU_nx383)) ;
    nand02 L1_4_L2_2_G4_MINI_ALU_ix382 (.Y (L1_4_L2_2_G4_MINI_ALU_nx381), .A0 (
           L1_4_L2_2_G4_MINI_ALU_BoothOperand_0), .A1 (nx8484)) ;
    xnor2 L1_4_L2_2_G4_MINI_ALU_ix384 (.Y (L1_4_L2_2_G4_MINI_ALU_nx383), .A0 (
          L1_4_L2_2_G4_MINI_ALU_BoothOperand_1), .A1 (
          L1_4_L2_2_G4_MINI_ALU_BoothP_1)) ;
    inv01 L1_4_L2_2_G4_MINI_ALU_ix388 (.Y (L1_4_L2_2_G4_MINI_ALU_nx387), .A (
          L1_4_L2_2_G4_MINI_ALU_BoothP_2)) ;
    xnor2 L1_4_L2_2_G4_MINI_ALU_ix390 (.Y (L1_4_L2_2_G4_MINI_ALU_nx389), .A0 (
          L1_4_L2_2_G4_MINI_ALU_nx391), .A1 (L1_4_L2_2_G4_MINI_ALU_nx395)) ;
    aoi32 L1_4_L2_2_G4_MINI_ALU_ix392 (.Y (L1_4_L2_2_G4_MINI_ALU_nx391), .A0 (
          L1_4_L2_2_G4_MINI_ALU_BoothOperand_0), .A1 (nx8484), .A2 (
          L1_4_L2_2_G4_MINI_ALU_nx154), .B0 (L1_4_L2_2_G4_MINI_ALU_BoothP_1), .B1 (
          L1_4_L2_2_G4_MINI_ALU_BoothOperand_1)) ;
    xnor2 L1_4_L2_2_G4_MINI_ALU_ix396 (.Y (L1_4_L2_2_G4_MINI_ALU_nx395), .A0 (
          L1_4_L2_2_G4_MINI_ALU_BoothOperand_2), .A1 (
          L1_4_L2_2_G4_MINI_ALU_BoothP_2)) ;
    inv01 L1_4_L2_2_G4_MINI_ALU_ix400 (.Y (L1_4_L2_2_G4_MINI_ALU_nx399), .A (
          L1_4_L2_2_G4_MINI_ALU_BoothP_3)) ;
    xnor2 L1_4_L2_2_G4_MINI_ALU_ix402 (.Y (L1_4_L2_2_G4_MINI_ALU_nx401), .A0 (
          L1_4_L2_2_G4_MINI_ALU_nx403), .A1 (L1_4_L2_2_G4_MINI_ALU_nx405)) ;
    xnor2 L1_4_L2_2_G4_MINI_ALU_ix406 (.Y (L1_4_L2_2_G4_MINI_ALU_nx405), .A0 (
          L1_4_L2_2_G4_MINI_ALU_BoothOperand_3), .A1 (
          L1_4_L2_2_G4_MINI_ALU_BoothP_3)) ;
    inv01 L1_4_L2_2_G4_MINI_ALU_ix410 (.Y (L1_4_L2_2_G4_MINI_ALU_nx409), .A (
          L1_4_L2_2_G4_MINI_ALU_BoothP_4)) ;
    xnor2 L1_4_L2_2_G4_MINI_ALU_ix412 (.Y (L1_4_L2_2_G4_MINI_ALU_nx411), .A0 (
          L1_4_L2_2_G4_MINI_ALU_nx413), .A1 (L1_4_L2_2_G4_MINI_ALU_nx415)) ;
    xnor2 L1_4_L2_2_G4_MINI_ALU_ix416 (.Y (L1_4_L2_2_G4_MINI_ALU_nx415), .A0 (
          L1_4_L2_2_G4_MINI_ALU_BoothOperand_4), .A1 (
          L1_4_L2_2_G4_MINI_ALU_BoothP_4)) ;
    inv01 L1_4_L2_2_G4_MINI_ALU_ix420 (.Y (L1_4_L2_2_G4_MINI_ALU_nx419), .A (
          L1_4_L2_2_G4_MINI_ALU_BoothP_5)) ;
    xnor2 L1_4_L2_2_G4_MINI_ALU_ix422 (.Y (L1_4_L2_2_G4_MINI_ALU_nx421), .A0 (
          L1_4_L2_2_G4_MINI_ALU_nx423), .A1 (L1_4_L2_2_G4_MINI_ALU_nx425)) ;
    xnor2 L1_4_L2_2_G4_MINI_ALU_ix426 (.Y (L1_4_L2_2_G4_MINI_ALU_nx425), .A0 (
          L1_4_L2_2_G4_MINI_ALU_BoothOperand_5), .A1 (
          L1_4_L2_2_G4_MINI_ALU_BoothP_5)) ;
    inv01 L1_4_L2_2_G4_MINI_ALU_ix430 (.Y (L1_4_L2_2_G4_MINI_ALU_nx429), .A (
          L1_4_L2_2_G4_MINI_ALU_BoothP_6)) ;
    xnor2 L1_4_L2_2_G4_MINI_ALU_ix432 (.Y (L1_4_L2_2_G4_MINI_ALU_nx431), .A0 (
          L1_4_L2_2_G4_MINI_ALU_nx433), .A1 (L1_4_L2_2_G4_MINI_ALU_nx435)) ;
    xnor2 L1_4_L2_2_G4_MINI_ALU_ix436 (.Y (L1_4_L2_2_G4_MINI_ALU_nx435), .A0 (
          L1_4_L2_2_G4_MINI_ALU_BoothOperand_6), .A1 (
          L1_4_L2_2_G4_MINI_ALU_BoothP_6)) ;
    inv01 L1_4_L2_2_G4_MINI_ALU_ix440 (.Y (L1_4_L2_2_G4_MINI_ALU_nx439), .A (
          L1_4_L2_2_G4_MINI_ALU_BoothP_7)) ;
    xnor2 L1_4_L2_2_G4_MINI_ALU_ix442 (.Y (L1_4_L2_2_G4_MINI_ALU_nx441), .A0 (
          L1_4_L2_2_G4_MINI_ALU_nx443), .A1 (L1_4_L2_2_G4_MINI_ALU_nx445)) ;
    xnor2 L1_4_L2_2_G4_MINI_ALU_ix446 (.Y (L1_4_L2_2_G4_MINI_ALU_nx445), .A0 (
          L1_4_L2_2_G4_MINI_ALU_BoothOperand_7), .A1 (
          L1_4_L2_2_G4_MINI_ALU_BoothP_7)) ;
    inv01 L1_4_L2_2_G4_MINI_ALU_ix450 (.Y (L1_4_L2_2_G4_MINI_ALU_nx449), .A (
          L1_4_L2_2_G4_MINI_ALU_BoothP_8)) ;
    xnor2 L1_4_L2_2_G4_MINI_ALU_ix452 (.Y (L1_4_L2_2_G4_MINI_ALU_nx451), .A0 (
          L1_4_L2_2_G4_MINI_ALU_nx453), .A1 (L1_4_L2_2_G4_MINI_ALU_nx455)) ;
    xnor2 L1_4_L2_2_G4_MINI_ALU_ix456 (.Y (L1_4_L2_2_G4_MINI_ALU_nx455), .A0 (
          L1_4_L2_2_G4_MINI_ALU_BoothOperand_8), .A1 (
          L1_4_L2_2_G4_MINI_ALU_BoothP_8)) ;
    xor2 L1_4_L2_2_G4_MINI_ALU_ix317 (.Y (L1_4_L2_2_G4_MINI_ALU_nx316), .A0 (
         L1_4_L2_2_G4_MINI_ALU_nx461), .A1 (L1_4_L2_2_G4_MINI_ALU_nx463)) ;
    xnor2 L1_4_L2_2_G4_MINI_ALU_ix464 (.Y (L1_4_L2_2_G4_MINI_ALU_nx463), .A0 (
          L1_4_L2_2_G4_MINI_ALU_BoothOperand_9), .A1 (
          L1_4_L2_2_G4_MINI_ALU_BoothP_9)) ;
    xor2 L1_4_L2_2_G4_MINI_ALU_ix337 (.Y (L1_4_L2_2_G4_MINI_ALU_nx336), .A0 (
         L1_4_L2_2_G4_MINI_ALU_nx467), .A1 (L1_4_L2_2_G4_MINI_ALU_nx471)) ;
    inv01 L1_4_L2_2_G4_MINI_ALU_ix470 (.Y (L1_4_L2_2_G4_MINI_ALU_nx469), .A (
          L1_4_L2_2_G4_MINI_ALU_BoothP_9)) ;
    xnor2 L1_4_L2_2_G4_MINI_ALU_ix472 (.Y (L1_4_L2_2_G4_MINI_ALU_nx471), .A0 (
          L1_4_L2_2_G4_MINI_ALU_BoothOperand_10), .A1 (
          L1_4_L2_2_G4_MINI_ALU_BoothP_10)) ;
    xor2 L1_4_L2_2_G4_MINI_ALU_ix357 (.Y (L1_4_L2_2_G4_MINI_ALU_nx356), .A0 (
         L1_4_L2_2_G4_MINI_ALU_nx475), .A1 (L1_4_L2_2_G4_MINI_ALU_nx479)) ;
    inv01 L1_4_L2_2_G4_MINI_ALU_ix478 (.Y (L1_4_L2_2_G4_MINI_ALU_nx477), .A (
          L1_4_L2_2_G4_MINI_ALU_BoothP_10)) ;
    xnor2 L1_4_L2_2_G4_MINI_ALU_ix480 (.Y (L1_4_L2_2_G4_MINI_ALU_nx479), .A0 (
          L1_4_L2_2_G4_MINI_ALU_BoothOperand_11), .A1 (
          L1_4_L2_2_G4_MINI_ALU_BoothP_11)) ;
    xor2 L1_4_L2_2_G4_MINI_ALU_ix377 (.Y (L1_4_L2_2_G4_MINI_ALU_nx376), .A0 (
         L1_4_L2_2_G4_MINI_ALU_nx483), .A1 (L1_4_L2_2_G4_MINI_ALU_nx487)) ;
    inv01 L1_4_L2_2_G4_MINI_ALU_ix486 (.Y (L1_4_L2_2_G4_MINI_ALU_nx485), .A (
          L1_4_L2_2_G4_MINI_ALU_BoothP_11)) ;
    xnor2 L1_4_L2_2_G4_MINI_ALU_ix488 (.Y (L1_4_L2_2_G4_MINI_ALU_nx487), .A0 (
          L1_4_L2_2_G4_MINI_ALU_BoothOperand_12), .A1 (
          L1_4_L2_2_G4_MINI_ALU_BoothP_12)) ;
    xor2 L1_4_L2_2_G4_MINI_ALU_ix397 (.Y (L1_4_L2_2_G4_MINI_ALU_nx396), .A0 (
         L1_4_L2_2_G4_MINI_ALU_nx491), .A1 (L1_4_L2_2_G4_MINI_ALU_nx495)) ;
    inv01 L1_4_L2_2_G4_MINI_ALU_ix494 (.Y (L1_4_L2_2_G4_MINI_ALU_nx493), .A (
          L1_4_L2_2_G4_MINI_ALU_BoothP_12)) ;
    xnor2 L1_4_L2_2_G4_MINI_ALU_ix496 (.Y (L1_4_L2_2_G4_MINI_ALU_nx495), .A0 (
          L1_4_L2_2_G4_MINI_ALU_BoothOperand_13), .A1 (
          L1_4_L2_2_G4_MINI_ALU_BoothP_13)) ;
    xor2 L1_4_L2_2_G4_MINI_ALU_ix417 (.Y (L1_4_L2_2_G4_MINI_ALU_nx416), .A0 (
         L1_4_L2_2_G4_MINI_ALU_nx499), .A1 (L1_4_L2_2_G4_MINI_ALU_nx503)) ;
    inv01 L1_4_L2_2_G4_MINI_ALU_ix502 (.Y (L1_4_L2_2_G4_MINI_ALU_nx501), .A (
          L1_4_L2_2_G4_MINI_ALU_BoothP_13)) ;
    xnor2 L1_4_L2_2_G4_MINI_ALU_ix504 (.Y (L1_4_L2_2_G4_MINI_ALU_nx503), .A0 (
          L1_4_L2_2_G4_MINI_ALU_BoothOperand_14), .A1 (
          L1_4_L2_2_G4_MINI_ALU_BoothP_14)) ;
    xor2 L1_4_L2_2_G4_MINI_ALU_ix437 (.Y (L1_4_L2_2_G4_MINI_ALU_nx436), .A0 (
         L1_4_L2_2_G4_MINI_ALU_nx507), .A1 (L1_4_L2_2_G4_MINI_ALU_nx511)) ;
    inv01 L1_4_L2_2_G4_MINI_ALU_ix510 (.Y (L1_4_L2_2_G4_MINI_ALU_nx509), .A (
          L1_4_L2_2_G4_MINI_ALU_BoothP_14)) ;
    xnor2 L1_4_L2_2_G4_MINI_ALU_ix512 (.Y (L1_4_L2_2_G4_MINI_ALU_nx511), .A0 (
          L1_4_L2_2_G4_MINI_ALU_BoothOperand_15), .A1 (
          L1_4_L2_2_G4_MINI_ALU_BoothP_15)) ;
    xnor2 L1_4_L2_2_G4_MINI_ALU_ix457 (.Y (L1_4_L2_2_G4_MINI_ALU_nx456), .A0 (
          L1_4_L2_2_G4_MINI_ALU_nx515), .A1 (L1_4_L2_2_G4_MINI_ALU_nx454)) ;
    inv01 L1_4_L2_2_G4_MINI_ALU_ix518 (.Y (L1_4_L2_2_G4_MINI_ALU_nx517), .A (
          L1_4_L2_2_G4_MINI_ALU_BoothP_15)) ;
    xor2 L1_4_L2_2_G4_MINI_ALU_ix455 (.Y (L1_4_L2_2_G4_MINI_ALU_nx454), .A0 (
         L1_4_L2_2_G4_MINI_ALU_BoothOperand_16), .A1 (
         L1_4_L2_2_G4_MINI_ALU_BoothP_16)) ;
    mux21_ni L1_4_L2_2_G4_MINI_ALU_ix91 (.Y (L1FirstOperands_3__0), .A0 (
             L1_4_L2_2_G4_MINI_ALU_BoothP_1), .A1 (WindowDin_4__2__0), .S0 (
             Instr)) ;
    mux21_ni L1_4_L2_2_G4_MINI_ALU_ix99 (.Y (L1FirstOperands_3__1), .A0 (
             L1_4_L2_2_G4_MINI_ALU_BoothP_2), .A1 (WindowDin_4__2__1), .S0 (
             Instr)) ;
    mux21_ni L1_4_L2_2_G4_MINI_ALU_ix107 (.Y (L1FirstOperands_3__2), .A0 (
             L1_4_L2_2_G4_MINI_ALU_BoothP_3), .A1 (WindowDin_4__2__2), .S0 (
             Instr)) ;
    mux21_ni L1_4_L2_2_G4_MINI_ALU_ix115 (.Y (L1FirstOperands_3__3), .A0 (
             L1_4_L2_2_G4_MINI_ALU_BoothP_4), .A1 (WindowDin_4__2__3), .S0 (
             Instr)) ;
    mux21_ni L1_4_L2_2_G4_MINI_ALU_ix123 (.Y (L1FirstOperands_3__4), .A0 (
             L1_4_L2_2_G4_MINI_ALU_BoothP_5), .A1 (WindowDin_4__2__4), .S0 (
             Instr)) ;
    mux21_ni L1_4_L2_2_G4_MINI_ALU_ix131 (.Y (L1FirstOperands_3__5), .A0 (
             L1_4_L2_2_G4_MINI_ALU_BoothP_6), .A1 (WindowDin_4__2__5), .S0 (
             Instr)) ;
    mux21_ni L1_4_L2_2_G4_MINI_ALU_ix139 (.Y (L1FirstOperands_3__6), .A0 (
             L1_4_L2_2_G4_MINI_ALU_BoothP_7), .A1 (WindowDin_4__2__6), .S0 (
             Instr)) ;
    mux21_ni L1_4_L2_2_G4_MINI_ALU_ix147 (.Y (L1FirstOperands_3__7), .A0 (
             L1_4_L2_2_G4_MINI_ALU_BoothP_8), .A1 (WindowDin_4__2__7), .S0 (
             Instr)) ;
    xor2 L1_4_L2_2_G4_MINI_ALU_ix77 (.Y (L4Results_0__1), .A0 (
         L1_4_L2_2_G4_MINI_ALU_nx529), .A1 (L1_4_L2_2_G4_MINI_ALU_nx531)) ;
    nand02 L1_4_L2_2_G4_MINI_ALU_ix530 (.Y (L1_4_L2_2_G4_MINI_ALU_nx529), .A0 (
           L3Results_1__0), .A1 (L3Results_0__0)) ;
    xnor2 L1_4_L2_2_G4_MINI_ALU_ix532 (.Y (L1_4_L2_2_G4_MINI_ALU_nx531), .A0 (
          L3Results_1__1), .A1 (L3Results_0__1)) ;
    xor2 L1_4_L2_2_G4_MINI_ALU_ix75 (.Y (L4Results_0__2), .A0 (
         L1_4_L2_2_G4_MINI_ALU_nx534), .A1 (L1_4_L2_2_G4_MINI_ALU_nx537)) ;
    aoi32 L1_4_L2_2_G4_MINI_ALU_ix535 (.Y (L1_4_L2_2_G4_MINI_ALU_nx534), .A0 (
          L3Results_1__0), .A1 (L3Results_0__0), .A2 (L1_4_L2_2_G4_MINI_ALU_nx30
          ), .B0 (L3Results_0__1), .B1 (L3Results_1__1)) ;
    xnor2 L1_4_L2_2_G4_MINI_ALU_ix538 (.Y (L1_4_L2_2_G4_MINI_ALU_nx537), .A0 (
          L3Results_1__2), .A1 (L3Results_0__2)) ;
    xor2 L1_4_L2_2_G4_MINI_ALU_ix73 (.Y (L4Results_0__3), .A0 (
         L1_4_L2_2_G4_MINI_ALU_nx540), .A1 (L1_4_L2_2_G4_MINI_ALU_nx544)) ;
    aoi22 L1_4_L2_2_G4_MINI_ALU_ix541 (.Y (L1_4_L2_2_G4_MINI_ALU_nx540), .A0 (
          L3Results_0__2), .A1 (L3Results_1__2), .B0 (L1_4_L2_2_G4_MINI_ALU_nx40
          ), .B1 (L1_4_L2_2_G4_MINI_ALU_nx24)) ;
    xnor2 L1_4_L2_2_G4_MINI_ALU_ix545 (.Y (L1_4_L2_2_G4_MINI_ALU_nx544), .A0 (
          L3Results_1__3), .A1 (L3Results_0__3)) ;
    xor2 L1_4_L2_2_G4_MINI_ALU_ix71 (.Y (L4Results_0__4), .A0 (
         L1_4_L2_2_G4_MINI_ALU_nx547), .A1 (L1_4_L2_2_G4_MINI_ALU_nx551)) ;
    aoi22 L1_4_L2_2_G4_MINI_ALU_ix548 (.Y (L1_4_L2_2_G4_MINI_ALU_nx547), .A0 (
          L3Results_0__3), .A1 (L3Results_1__3), .B0 (L1_4_L2_2_G4_MINI_ALU_nx44
          ), .B1 (L1_4_L2_2_G4_MINI_ALU_nx18)) ;
    xnor2 L1_4_L2_2_G4_MINI_ALU_ix552 (.Y (L1_4_L2_2_G4_MINI_ALU_nx551), .A0 (
          L3Results_1__4), .A1 (L3Results_0__4)) ;
    xor2 L1_4_L2_2_G4_MINI_ALU_ix69 (.Y (L4Results_0__5), .A0 (
         L1_4_L2_2_G4_MINI_ALU_nx554), .A1 (L1_4_L2_2_G4_MINI_ALU_nx558)) ;
    aoi22 L1_4_L2_2_G4_MINI_ALU_ix555 (.Y (L1_4_L2_2_G4_MINI_ALU_nx554), .A0 (
          L3Results_0__4), .A1 (L3Results_1__4), .B0 (L1_4_L2_2_G4_MINI_ALU_nx48
          ), .B1 (L1_4_L2_2_G4_MINI_ALU_nx12)) ;
    xnor2 L1_4_L2_2_G4_MINI_ALU_ix559 (.Y (L1_4_L2_2_G4_MINI_ALU_nx558), .A0 (
          L3Results_1__5), .A1 (L3Results_0__5)) ;
    xor2 L1_4_L2_2_G4_MINI_ALU_ix67 (.Y (L4Results_0__6), .A0 (
         L1_4_L2_2_G4_MINI_ALU_nx561), .A1 (L1_4_L2_2_G4_MINI_ALU_nx565)) ;
    aoi22 L1_4_L2_2_G4_MINI_ALU_ix562 (.Y (L1_4_L2_2_G4_MINI_ALU_nx561), .A0 (
          L3Results_0__5), .A1 (L3Results_1__5), .B0 (L1_4_L2_2_G4_MINI_ALU_nx52
          ), .B1 (L1_4_L2_2_G4_MINI_ALU_nx6)) ;
    xnor2 L1_4_L2_2_G4_MINI_ALU_ix566 (.Y (L1_4_L2_2_G4_MINI_ALU_nx565), .A0 (
          L3Results_1__6), .A1 (L3Results_0__6)) ;
    xnor2 L1_4_L2_2_G4_MINI_ALU_ix65 (.Y (L4Results_0__7), .A0 (
          L1_4_L2_2_G4_MINI_ALU_nx568), .A1 (L1_4_L2_2_G4_MINI_ALU_nx62)) ;
    aoi22 L1_4_L2_2_G4_MINI_ALU_ix569 (.Y (L1_4_L2_2_G4_MINI_ALU_nx568), .A0 (
          L3Results_0__6), .A1 (L3Results_1__6), .B0 (L1_4_L2_2_G4_MINI_ALU_nx56
          ), .B1 (L1_4_L2_2_G4_MINI_ALU_nx0)) ;
    xor2 L1_4_L2_2_G4_MINI_ALU_ix63 (.Y (L1_4_L2_2_G4_MINI_ALU_nx62), .A0 (
         L3Results_1__7), .A1 (L3Results_0__7)) ;
    inv01 L1_4_L2_2_G4_MINI_ALU_ix155 (.Y (L1_4_L2_2_G4_MINI_ALU_nx154), .A (
          L1_4_L2_2_G4_MINI_ALU_nx383)) ;
    inv01 L1_4_L2_2_G4_MINI_ALU_ix57 (.Y (L1_4_L2_2_G4_MINI_ALU_nx56), .A (
          L1_4_L2_2_G4_MINI_ALU_nx561)) ;
    inv01 L1_4_L2_2_G4_MINI_ALU_ix53 (.Y (L1_4_L2_2_G4_MINI_ALU_nx52), .A (
          L1_4_L2_2_G4_MINI_ALU_nx554)) ;
    inv01 L1_4_L2_2_G4_MINI_ALU_ix49 (.Y (L1_4_L2_2_G4_MINI_ALU_nx48), .A (
          L1_4_L2_2_G4_MINI_ALU_nx547)) ;
    inv01 L1_4_L2_2_G4_MINI_ALU_ix45 (.Y (L1_4_L2_2_G4_MINI_ALU_nx44), .A (
          L1_4_L2_2_G4_MINI_ALU_nx540)) ;
    inv01 L1_4_L2_2_G4_MINI_ALU_ix41 (.Y (L1_4_L2_2_G4_MINI_ALU_nx40), .A (
          L1_4_L2_2_G4_MINI_ALU_nx534)) ;
    inv01 L1_4_L2_2_G4_MINI_ALU_ix31 (.Y (L1_4_L2_2_G4_MINI_ALU_nx30), .A (
          L1_4_L2_2_G4_MINI_ALU_nx531)) ;
    inv01 L1_4_L2_2_G4_MINI_ALU_ix25 (.Y (L1_4_L2_2_G4_MINI_ALU_nx24), .A (
          L1_4_L2_2_G4_MINI_ALU_nx537)) ;
    inv01 L1_4_L2_2_G4_MINI_ALU_ix19 (.Y (L1_4_L2_2_G4_MINI_ALU_nx18), .A (
          L1_4_L2_2_G4_MINI_ALU_nx544)) ;
    inv01 L1_4_L2_2_G4_MINI_ALU_ix13 (.Y (L1_4_L2_2_G4_MINI_ALU_nx12), .A (
          L1_4_L2_2_G4_MINI_ALU_nx551)) ;
    inv01 L1_4_L2_2_G4_MINI_ALU_ix7 (.Y (L1_4_L2_2_G4_MINI_ALU_nx6), .A (
          L1_4_L2_2_G4_MINI_ALU_nx558)) ;
    inv01 L1_4_L2_2_G4_MINI_ALU_ix1 (.Y (L1_4_L2_2_G4_MINI_ALU_nx0), .A (
          L1_4_L2_2_G4_MINI_ALU_nx565)) ;
    fake_gnd L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix216 (.Y (
             L1_4_L2_2_G4_MINI_ALU_WindowCellShiftedLeft_16)) ;
    nor02ii L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix81 (.Y (
            L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_nx80), .A0 (Instr), .A1 (Start)) ;
    aoi21 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix77 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDin_10), .A0 (
          FilterDin_4__2__1), .A1 (FilterDin_4__2__0), .B0 (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_nx4)) ;
    nor02_2x L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix5 (.Y (
             L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_nx4), .A0 (FilterDin_4__2__0), .A1 (
             FilterDin_4__2__1)) ;
    aoi21 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix67 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDin_11), .A0 (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_nx328), .A1 (FilterDin_4__2__2), .B0 (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_nx8)) ;
    nor03_2x L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix9 (.Y (
             L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_nx8), .A0 (FilterDin_4__2__2), .A1 (
             FilterDin_4__2__0), .A2 (FilterDin_4__2__1)) ;
    xnor2 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix59 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDin_12), .A0 (
          FilterDin_4__2__3), .A1 (L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_nx8)) ;
    xnor2 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix51 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDin_13), .A0 (
          FilterDin_4__2__4), .A1 (L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_nx12)) ;
    nor04 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix13 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_nx12), .A0 (FilterDin_4__2__3), .A1 (
          FilterDin_4__2__2), .A2 (FilterDin_4__2__0), .A3 (FilterDin_4__2__1)
          ) ;
    xnor2 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix43 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDin_14), .A0 (
          FilterDin_4__2__5), .A1 (L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_nx16)) ;
    nor02ii L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix17 (.Y (
            L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_nx16), .A0 (FilterDin_4__2__4), .A1 (
            L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_nx12)) ;
    xnor2 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix35 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDin_15), .A0 (
          FilterDin_4__2__6), .A1 (L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_nx20)) ;
    nor02ii L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix21 (.Y (
            L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_nx20), .A0 (FilterDin_4__2__5), .A1 (
            L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_nx16)) ;
    xnor2 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix27 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDin_16), .A0 (
          FilterDin_4__2__7), .A1 (L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_nx24)) ;
    nor02ii L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix25 (.Y (
            L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_nx24), .A0 (FilterDin_4__2__6), .A1 (
            L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_nx20)) ;
    inv01 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix329 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_nx328), .A (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_nx4)) ;
    inv02 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix383 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_nx384), .A (
          L1_4_L2_2_G4_MINI_ALU_BoothP_0)) ;
    dff L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_0 (.Q (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_0), .QB (\$dummy [1126])
        , .D (L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .CLK (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    nor02_2x L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix567 (.Y (
             L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566), .A0 (RST), .A1 (
             L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644)) ;
    dff L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_1 (.Q (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_1), .QB (\$dummy [1127])
        , .D (L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .CLK (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_2 (.Q (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_2), .QB (\$dummy [1128])
        , .D (L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .CLK (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_3 (.Q (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_3), .QB (\$dummy [1129])
        , .D (L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .CLK (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_4 (.Q (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_4), .QB (\$dummy [1130])
        , .D (L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .CLK (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_5 (.Q (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_5), .QB (\$dummy [1131])
        , .D (L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .CLK (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_6 (.Q (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_6), .QB (\$dummy [1132])
        , .D (L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .CLK (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_7 (.Q (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_7), .QB (\$dummy [1133])
        , .D (L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .CLK (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_8 (.Q (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_8), .QB (\$dummy [1134])
        , .D (L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .CLK (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_9 (.Q (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_9), .QB (\$dummy [1135])
        , .D (L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .CLK (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_10 (.Q (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_10), .QB (\$dummy [1136])
        , .D (L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .CLK (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_11 (.Q (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_11), .QB (\$dummy [1137])
        , .D (L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .CLK (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_12 (.Q (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_12), .QB (\$dummy [1138])
        , .D (L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .CLK (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_13 (.Q (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_13), .QB (\$dummy [1139])
        , .D (L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .CLK (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_14 (.Q (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_14), .QB (\$dummy [1140])
        , .D (L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .CLK (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_15 (.Q (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_15), .QB (\$dummy [1141])
        , .D (L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .CLK (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_16 (.Q (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_16), .QB (\$dummy [1142])
        , .D (L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .CLK (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    inv02 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix623 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624), .A (CLK)) ;
    inv02 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix625 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626), .A (CLK)) ;
    inv02 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix627 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628), .A (CLK)) ;
    inv02 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix643 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644), .A (nx8498)) ;
    dff L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_0 (.Q (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_0), .QB (\$dummy [1143])
        , .D (L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .CLK (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    nor02_2x L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix567 (.Y (
             L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566), .A0 (RST), .A1 (
             L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644)) ;
    dff L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_1 (.Q (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_1), .QB (\$dummy [1144])
        , .D (L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .CLK (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_2 (.Q (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_2), .QB (\$dummy [1145])
        , .D (L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .CLK (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_3 (.Q (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_3), .QB (\$dummy [1146])
        , .D (L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .CLK (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_4 (.Q (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_4), .QB (\$dummy [1147])
        , .D (L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .CLK (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_5 (.Q (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_5), .QB (\$dummy [1148])
        , .D (L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .CLK (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_6 (.Q (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_6), .QB (\$dummy [1149])
        , .D (L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .CLK (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_7 (.Q (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_7), .QB (\$dummy [1150])
        , .D (L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .CLK (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_8 (.Q (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_8), .QB (\$dummy [1151])
        , .D (L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .CLK (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_9 (.Q (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_9), .QB (\$dummy [1152])
        , .D (L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .CLK (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_10 (.Q (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_10), .QB (\$dummy [1153])
        , .D (L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .CLK (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_11 (.Q (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_11), .QB (\$dummy [1154])
        , .D (L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .CLK (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_12 (.Q (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_12), .QB (\$dummy [1155])
        , .D (L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .CLK (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_13 (.Q (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_13), .QB (\$dummy [1156])
        , .D (L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .CLK (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_14 (.Q (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_14), .QB (\$dummy [1157])
        , .D (L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .CLK (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_15 (.Q (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_15), .QB (\$dummy [1158])
        , .D (L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .CLK (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_16 (.Q (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_16), .QB (\$dummy [1159])
        , .D (L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .CLK (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    inv02 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix623 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624), .A (CLK)) ;
    inv02 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix625 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626), .A (CLK)) ;
    inv02 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix627 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628), .A (CLK)) ;
    inv02 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix643 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644), .A (nx8504)) ;
    dff L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_0 (.Q (
        L1_4_L2_2_G4_MINI_ALU_BoothP_0), .QB (\$dummy [1160]), .D (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .CLK (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    nor02_2x L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix567 (.Y (
             L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566), .A0 (RST), .A1 (
             L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    dff L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_1 (.Q (
        L1_4_L2_2_G4_MINI_ALU_BoothP_1), .QB (\$dummy [1161]), .D (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .CLK (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_2 (.Q (
        L1_4_L2_2_G4_MINI_ALU_BoothP_2), .QB (\$dummy [1162]), .D (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .CLK (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_3 (.Q (
        L1_4_L2_2_G4_MINI_ALU_BoothP_3), .QB (\$dummy [1163]), .D (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .CLK (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_4 (.Q (
        L1_4_L2_2_G4_MINI_ALU_BoothP_4), .QB (\$dummy [1164]), .D (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .CLK (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_5 (.Q (
        L1_4_L2_2_G4_MINI_ALU_BoothP_5), .QB (\$dummy [1165]), .D (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .CLK (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_6 (.Q (
        L1_4_L2_2_G4_MINI_ALU_BoothP_6), .QB (\$dummy [1166]), .D (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .CLK (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_7 (.Q (
        L1_4_L2_2_G4_MINI_ALU_BoothP_7), .QB (\$dummy [1167]), .D (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .CLK (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_8 (.Q (
        L1_4_L2_2_G4_MINI_ALU_BoothP_8), .QB (\$dummy [1168]), .D (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .CLK (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_9 (.Q (
        L1_4_L2_2_G4_MINI_ALU_BoothP_9), .QB (\$dummy [1169]), .D (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .CLK (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_10 (.Q (
        L1_4_L2_2_G4_MINI_ALU_BoothP_10), .QB (\$dummy [1170]), .D (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .CLK (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_11 (.Q (
        L1_4_L2_2_G4_MINI_ALU_BoothP_11), .QB (\$dummy [1171]), .D (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .CLK (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_12 (.Q (
        L1_4_L2_2_G4_MINI_ALU_BoothP_12), .QB (\$dummy [1172]), .D (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .CLK (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_13 (.Q (
        L1_4_L2_2_G4_MINI_ALU_BoothP_13), .QB (\$dummy [1173]), .D (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .CLK (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_14 (.Q (
        L1_4_L2_2_G4_MINI_ALU_BoothP_14), .QB (\$dummy [1174]), .D (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .CLK (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_15 (.Q (
        L1_4_L2_2_G4_MINI_ALU_BoothP_15), .QB (\$dummy [1175]), .D (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .CLK (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_16 (.Q (
        L1_4_L2_2_G4_MINI_ALU_BoothP_16), .QB (\$dummy [1176]), .D (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .CLK (
        L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    inv02 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix623 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624), .A (CLK)) ;
    inv02 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix625 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626), .A (CLK)) ;
    inv02 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix627 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628), .A (CLK)) ;
    inv02 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix643 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644), .A (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642)) ;
    xor2 L1_4_L2_3_G5_MINI_ALU_ix83 (.Y (L5FirstOperands_1__0), .A0 (
         L3Results_2__0), .A1 (L4Results_0__0)) ;
    xnor2 L1_4_L2_3_G5_MINI_ALU_ix380 (.Y (L1_4_L2_3_G5_MINI_ALU_nx379), .A0 (
          L1_4_L2_3_G5_MINI_ALU_nx381), .A1 (L1_4_L2_3_G5_MINI_ALU_nx383)) ;
    nand02 L1_4_L2_3_G5_MINI_ALU_ix382 (.Y (L1_4_L2_3_G5_MINI_ALU_nx381), .A0 (
           L1_4_L2_3_G5_MINI_ALU_BoothOperand_0), .A1 (nx8524)) ;
    xnor2 L1_4_L2_3_G5_MINI_ALU_ix384 (.Y (L1_4_L2_3_G5_MINI_ALU_nx383), .A0 (
          L1_4_L2_3_G5_MINI_ALU_BoothOperand_1), .A1 (
          L1_4_L2_3_G5_MINI_ALU_BoothP_1)) ;
    inv01 L1_4_L2_3_G5_MINI_ALU_ix388 (.Y (L1_4_L2_3_G5_MINI_ALU_nx387), .A (
          L1_4_L2_3_G5_MINI_ALU_BoothP_2)) ;
    xnor2 L1_4_L2_3_G5_MINI_ALU_ix390 (.Y (L1_4_L2_3_G5_MINI_ALU_nx389), .A0 (
          L1_4_L2_3_G5_MINI_ALU_nx391), .A1 (L1_4_L2_3_G5_MINI_ALU_nx395)) ;
    aoi32 L1_4_L2_3_G5_MINI_ALU_ix392 (.Y (L1_4_L2_3_G5_MINI_ALU_nx391), .A0 (
          L1_4_L2_3_G5_MINI_ALU_BoothOperand_0), .A1 (nx8524), .A2 (
          L1_4_L2_3_G5_MINI_ALU_nx154), .B0 (L1_4_L2_3_G5_MINI_ALU_BoothP_1), .B1 (
          L1_4_L2_3_G5_MINI_ALU_BoothOperand_1)) ;
    xnor2 L1_4_L2_3_G5_MINI_ALU_ix396 (.Y (L1_4_L2_3_G5_MINI_ALU_nx395), .A0 (
          L1_4_L2_3_G5_MINI_ALU_BoothOperand_2), .A1 (
          L1_4_L2_3_G5_MINI_ALU_BoothP_2)) ;
    inv01 L1_4_L2_3_G5_MINI_ALU_ix400 (.Y (L1_4_L2_3_G5_MINI_ALU_nx399), .A (
          L1_4_L2_3_G5_MINI_ALU_BoothP_3)) ;
    xnor2 L1_4_L2_3_G5_MINI_ALU_ix402 (.Y (L1_4_L2_3_G5_MINI_ALU_nx401), .A0 (
          L1_4_L2_3_G5_MINI_ALU_nx403), .A1 (L1_4_L2_3_G5_MINI_ALU_nx405)) ;
    xnor2 L1_4_L2_3_G5_MINI_ALU_ix406 (.Y (L1_4_L2_3_G5_MINI_ALU_nx405), .A0 (
          L1_4_L2_3_G5_MINI_ALU_BoothOperand_3), .A1 (
          L1_4_L2_3_G5_MINI_ALU_BoothP_3)) ;
    inv01 L1_4_L2_3_G5_MINI_ALU_ix410 (.Y (L1_4_L2_3_G5_MINI_ALU_nx409), .A (
          L1_4_L2_3_G5_MINI_ALU_BoothP_4)) ;
    xnor2 L1_4_L2_3_G5_MINI_ALU_ix412 (.Y (L1_4_L2_3_G5_MINI_ALU_nx411), .A0 (
          L1_4_L2_3_G5_MINI_ALU_nx413), .A1 (L1_4_L2_3_G5_MINI_ALU_nx415)) ;
    xnor2 L1_4_L2_3_G5_MINI_ALU_ix416 (.Y (L1_4_L2_3_G5_MINI_ALU_nx415), .A0 (
          L1_4_L2_3_G5_MINI_ALU_BoothOperand_4), .A1 (
          L1_4_L2_3_G5_MINI_ALU_BoothP_4)) ;
    inv01 L1_4_L2_3_G5_MINI_ALU_ix420 (.Y (L1_4_L2_3_G5_MINI_ALU_nx419), .A (
          L1_4_L2_3_G5_MINI_ALU_BoothP_5)) ;
    xnor2 L1_4_L2_3_G5_MINI_ALU_ix422 (.Y (L1_4_L2_3_G5_MINI_ALU_nx421), .A0 (
          L1_4_L2_3_G5_MINI_ALU_nx423), .A1 (L1_4_L2_3_G5_MINI_ALU_nx425)) ;
    xnor2 L1_4_L2_3_G5_MINI_ALU_ix426 (.Y (L1_4_L2_3_G5_MINI_ALU_nx425), .A0 (
          L1_4_L2_3_G5_MINI_ALU_BoothOperand_5), .A1 (
          L1_4_L2_3_G5_MINI_ALU_BoothP_5)) ;
    inv01 L1_4_L2_3_G5_MINI_ALU_ix430 (.Y (L1_4_L2_3_G5_MINI_ALU_nx429), .A (
          L1_4_L2_3_G5_MINI_ALU_BoothP_6)) ;
    xnor2 L1_4_L2_3_G5_MINI_ALU_ix432 (.Y (L1_4_L2_3_G5_MINI_ALU_nx431), .A0 (
          L1_4_L2_3_G5_MINI_ALU_nx433), .A1 (L1_4_L2_3_G5_MINI_ALU_nx435)) ;
    xnor2 L1_4_L2_3_G5_MINI_ALU_ix436 (.Y (L1_4_L2_3_G5_MINI_ALU_nx435), .A0 (
          L1_4_L2_3_G5_MINI_ALU_BoothOperand_6), .A1 (
          L1_4_L2_3_G5_MINI_ALU_BoothP_6)) ;
    inv01 L1_4_L2_3_G5_MINI_ALU_ix440 (.Y (L1_4_L2_3_G5_MINI_ALU_nx439), .A (
          L1_4_L2_3_G5_MINI_ALU_BoothP_7)) ;
    xnor2 L1_4_L2_3_G5_MINI_ALU_ix442 (.Y (L1_4_L2_3_G5_MINI_ALU_nx441), .A0 (
          L1_4_L2_3_G5_MINI_ALU_nx443), .A1 (L1_4_L2_3_G5_MINI_ALU_nx445)) ;
    xnor2 L1_4_L2_3_G5_MINI_ALU_ix446 (.Y (L1_4_L2_3_G5_MINI_ALU_nx445), .A0 (
          L1_4_L2_3_G5_MINI_ALU_BoothOperand_7), .A1 (
          L1_4_L2_3_G5_MINI_ALU_BoothP_7)) ;
    inv01 L1_4_L2_3_G5_MINI_ALU_ix450 (.Y (L1_4_L2_3_G5_MINI_ALU_nx449), .A (
          L1_4_L2_3_G5_MINI_ALU_BoothP_8)) ;
    xnor2 L1_4_L2_3_G5_MINI_ALU_ix452 (.Y (L1_4_L2_3_G5_MINI_ALU_nx451), .A0 (
          L1_4_L2_3_G5_MINI_ALU_nx453), .A1 (L1_4_L2_3_G5_MINI_ALU_nx455)) ;
    xnor2 L1_4_L2_3_G5_MINI_ALU_ix456 (.Y (L1_4_L2_3_G5_MINI_ALU_nx455), .A0 (
          L1_4_L2_3_G5_MINI_ALU_BoothOperand_8), .A1 (
          L1_4_L2_3_G5_MINI_ALU_BoothP_8)) ;
    xor2 L1_4_L2_3_G5_MINI_ALU_ix317 (.Y (L1_4_L2_3_G5_MINI_ALU_nx316), .A0 (
         L1_4_L2_3_G5_MINI_ALU_nx461), .A1 (L1_4_L2_3_G5_MINI_ALU_nx463)) ;
    xnor2 L1_4_L2_3_G5_MINI_ALU_ix464 (.Y (L1_4_L2_3_G5_MINI_ALU_nx463), .A0 (
          L1_4_L2_3_G5_MINI_ALU_BoothOperand_9), .A1 (
          L1_4_L2_3_G5_MINI_ALU_BoothP_9)) ;
    xor2 L1_4_L2_3_G5_MINI_ALU_ix337 (.Y (L1_4_L2_3_G5_MINI_ALU_nx336), .A0 (
         L1_4_L2_3_G5_MINI_ALU_nx467), .A1 (L1_4_L2_3_G5_MINI_ALU_nx471)) ;
    inv01 L1_4_L2_3_G5_MINI_ALU_ix470 (.Y (L1_4_L2_3_G5_MINI_ALU_nx469), .A (
          L1_4_L2_3_G5_MINI_ALU_BoothP_9)) ;
    xnor2 L1_4_L2_3_G5_MINI_ALU_ix472 (.Y (L1_4_L2_3_G5_MINI_ALU_nx471), .A0 (
          L1_4_L2_3_G5_MINI_ALU_BoothOperand_10), .A1 (
          L1_4_L2_3_G5_MINI_ALU_BoothP_10)) ;
    xor2 L1_4_L2_3_G5_MINI_ALU_ix357 (.Y (L1_4_L2_3_G5_MINI_ALU_nx356), .A0 (
         L1_4_L2_3_G5_MINI_ALU_nx475), .A1 (L1_4_L2_3_G5_MINI_ALU_nx479)) ;
    inv01 L1_4_L2_3_G5_MINI_ALU_ix478 (.Y (L1_4_L2_3_G5_MINI_ALU_nx477), .A (
          L1_4_L2_3_G5_MINI_ALU_BoothP_10)) ;
    xnor2 L1_4_L2_3_G5_MINI_ALU_ix480 (.Y (L1_4_L2_3_G5_MINI_ALU_nx479), .A0 (
          L1_4_L2_3_G5_MINI_ALU_BoothOperand_11), .A1 (
          L1_4_L2_3_G5_MINI_ALU_BoothP_11)) ;
    xor2 L1_4_L2_3_G5_MINI_ALU_ix377 (.Y (L1_4_L2_3_G5_MINI_ALU_nx376), .A0 (
         L1_4_L2_3_G5_MINI_ALU_nx483), .A1 (L1_4_L2_3_G5_MINI_ALU_nx487)) ;
    inv01 L1_4_L2_3_G5_MINI_ALU_ix486 (.Y (L1_4_L2_3_G5_MINI_ALU_nx485), .A (
          L1_4_L2_3_G5_MINI_ALU_BoothP_11)) ;
    xnor2 L1_4_L2_3_G5_MINI_ALU_ix488 (.Y (L1_4_L2_3_G5_MINI_ALU_nx487), .A0 (
          L1_4_L2_3_G5_MINI_ALU_BoothOperand_12), .A1 (
          L1_4_L2_3_G5_MINI_ALU_BoothP_12)) ;
    xor2 L1_4_L2_3_G5_MINI_ALU_ix397 (.Y (L1_4_L2_3_G5_MINI_ALU_nx396), .A0 (
         L1_4_L2_3_G5_MINI_ALU_nx491), .A1 (L1_4_L2_3_G5_MINI_ALU_nx495)) ;
    inv01 L1_4_L2_3_G5_MINI_ALU_ix494 (.Y (L1_4_L2_3_G5_MINI_ALU_nx493), .A (
          L1_4_L2_3_G5_MINI_ALU_BoothP_12)) ;
    xnor2 L1_4_L2_3_G5_MINI_ALU_ix496 (.Y (L1_4_L2_3_G5_MINI_ALU_nx495), .A0 (
          L1_4_L2_3_G5_MINI_ALU_BoothOperand_13), .A1 (
          L1_4_L2_3_G5_MINI_ALU_BoothP_13)) ;
    xor2 L1_4_L2_3_G5_MINI_ALU_ix417 (.Y (L1_4_L2_3_G5_MINI_ALU_nx416), .A0 (
         L1_4_L2_3_G5_MINI_ALU_nx499), .A1 (L1_4_L2_3_G5_MINI_ALU_nx503)) ;
    inv01 L1_4_L2_3_G5_MINI_ALU_ix502 (.Y (L1_4_L2_3_G5_MINI_ALU_nx501), .A (
          L1_4_L2_3_G5_MINI_ALU_BoothP_13)) ;
    xnor2 L1_4_L2_3_G5_MINI_ALU_ix504 (.Y (L1_4_L2_3_G5_MINI_ALU_nx503), .A0 (
          L1_4_L2_3_G5_MINI_ALU_BoothOperand_14), .A1 (
          L1_4_L2_3_G5_MINI_ALU_BoothP_14)) ;
    xor2 L1_4_L2_3_G5_MINI_ALU_ix437 (.Y (L1_4_L2_3_G5_MINI_ALU_nx436), .A0 (
         L1_4_L2_3_G5_MINI_ALU_nx507), .A1 (L1_4_L2_3_G5_MINI_ALU_nx511)) ;
    inv01 L1_4_L2_3_G5_MINI_ALU_ix510 (.Y (L1_4_L2_3_G5_MINI_ALU_nx509), .A (
          L1_4_L2_3_G5_MINI_ALU_BoothP_14)) ;
    xnor2 L1_4_L2_3_G5_MINI_ALU_ix512 (.Y (L1_4_L2_3_G5_MINI_ALU_nx511), .A0 (
          L1_4_L2_3_G5_MINI_ALU_BoothOperand_15), .A1 (
          L1_4_L2_3_G5_MINI_ALU_BoothP_15)) ;
    xnor2 L1_4_L2_3_G5_MINI_ALU_ix457 (.Y (L1_4_L2_3_G5_MINI_ALU_nx456), .A0 (
          L1_4_L2_3_G5_MINI_ALU_nx515), .A1 (L1_4_L2_3_G5_MINI_ALU_nx454)) ;
    inv01 L1_4_L2_3_G5_MINI_ALU_ix518 (.Y (L1_4_L2_3_G5_MINI_ALU_nx517), .A (
          L1_4_L2_3_G5_MINI_ALU_BoothP_15)) ;
    xor2 L1_4_L2_3_G5_MINI_ALU_ix455 (.Y (L1_4_L2_3_G5_MINI_ALU_nx454), .A0 (
         L1_4_L2_3_G5_MINI_ALU_BoothOperand_16), .A1 (
         L1_4_L2_3_G5_MINI_ALU_BoothP_16)) ;
    mux21_ni L1_4_L2_3_G5_MINI_ALU_ix91 (.Y (L1FirstOperands_7__0), .A0 (
             L1_4_L2_3_G5_MINI_ALU_BoothP_1), .A1 (WindowDin_4__3__0), .S0 (
             Instr)) ;
    mux21_ni L1_4_L2_3_G5_MINI_ALU_ix99 (.Y (L1FirstOperands_7__1), .A0 (
             L1_4_L2_3_G5_MINI_ALU_BoothP_2), .A1 (WindowDin_4__3__1), .S0 (
             Instr)) ;
    mux21_ni L1_4_L2_3_G5_MINI_ALU_ix107 (.Y (L1FirstOperands_7__2), .A0 (
             L1_4_L2_3_G5_MINI_ALU_BoothP_3), .A1 (WindowDin_4__3__2), .S0 (
             Instr)) ;
    mux21_ni L1_4_L2_3_G5_MINI_ALU_ix115 (.Y (L1FirstOperands_7__3), .A0 (
             L1_4_L2_3_G5_MINI_ALU_BoothP_4), .A1 (WindowDin_4__3__3), .S0 (
             Instr)) ;
    mux21_ni L1_4_L2_3_G5_MINI_ALU_ix123 (.Y (L1FirstOperands_7__4), .A0 (
             L1_4_L2_3_G5_MINI_ALU_BoothP_5), .A1 (WindowDin_4__3__4), .S0 (
             Instr)) ;
    mux21_ni L1_4_L2_3_G5_MINI_ALU_ix131 (.Y (L1FirstOperands_7__5), .A0 (
             L1_4_L2_3_G5_MINI_ALU_BoothP_6), .A1 (WindowDin_4__3__5), .S0 (
             Instr)) ;
    mux21_ni L1_4_L2_3_G5_MINI_ALU_ix139 (.Y (L1FirstOperands_7__6), .A0 (
             L1_4_L2_3_G5_MINI_ALU_BoothP_7), .A1 (WindowDin_4__3__6), .S0 (
             Instr)) ;
    mux21_ni L1_4_L2_3_G5_MINI_ALU_ix147 (.Y (L1FirstOperands_7__7), .A0 (
             L1_4_L2_3_G5_MINI_ALU_BoothP_8), .A1 (WindowDin_4__3__7), .S0 (
             Instr)) ;
    xor2 L1_4_L2_3_G5_MINI_ALU_ix77 (.Y (L5FirstOperands_1__1), .A0 (
         L1_4_L2_3_G5_MINI_ALU_nx529), .A1 (L1_4_L2_3_G5_MINI_ALU_nx531)) ;
    nand02 L1_4_L2_3_G5_MINI_ALU_ix530 (.Y (L1_4_L2_3_G5_MINI_ALU_nx529), .A0 (
           L3Results_2__0), .A1 (L4Results_0__0)) ;
    xnor2 L1_4_L2_3_G5_MINI_ALU_ix532 (.Y (L1_4_L2_3_G5_MINI_ALU_nx531), .A0 (
          L3Results_2__1), .A1 (L4Results_0__1)) ;
    xor2 L1_4_L2_3_G5_MINI_ALU_ix75 (.Y (L5FirstOperands_1__2), .A0 (
         L1_4_L2_3_G5_MINI_ALU_nx534), .A1 (L1_4_L2_3_G5_MINI_ALU_nx537)) ;
    aoi32 L1_4_L2_3_G5_MINI_ALU_ix535 (.Y (L1_4_L2_3_G5_MINI_ALU_nx534), .A0 (
          L3Results_2__0), .A1 (L4Results_0__0), .A2 (L1_4_L2_3_G5_MINI_ALU_nx30
          ), .B0 (L4Results_0__1), .B1 (L3Results_2__1)) ;
    xnor2 L1_4_L2_3_G5_MINI_ALU_ix538 (.Y (L1_4_L2_3_G5_MINI_ALU_nx537), .A0 (
          L3Results_2__2), .A1 (L4Results_0__2)) ;
    xor2 L1_4_L2_3_G5_MINI_ALU_ix73 (.Y (L5FirstOperands_1__3), .A0 (
         L1_4_L2_3_G5_MINI_ALU_nx540), .A1 (L1_4_L2_3_G5_MINI_ALU_nx544)) ;
    aoi22 L1_4_L2_3_G5_MINI_ALU_ix541 (.Y (L1_4_L2_3_G5_MINI_ALU_nx540), .A0 (
          L4Results_0__2), .A1 (L3Results_2__2), .B0 (L1_4_L2_3_G5_MINI_ALU_nx40
          ), .B1 (L1_4_L2_3_G5_MINI_ALU_nx24)) ;
    xnor2 L1_4_L2_3_G5_MINI_ALU_ix545 (.Y (L1_4_L2_3_G5_MINI_ALU_nx544), .A0 (
          L3Results_2__3), .A1 (L4Results_0__3)) ;
    xor2 L1_4_L2_3_G5_MINI_ALU_ix71 (.Y (L5FirstOperands_1__4), .A0 (
         L1_4_L2_3_G5_MINI_ALU_nx547), .A1 (L1_4_L2_3_G5_MINI_ALU_nx551)) ;
    aoi22 L1_4_L2_3_G5_MINI_ALU_ix548 (.Y (L1_4_L2_3_G5_MINI_ALU_nx547), .A0 (
          L4Results_0__3), .A1 (L3Results_2__3), .B0 (L1_4_L2_3_G5_MINI_ALU_nx44
          ), .B1 (L1_4_L2_3_G5_MINI_ALU_nx18)) ;
    xnor2 L1_4_L2_3_G5_MINI_ALU_ix552 (.Y (L1_4_L2_3_G5_MINI_ALU_nx551), .A0 (
          L3Results_2__4), .A1 (L4Results_0__4)) ;
    xor2 L1_4_L2_3_G5_MINI_ALU_ix69 (.Y (L5FirstOperands_1__5), .A0 (
         L1_4_L2_3_G5_MINI_ALU_nx554), .A1 (L1_4_L2_3_G5_MINI_ALU_nx558)) ;
    aoi22 L1_4_L2_3_G5_MINI_ALU_ix555 (.Y (L1_4_L2_3_G5_MINI_ALU_nx554), .A0 (
          L4Results_0__4), .A1 (L3Results_2__4), .B0 (L1_4_L2_3_G5_MINI_ALU_nx48
          ), .B1 (L1_4_L2_3_G5_MINI_ALU_nx12)) ;
    xnor2 L1_4_L2_3_G5_MINI_ALU_ix559 (.Y (L1_4_L2_3_G5_MINI_ALU_nx558), .A0 (
          L3Results_2__5), .A1 (L4Results_0__5)) ;
    xor2 L1_4_L2_3_G5_MINI_ALU_ix67 (.Y (L5FirstOperands_1__6), .A0 (
         L1_4_L2_3_G5_MINI_ALU_nx561), .A1 (L1_4_L2_3_G5_MINI_ALU_nx565)) ;
    aoi22 L1_4_L2_3_G5_MINI_ALU_ix562 (.Y (L1_4_L2_3_G5_MINI_ALU_nx561), .A0 (
          L4Results_0__5), .A1 (L3Results_2__5), .B0 (L1_4_L2_3_G5_MINI_ALU_nx52
          ), .B1 (L1_4_L2_3_G5_MINI_ALU_nx6)) ;
    xnor2 L1_4_L2_3_G5_MINI_ALU_ix566 (.Y (L1_4_L2_3_G5_MINI_ALU_nx565), .A0 (
          L3Results_2__6), .A1 (L4Results_0__6)) ;
    xnor2 L1_4_L2_3_G5_MINI_ALU_ix65 (.Y (L5FirstOperands_1__7), .A0 (
          L1_4_L2_3_G5_MINI_ALU_nx568), .A1 (L1_4_L2_3_G5_MINI_ALU_nx62)) ;
    aoi22 L1_4_L2_3_G5_MINI_ALU_ix569 (.Y (L1_4_L2_3_G5_MINI_ALU_nx568), .A0 (
          L4Results_0__6), .A1 (L3Results_2__6), .B0 (L1_4_L2_3_G5_MINI_ALU_nx56
          ), .B1 (L1_4_L2_3_G5_MINI_ALU_nx0)) ;
    xor2 L1_4_L2_3_G5_MINI_ALU_ix63 (.Y (L1_4_L2_3_G5_MINI_ALU_nx62), .A0 (
         L3Results_2__7), .A1 (L4Results_0__7)) ;
    inv01 L1_4_L2_3_G5_MINI_ALU_ix155 (.Y (L1_4_L2_3_G5_MINI_ALU_nx154), .A (
          L1_4_L2_3_G5_MINI_ALU_nx383)) ;
    inv01 L1_4_L2_3_G5_MINI_ALU_ix57 (.Y (L1_4_L2_3_G5_MINI_ALU_nx56), .A (
          L1_4_L2_3_G5_MINI_ALU_nx561)) ;
    inv01 L1_4_L2_3_G5_MINI_ALU_ix53 (.Y (L1_4_L2_3_G5_MINI_ALU_nx52), .A (
          L1_4_L2_3_G5_MINI_ALU_nx554)) ;
    inv01 L1_4_L2_3_G5_MINI_ALU_ix49 (.Y (L1_4_L2_3_G5_MINI_ALU_nx48), .A (
          L1_4_L2_3_G5_MINI_ALU_nx547)) ;
    inv01 L1_4_L2_3_G5_MINI_ALU_ix45 (.Y (L1_4_L2_3_G5_MINI_ALU_nx44), .A (
          L1_4_L2_3_G5_MINI_ALU_nx540)) ;
    inv01 L1_4_L2_3_G5_MINI_ALU_ix41 (.Y (L1_4_L2_3_G5_MINI_ALU_nx40), .A (
          L1_4_L2_3_G5_MINI_ALU_nx534)) ;
    inv01 L1_4_L2_3_G5_MINI_ALU_ix31 (.Y (L1_4_L2_3_G5_MINI_ALU_nx30), .A (
          L1_4_L2_3_G5_MINI_ALU_nx531)) ;
    inv01 L1_4_L2_3_G5_MINI_ALU_ix25 (.Y (L1_4_L2_3_G5_MINI_ALU_nx24), .A (
          L1_4_L2_3_G5_MINI_ALU_nx537)) ;
    inv01 L1_4_L2_3_G5_MINI_ALU_ix19 (.Y (L1_4_L2_3_G5_MINI_ALU_nx18), .A (
          L1_4_L2_3_G5_MINI_ALU_nx544)) ;
    inv01 L1_4_L2_3_G5_MINI_ALU_ix13 (.Y (L1_4_L2_3_G5_MINI_ALU_nx12), .A (
          L1_4_L2_3_G5_MINI_ALU_nx551)) ;
    inv01 L1_4_L2_3_G5_MINI_ALU_ix7 (.Y (L1_4_L2_3_G5_MINI_ALU_nx6), .A (
          L1_4_L2_3_G5_MINI_ALU_nx558)) ;
    inv01 L1_4_L2_3_G5_MINI_ALU_ix1 (.Y (L1_4_L2_3_G5_MINI_ALU_nx0), .A (
          L1_4_L2_3_G5_MINI_ALU_nx565)) ;
    fake_gnd L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix216 (.Y (
             L1_4_L2_3_G5_MINI_ALU_WindowCellShiftedLeft_16)) ;
    nor02ii L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix81 (.Y (
            L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_nx80), .A0 (Instr), .A1 (Start)) ;
    aoi21 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix77 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_10), .A0 (
          FilterDin_4__3__1), .A1 (FilterDin_4__3__0), .B0 (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_nx4)) ;
    nor02_2x L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix5 (.Y (
             L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_nx4), .A0 (FilterDin_4__3__0), .A1 (
             FilterDin_4__3__1)) ;
    aoi21 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix67 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_11), .A0 (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_nx328), .A1 (FilterDin_4__3__2), .B0 (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_nx8)) ;
    nor03_2x L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix9 (.Y (
             L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_nx8), .A0 (FilterDin_4__3__2), .A1 (
             FilterDin_4__3__0), .A2 (FilterDin_4__3__1)) ;
    xnor2 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix59 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_12), .A0 (
          FilterDin_4__3__3), .A1 (L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_nx8)) ;
    xnor2 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix51 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_13), .A0 (
          FilterDin_4__3__4), .A1 (L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_nx12)) ;
    nor04 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix13 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_nx12), .A0 (FilterDin_4__3__3), .A1 (
          FilterDin_4__3__2), .A2 (FilterDin_4__3__0), .A3 (FilterDin_4__3__1)
          ) ;
    xnor2 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix43 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_14), .A0 (
          FilterDin_4__3__5), .A1 (L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_nx16)) ;
    nor02ii L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix17 (.Y (
            L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_nx16), .A0 (FilterDin_4__3__4), .A1 (
            L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_nx12)) ;
    xnor2 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix35 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_15), .A0 (
          FilterDin_4__3__6), .A1 (L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_nx20)) ;
    nor02ii L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix21 (.Y (
            L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_nx20), .A0 (FilterDin_4__3__5), .A1 (
            L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_nx16)) ;
    xnor2 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix27 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_16), .A0 (
          FilterDin_4__3__7), .A1 (L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_nx24)) ;
    nor02ii L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix25 (.Y (
            L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_nx24), .A0 (FilterDin_4__3__6), .A1 (
            L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_nx20)) ;
    inv01 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix329 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_nx328), .A (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_nx4)) ;
    inv02 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix383 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_nx384), .A (
          L1_4_L2_3_G5_MINI_ALU_BoothP_0)) ;
    dff L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_0 (.Q (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_0), .QB (\$dummy [1177])
        , .D (L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .CLK (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    nor02_2x L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix567 (.Y (
             L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566), .A0 (RST), .A1 (
             L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644)) ;
    dff L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_1 (.Q (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_1), .QB (\$dummy [1178])
        , .D (L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .CLK (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_2 (.Q (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_2), .QB (\$dummy [1179])
        , .D (L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .CLK (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_3 (.Q (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_3), .QB (\$dummy [1180])
        , .D (L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .CLK (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_4 (.Q (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_4), .QB (\$dummy [1181])
        , .D (L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .CLK (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_5 (.Q (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_5), .QB (\$dummy [1182])
        , .D (L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .CLK (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_6 (.Q (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_6), .QB (\$dummy [1183])
        , .D (L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .CLK (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_7 (.Q (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_7), .QB (\$dummy [1184])
        , .D (L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .CLK (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_8 (.Q (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_8), .QB (\$dummy [1185])
        , .D (L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .CLK (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_9 (.Q (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_9), .QB (\$dummy [1186])
        , .D (L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .CLK (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_10 (.Q (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_10), .QB (\$dummy [1187])
        , .D (L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .CLK (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_11 (.Q (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_11), .QB (\$dummy [1188])
        , .D (L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .CLK (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_12 (.Q (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_12), .QB (\$dummy [1189])
        , .D (L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .CLK (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_13 (.Q (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_13), .QB (\$dummy [1190])
        , .D (L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .CLK (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_14 (.Q (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_14), .QB (\$dummy [1191])
        , .D (L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .CLK (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_15 (.Q (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_15), .QB (\$dummy [1192])
        , .D (L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .CLK (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_16 (.Q (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_16), .QB (\$dummy [1193])
        , .D (L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .CLK (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    inv02 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix623 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624), .A (CLK)) ;
    inv02 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix625 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626), .A (CLK)) ;
    inv02 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix627 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628), .A (CLK)) ;
    inv02 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix643 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644), .A (nx8538)) ;
    dff L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_0 (.Q (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_0), .QB (\$dummy [1194])
        , .D (L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .CLK (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    nor02_2x L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix567 (.Y (
             L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566), .A0 (RST), .A1 (
             L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644)) ;
    dff L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_1 (.Q (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_1), .QB (\$dummy [1195])
        , .D (L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .CLK (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_2 (.Q (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_2), .QB (\$dummy [1196])
        , .D (L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .CLK (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_3 (.Q (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_3), .QB (\$dummy [1197])
        , .D (L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .CLK (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_4 (.Q (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_4), .QB (\$dummy [1198])
        , .D (L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .CLK (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_5 (.Q (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_5), .QB (\$dummy [1199])
        , .D (L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .CLK (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_6 (.Q (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_6), .QB (\$dummy [1200])
        , .D (L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .CLK (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_7 (.Q (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_7), .QB (\$dummy [1201])
        , .D (L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .CLK (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_8 (.Q (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_8), .QB (\$dummy [1202])
        , .D (L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .CLK (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_9 (.Q (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_9), .QB (\$dummy [1203])
        , .D (L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .CLK (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_10 (.Q (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_10), .QB (\$dummy [1204])
        , .D (L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .CLK (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_11 (.Q (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_11), .QB (\$dummy [1205])
        , .D (L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .CLK (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_12 (.Q (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_12), .QB (\$dummy [1206])
        , .D (L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .CLK (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_13 (.Q (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_13), .QB (\$dummy [1207])
        , .D (L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .CLK (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_14 (.Q (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_14), .QB (\$dummy [1208])
        , .D (L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .CLK (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_15 (.Q (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_15), .QB (\$dummy [1209])
        , .D (L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .CLK (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_16 (.Q (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_16), .QB (\$dummy [1210])
        , .D (L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .CLK (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    inv02 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix623 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624), .A (CLK)) ;
    inv02 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix625 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626), .A (CLK)) ;
    inv02 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix627 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628), .A (CLK)) ;
    inv02 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix643 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644), .A (nx8544)) ;
    dff L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_0 (.Q (
        L1_4_L2_3_G5_MINI_ALU_BoothP_0), .QB (\$dummy [1211]), .D (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .CLK (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    nor02_2x L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix567 (.Y (
             L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566), .A0 (RST), .A1 (
             L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    dff L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_1 (.Q (
        L1_4_L2_3_G5_MINI_ALU_BoothP_1), .QB (\$dummy [1212]), .D (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .CLK (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_2 (.Q (
        L1_4_L2_3_G5_MINI_ALU_BoothP_2), .QB (\$dummy [1213]), .D (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .CLK (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_3 (.Q (
        L1_4_L2_3_G5_MINI_ALU_BoothP_3), .QB (\$dummy [1214]), .D (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .CLK (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_4 (.Q (
        L1_4_L2_3_G5_MINI_ALU_BoothP_4), .QB (\$dummy [1215]), .D (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .CLK (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_5 (.Q (
        L1_4_L2_3_G5_MINI_ALU_BoothP_5), .QB (\$dummy [1216]), .D (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .CLK (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_6 (.Q (
        L1_4_L2_3_G5_MINI_ALU_BoothP_6), .QB (\$dummy [1217]), .D (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .CLK (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_7 (.Q (
        L1_4_L2_3_G5_MINI_ALU_BoothP_7), .QB (\$dummy [1218]), .D (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .CLK (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_8 (.Q (
        L1_4_L2_3_G5_MINI_ALU_BoothP_8), .QB (\$dummy [1219]), .D (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .CLK (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_9 (.Q (
        L1_4_L2_3_G5_MINI_ALU_BoothP_9), .QB (\$dummy [1220]), .D (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .CLK (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_10 (.Q (
        L1_4_L2_3_G5_MINI_ALU_BoothP_10), .QB (\$dummy [1221]), .D (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .CLK (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_11 (.Q (
        L1_4_L2_3_G5_MINI_ALU_BoothP_11), .QB (\$dummy [1222]), .D (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .CLK (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_12 (.Q (
        L1_4_L2_3_G5_MINI_ALU_BoothP_12), .QB (\$dummy [1223]), .D (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .CLK (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_13 (.Q (
        L1_4_L2_3_G5_MINI_ALU_BoothP_13), .QB (\$dummy [1224]), .D (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .CLK (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_14 (.Q (
        L1_4_L2_3_G5_MINI_ALU_BoothP_14), .QB (\$dummy [1225]), .D (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .CLK (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_15 (.Q (
        L1_4_L2_3_G5_MINI_ALU_BoothP_15), .QB (\$dummy [1226]), .D (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .CLK (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_16 (.Q (
        L1_4_L2_3_G5_MINI_ALU_BoothP_16), .QB (\$dummy [1227]), .D (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .CLK (
        L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    inv02 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix623 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624), .A (CLK)) ;
    inv02 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix625 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626), .A (CLK)) ;
    inv02 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix627 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628), .A (CLK)) ;
    inv02 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix643 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644), .A (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642)) ;
    xor2 L1_4_L2_4_G5_MINI_ALU_ix83 (.Y (L5Results_1__0), .A0 (
         L5SecondOperands_1__0), .A1 (L5FirstOperands_1__0)) ;
    xnor2 L1_4_L2_4_G5_MINI_ALU_ix380 (.Y (L1_4_L2_4_G5_MINI_ALU_nx379), .A0 (
          L1_4_L2_4_G5_MINI_ALU_nx381), .A1 (L1_4_L2_4_G5_MINI_ALU_nx383)) ;
    nand02 L1_4_L2_4_G5_MINI_ALU_ix382 (.Y (L1_4_L2_4_G5_MINI_ALU_nx381), .A0 (
           L1_4_L2_4_G5_MINI_ALU_BoothOperand_0), .A1 (nx8564)) ;
    xnor2 L1_4_L2_4_G5_MINI_ALU_ix384 (.Y (L1_4_L2_4_G5_MINI_ALU_nx383), .A0 (
          L1_4_L2_4_G5_MINI_ALU_BoothOperand_1), .A1 (
          L1_4_L2_4_G5_MINI_ALU_BoothP_1)) ;
    inv01 L1_4_L2_4_G5_MINI_ALU_ix388 (.Y (L1_4_L2_4_G5_MINI_ALU_nx387), .A (
          L1_4_L2_4_G5_MINI_ALU_BoothP_2)) ;
    xnor2 L1_4_L2_4_G5_MINI_ALU_ix390 (.Y (L1_4_L2_4_G5_MINI_ALU_nx389), .A0 (
          L1_4_L2_4_G5_MINI_ALU_nx391), .A1 (L1_4_L2_4_G5_MINI_ALU_nx395)) ;
    aoi32 L1_4_L2_4_G5_MINI_ALU_ix392 (.Y (L1_4_L2_4_G5_MINI_ALU_nx391), .A0 (
          L1_4_L2_4_G5_MINI_ALU_BoothOperand_0), .A1 (nx8564), .A2 (
          L1_4_L2_4_G5_MINI_ALU_nx154), .B0 (L1_4_L2_4_G5_MINI_ALU_BoothP_1), .B1 (
          L1_4_L2_4_G5_MINI_ALU_BoothOperand_1)) ;
    xnor2 L1_4_L2_4_G5_MINI_ALU_ix396 (.Y (L1_4_L2_4_G5_MINI_ALU_nx395), .A0 (
          L1_4_L2_4_G5_MINI_ALU_BoothOperand_2), .A1 (
          L1_4_L2_4_G5_MINI_ALU_BoothP_2)) ;
    inv01 L1_4_L2_4_G5_MINI_ALU_ix400 (.Y (L1_4_L2_4_G5_MINI_ALU_nx399), .A (
          L1_4_L2_4_G5_MINI_ALU_BoothP_3)) ;
    xnor2 L1_4_L2_4_G5_MINI_ALU_ix402 (.Y (L1_4_L2_4_G5_MINI_ALU_nx401), .A0 (
          L1_4_L2_4_G5_MINI_ALU_nx403), .A1 (L1_4_L2_4_G5_MINI_ALU_nx405)) ;
    xnor2 L1_4_L2_4_G5_MINI_ALU_ix406 (.Y (L1_4_L2_4_G5_MINI_ALU_nx405), .A0 (
          L1_4_L2_4_G5_MINI_ALU_BoothOperand_3), .A1 (
          L1_4_L2_4_G5_MINI_ALU_BoothP_3)) ;
    inv01 L1_4_L2_4_G5_MINI_ALU_ix410 (.Y (L1_4_L2_4_G5_MINI_ALU_nx409), .A (
          L1_4_L2_4_G5_MINI_ALU_BoothP_4)) ;
    xnor2 L1_4_L2_4_G5_MINI_ALU_ix412 (.Y (L1_4_L2_4_G5_MINI_ALU_nx411), .A0 (
          L1_4_L2_4_G5_MINI_ALU_nx413), .A1 (L1_4_L2_4_G5_MINI_ALU_nx415)) ;
    xnor2 L1_4_L2_4_G5_MINI_ALU_ix416 (.Y (L1_4_L2_4_G5_MINI_ALU_nx415), .A0 (
          L1_4_L2_4_G5_MINI_ALU_BoothOperand_4), .A1 (
          L1_4_L2_4_G5_MINI_ALU_BoothP_4)) ;
    inv01 L1_4_L2_4_G5_MINI_ALU_ix420 (.Y (L1_4_L2_4_G5_MINI_ALU_nx419), .A (
          L1_4_L2_4_G5_MINI_ALU_BoothP_5)) ;
    xnor2 L1_4_L2_4_G5_MINI_ALU_ix422 (.Y (L1_4_L2_4_G5_MINI_ALU_nx421), .A0 (
          L1_4_L2_4_G5_MINI_ALU_nx423), .A1 (L1_4_L2_4_G5_MINI_ALU_nx425)) ;
    xnor2 L1_4_L2_4_G5_MINI_ALU_ix426 (.Y (L1_4_L2_4_G5_MINI_ALU_nx425), .A0 (
          L1_4_L2_4_G5_MINI_ALU_BoothOperand_5), .A1 (
          L1_4_L2_4_G5_MINI_ALU_BoothP_5)) ;
    inv01 L1_4_L2_4_G5_MINI_ALU_ix430 (.Y (L1_4_L2_4_G5_MINI_ALU_nx429), .A (
          L1_4_L2_4_G5_MINI_ALU_BoothP_6)) ;
    xnor2 L1_4_L2_4_G5_MINI_ALU_ix432 (.Y (L1_4_L2_4_G5_MINI_ALU_nx431), .A0 (
          L1_4_L2_4_G5_MINI_ALU_nx433), .A1 (L1_4_L2_4_G5_MINI_ALU_nx435)) ;
    xnor2 L1_4_L2_4_G5_MINI_ALU_ix436 (.Y (L1_4_L2_4_G5_MINI_ALU_nx435), .A0 (
          L1_4_L2_4_G5_MINI_ALU_BoothOperand_6), .A1 (
          L1_4_L2_4_G5_MINI_ALU_BoothP_6)) ;
    inv01 L1_4_L2_4_G5_MINI_ALU_ix440 (.Y (L1_4_L2_4_G5_MINI_ALU_nx439), .A (
          L1_4_L2_4_G5_MINI_ALU_BoothP_7)) ;
    xnor2 L1_4_L2_4_G5_MINI_ALU_ix442 (.Y (L1_4_L2_4_G5_MINI_ALU_nx441), .A0 (
          L1_4_L2_4_G5_MINI_ALU_nx443), .A1 (L1_4_L2_4_G5_MINI_ALU_nx445)) ;
    xnor2 L1_4_L2_4_G5_MINI_ALU_ix446 (.Y (L1_4_L2_4_G5_MINI_ALU_nx445), .A0 (
          L1_4_L2_4_G5_MINI_ALU_BoothOperand_7), .A1 (
          L1_4_L2_4_G5_MINI_ALU_BoothP_7)) ;
    inv01 L1_4_L2_4_G5_MINI_ALU_ix450 (.Y (L1_4_L2_4_G5_MINI_ALU_nx449), .A (
          L1_4_L2_4_G5_MINI_ALU_BoothP_8)) ;
    xnor2 L1_4_L2_4_G5_MINI_ALU_ix452 (.Y (L1_4_L2_4_G5_MINI_ALU_nx451), .A0 (
          L1_4_L2_4_G5_MINI_ALU_nx453), .A1 (L1_4_L2_4_G5_MINI_ALU_nx455)) ;
    xnor2 L1_4_L2_4_G5_MINI_ALU_ix456 (.Y (L1_4_L2_4_G5_MINI_ALU_nx455), .A0 (
          L1_4_L2_4_G5_MINI_ALU_BoothOperand_8), .A1 (
          L1_4_L2_4_G5_MINI_ALU_BoothP_8)) ;
    xor2 L1_4_L2_4_G5_MINI_ALU_ix317 (.Y (L1_4_L2_4_G5_MINI_ALU_nx316), .A0 (
         L1_4_L2_4_G5_MINI_ALU_nx461), .A1 (L1_4_L2_4_G5_MINI_ALU_nx463)) ;
    xnor2 L1_4_L2_4_G5_MINI_ALU_ix464 (.Y (L1_4_L2_4_G5_MINI_ALU_nx463), .A0 (
          L1_4_L2_4_G5_MINI_ALU_BoothOperand_9), .A1 (
          L1_4_L2_4_G5_MINI_ALU_BoothP_9)) ;
    xor2 L1_4_L2_4_G5_MINI_ALU_ix337 (.Y (L1_4_L2_4_G5_MINI_ALU_nx336), .A0 (
         L1_4_L2_4_G5_MINI_ALU_nx467), .A1 (L1_4_L2_4_G5_MINI_ALU_nx471)) ;
    inv01 L1_4_L2_4_G5_MINI_ALU_ix470 (.Y (L1_4_L2_4_G5_MINI_ALU_nx469), .A (
          L1_4_L2_4_G5_MINI_ALU_BoothP_9)) ;
    xnor2 L1_4_L2_4_G5_MINI_ALU_ix472 (.Y (L1_4_L2_4_G5_MINI_ALU_nx471), .A0 (
          L1_4_L2_4_G5_MINI_ALU_BoothOperand_10), .A1 (
          L1_4_L2_4_G5_MINI_ALU_BoothP_10)) ;
    xor2 L1_4_L2_4_G5_MINI_ALU_ix357 (.Y (L1_4_L2_4_G5_MINI_ALU_nx356), .A0 (
         L1_4_L2_4_G5_MINI_ALU_nx475), .A1 (L1_4_L2_4_G5_MINI_ALU_nx479)) ;
    inv01 L1_4_L2_4_G5_MINI_ALU_ix478 (.Y (L1_4_L2_4_G5_MINI_ALU_nx477), .A (
          L1_4_L2_4_G5_MINI_ALU_BoothP_10)) ;
    xnor2 L1_4_L2_4_G5_MINI_ALU_ix480 (.Y (L1_4_L2_4_G5_MINI_ALU_nx479), .A0 (
          L1_4_L2_4_G5_MINI_ALU_BoothOperand_11), .A1 (
          L1_4_L2_4_G5_MINI_ALU_BoothP_11)) ;
    xor2 L1_4_L2_4_G5_MINI_ALU_ix377 (.Y (L1_4_L2_4_G5_MINI_ALU_nx376), .A0 (
         L1_4_L2_4_G5_MINI_ALU_nx483), .A1 (L1_4_L2_4_G5_MINI_ALU_nx487)) ;
    inv01 L1_4_L2_4_G5_MINI_ALU_ix486 (.Y (L1_4_L2_4_G5_MINI_ALU_nx485), .A (
          L1_4_L2_4_G5_MINI_ALU_BoothP_11)) ;
    xnor2 L1_4_L2_4_G5_MINI_ALU_ix488 (.Y (L1_4_L2_4_G5_MINI_ALU_nx487), .A0 (
          L1_4_L2_4_G5_MINI_ALU_BoothOperand_12), .A1 (
          L1_4_L2_4_G5_MINI_ALU_BoothP_12)) ;
    xor2 L1_4_L2_4_G5_MINI_ALU_ix397 (.Y (L1_4_L2_4_G5_MINI_ALU_nx396), .A0 (
         L1_4_L2_4_G5_MINI_ALU_nx491), .A1 (L1_4_L2_4_G5_MINI_ALU_nx495)) ;
    inv01 L1_4_L2_4_G5_MINI_ALU_ix494 (.Y (L1_4_L2_4_G5_MINI_ALU_nx493), .A (
          L1_4_L2_4_G5_MINI_ALU_BoothP_12)) ;
    xnor2 L1_4_L2_4_G5_MINI_ALU_ix496 (.Y (L1_4_L2_4_G5_MINI_ALU_nx495), .A0 (
          L1_4_L2_4_G5_MINI_ALU_BoothOperand_13), .A1 (
          L1_4_L2_4_G5_MINI_ALU_BoothP_13)) ;
    xor2 L1_4_L2_4_G5_MINI_ALU_ix417 (.Y (L1_4_L2_4_G5_MINI_ALU_nx416), .A0 (
         L1_4_L2_4_G5_MINI_ALU_nx499), .A1 (L1_4_L2_4_G5_MINI_ALU_nx503)) ;
    inv01 L1_4_L2_4_G5_MINI_ALU_ix502 (.Y (L1_4_L2_4_G5_MINI_ALU_nx501), .A (
          L1_4_L2_4_G5_MINI_ALU_BoothP_13)) ;
    xnor2 L1_4_L2_4_G5_MINI_ALU_ix504 (.Y (L1_4_L2_4_G5_MINI_ALU_nx503), .A0 (
          L1_4_L2_4_G5_MINI_ALU_BoothOperand_14), .A1 (
          L1_4_L2_4_G5_MINI_ALU_BoothP_14)) ;
    xor2 L1_4_L2_4_G5_MINI_ALU_ix437 (.Y (L1_4_L2_4_G5_MINI_ALU_nx436), .A0 (
         L1_4_L2_4_G5_MINI_ALU_nx507), .A1 (L1_4_L2_4_G5_MINI_ALU_nx511)) ;
    inv01 L1_4_L2_4_G5_MINI_ALU_ix510 (.Y (L1_4_L2_4_G5_MINI_ALU_nx509), .A (
          L1_4_L2_4_G5_MINI_ALU_BoothP_14)) ;
    xnor2 L1_4_L2_4_G5_MINI_ALU_ix512 (.Y (L1_4_L2_4_G5_MINI_ALU_nx511), .A0 (
          L1_4_L2_4_G5_MINI_ALU_BoothOperand_15), .A1 (
          L1_4_L2_4_G5_MINI_ALU_BoothP_15)) ;
    xnor2 L1_4_L2_4_G5_MINI_ALU_ix457 (.Y (L1_4_L2_4_G5_MINI_ALU_nx456), .A0 (
          L1_4_L2_4_G5_MINI_ALU_nx515), .A1 (L1_4_L2_4_G5_MINI_ALU_nx454)) ;
    inv01 L1_4_L2_4_G5_MINI_ALU_ix518 (.Y (L1_4_L2_4_G5_MINI_ALU_nx517), .A (
          L1_4_L2_4_G5_MINI_ALU_BoothP_15)) ;
    xor2 L1_4_L2_4_G5_MINI_ALU_ix455 (.Y (L1_4_L2_4_G5_MINI_ALU_nx454), .A0 (
         L1_4_L2_4_G5_MINI_ALU_BoothOperand_16), .A1 (
         L1_4_L2_4_G5_MINI_ALU_BoothP_16)) ;
    mux21_ni L1_4_L2_4_G5_MINI_ALU_ix91 (.Y (L5SecondOperands_1__0), .A0 (
             L1_4_L2_4_G5_MINI_ALU_BoothP_1), .A1 (WindowDin_4__4__0), .S0 (
             Instr)) ;
    mux21_ni L1_4_L2_4_G5_MINI_ALU_ix99 (.Y (L5SecondOperands_1__1), .A0 (
             L1_4_L2_4_G5_MINI_ALU_BoothP_2), .A1 (WindowDin_4__4__1), .S0 (
             Instr)) ;
    mux21_ni L1_4_L2_4_G5_MINI_ALU_ix107 (.Y (L5SecondOperands_1__2), .A0 (
             L1_4_L2_4_G5_MINI_ALU_BoothP_3), .A1 (WindowDin_4__4__2), .S0 (
             Instr)) ;
    mux21_ni L1_4_L2_4_G5_MINI_ALU_ix115 (.Y (L5SecondOperands_1__3), .A0 (
             L1_4_L2_4_G5_MINI_ALU_BoothP_4), .A1 (WindowDin_4__4__3), .S0 (
             Instr)) ;
    mux21_ni L1_4_L2_4_G5_MINI_ALU_ix123 (.Y (L5SecondOperands_1__4), .A0 (
             L1_4_L2_4_G5_MINI_ALU_BoothP_5), .A1 (WindowDin_4__4__4), .S0 (
             Instr)) ;
    mux21_ni L1_4_L2_4_G5_MINI_ALU_ix131 (.Y (L5SecondOperands_1__5), .A0 (
             L1_4_L2_4_G5_MINI_ALU_BoothP_6), .A1 (WindowDin_4__4__5), .S0 (
             Instr)) ;
    mux21_ni L1_4_L2_4_G5_MINI_ALU_ix139 (.Y (L5SecondOperands_1__6), .A0 (
             L1_4_L2_4_G5_MINI_ALU_BoothP_7), .A1 (WindowDin_4__4__6), .S0 (
             Instr)) ;
    mux21_ni L1_4_L2_4_G5_MINI_ALU_ix147 (.Y (L5SecondOperands_1__7), .A0 (
             L1_4_L2_4_G5_MINI_ALU_BoothP_8), .A1 (WindowDin_4__4__7), .S0 (
             Instr)) ;
    xor2 L1_4_L2_4_G5_MINI_ALU_ix77 (.Y (L5Results_1__1), .A0 (
         L1_4_L2_4_G5_MINI_ALU_nx529), .A1 (L1_4_L2_4_G5_MINI_ALU_nx531)) ;
    nand02 L1_4_L2_4_G5_MINI_ALU_ix530 (.Y (L1_4_L2_4_G5_MINI_ALU_nx529), .A0 (
           L5SecondOperands_1__0), .A1 (L5FirstOperands_1__0)) ;
    xnor2 L1_4_L2_4_G5_MINI_ALU_ix532 (.Y (L1_4_L2_4_G5_MINI_ALU_nx531), .A0 (
          L5SecondOperands_1__1), .A1 (L5FirstOperands_1__1)) ;
    xor2 L1_4_L2_4_G5_MINI_ALU_ix75 (.Y (L5Results_1__2), .A0 (
         L1_4_L2_4_G5_MINI_ALU_nx534), .A1 (L1_4_L2_4_G5_MINI_ALU_nx537)) ;
    aoi32 L1_4_L2_4_G5_MINI_ALU_ix535 (.Y (L1_4_L2_4_G5_MINI_ALU_nx534), .A0 (
          L5SecondOperands_1__0), .A1 (L5FirstOperands_1__0), .A2 (
          L1_4_L2_4_G5_MINI_ALU_nx30), .B0 (L5FirstOperands_1__1), .B1 (
          L5SecondOperands_1__1)) ;
    xnor2 L1_4_L2_4_G5_MINI_ALU_ix538 (.Y (L1_4_L2_4_G5_MINI_ALU_nx537), .A0 (
          L5SecondOperands_1__2), .A1 (L5FirstOperands_1__2)) ;
    xor2 L1_4_L2_4_G5_MINI_ALU_ix73 (.Y (L5Results_1__3), .A0 (
         L1_4_L2_4_G5_MINI_ALU_nx540), .A1 (L1_4_L2_4_G5_MINI_ALU_nx544)) ;
    aoi22 L1_4_L2_4_G5_MINI_ALU_ix541 (.Y (L1_4_L2_4_G5_MINI_ALU_nx540), .A0 (
          L5FirstOperands_1__2), .A1 (L5SecondOperands_1__2), .B0 (
          L1_4_L2_4_G5_MINI_ALU_nx40), .B1 (L1_4_L2_4_G5_MINI_ALU_nx24)) ;
    xnor2 L1_4_L2_4_G5_MINI_ALU_ix545 (.Y (L1_4_L2_4_G5_MINI_ALU_nx544), .A0 (
          L5SecondOperands_1__3), .A1 (L5FirstOperands_1__3)) ;
    xor2 L1_4_L2_4_G5_MINI_ALU_ix71 (.Y (L5Results_1__4), .A0 (
         L1_4_L2_4_G5_MINI_ALU_nx547), .A1 (L1_4_L2_4_G5_MINI_ALU_nx551)) ;
    aoi22 L1_4_L2_4_G5_MINI_ALU_ix548 (.Y (L1_4_L2_4_G5_MINI_ALU_nx547), .A0 (
          L5FirstOperands_1__3), .A1 (L5SecondOperands_1__3), .B0 (
          L1_4_L2_4_G5_MINI_ALU_nx44), .B1 (L1_4_L2_4_G5_MINI_ALU_nx18)) ;
    xnor2 L1_4_L2_4_G5_MINI_ALU_ix552 (.Y (L1_4_L2_4_G5_MINI_ALU_nx551), .A0 (
          L5SecondOperands_1__4), .A1 (L5FirstOperands_1__4)) ;
    xor2 L1_4_L2_4_G5_MINI_ALU_ix69 (.Y (L5Results_1__5), .A0 (
         L1_4_L2_4_G5_MINI_ALU_nx554), .A1 (L1_4_L2_4_G5_MINI_ALU_nx558)) ;
    aoi22 L1_4_L2_4_G5_MINI_ALU_ix555 (.Y (L1_4_L2_4_G5_MINI_ALU_nx554), .A0 (
          L5FirstOperands_1__4), .A1 (L5SecondOperands_1__4), .B0 (
          L1_4_L2_4_G5_MINI_ALU_nx48), .B1 (L1_4_L2_4_G5_MINI_ALU_nx12)) ;
    xnor2 L1_4_L2_4_G5_MINI_ALU_ix559 (.Y (L1_4_L2_4_G5_MINI_ALU_nx558), .A0 (
          L5SecondOperands_1__5), .A1 (L5FirstOperands_1__5)) ;
    xor2 L1_4_L2_4_G5_MINI_ALU_ix67 (.Y (L5Results_1__6), .A0 (
         L1_4_L2_4_G5_MINI_ALU_nx561), .A1 (L1_4_L2_4_G5_MINI_ALU_nx565)) ;
    aoi22 L1_4_L2_4_G5_MINI_ALU_ix562 (.Y (L1_4_L2_4_G5_MINI_ALU_nx561), .A0 (
          L5FirstOperands_1__5), .A1 (L5SecondOperands_1__5), .B0 (
          L1_4_L2_4_G5_MINI_ALU_nx52), .B1 (L1_4_L2_4_G5_MINI_ALU_nx6)) ;
    xnor2 L1_4_L2_4_G5_MINI_ALU_ix566 (.Y (L1_4_L2_4_G5_MINI_ALU_nx565), .A0 (
          L5SecondOperands_1__6), .A1 (L5FirstOperands_1__6)) ;
    xnor2 L1_4_L2_4_G5_MINI_ALU_ix65 (.Y (L5Results_1__7), .A0 (
          L1_4_L2_4_G5_MINI_ALU_nx568), .A1 (L1_4_L2_4_G5_MINI_ALU_nx62)) ;
    aoi22 L1_4_L2_4_G5_MINI_ALU_ix569 (.Y (L1_4_L2_4_G5_MINI_ALU_nx568), .A0 (
          L5FirstOperands_1__6), .A1 (L5SecondOperands_1__6), .B0 (
          L1_4_L2_4_G5_MINI_ALU_nx56), .B1 (L1_4_L2_4_G5_MINI_ALU_nx0)) ;
    xor2 L1_4_L2_4_G5_MINI_ALU_ix63 (.Y (L1_4_L2_4_G5_MINI_ALU_nx62), .A0 (
         L5SecondOperands_1__7), .A1 (L5FirstOperands_1__7)) ;
    inv01 L1_4_L2_4_G5_MINI_ALU_ix155 (.Y (L1_4_L2_4_G5_MINI_ALU_nx154), .A (
          L1_4_L2_4_G5_MINI_ALU_nx383)) ;
    inv01 L1_4_L2_4_G5_MINI_ALU_ix57 (.Y (L1_4_L2_4_G5_MINI_ALU_nx56), .A (
          L1_4_L2_4_G5_MINI_ALU_nx561)) ;
    inv01 L1_4_L2_4_G5_MINI_ALU_ix53 (.Y (L1_4_L2_4_G5_MINI_ALU_nx52), .A (
          L1_4_L2_4_G5_MINI_ALU_nx554)) ;
    inv01 L1_4_L2_4_G5_MINI_ALU_ix49 (.Y (L1_4_L2_4_G5_MINI_ALU_nx48), .A (
          L1_4_L2_4_G5_MINI_ALU_nx547)) ;
    inv01 L1_4_L2_4_G5_MINI_ALU_ix45 (.Y (L1_4_L2_4_G5_MINI_ALU_nx44), .A (
          L1_4_L2_4_G5_MINI_ALU_nx540)) ;
    inv01 L1_4_L2_4_G5_MINI_ALU_ix41 (.Y (L1_4_L2_4_G5_MINI_ALU_nx40), .A (
          L1_4_L2_4_G5_MINI_ALU_nx534)) ;
    inv01 L1_4_L2_4_G5_MINI_ALU_ix31 (.Y (L1_4_L2_4_G5_MINI_ALU_nx30), .A (
          L1_4_L2_4_G5_MINI_ALU_nx531)) ;
    inv01 L1_4_L2_4_G5_MINI_ALU_ix25 (.Y (L1_4_L2_4_G5_MINI_ALU_nx24), .A (
          L1_4_L2_4_G5_MINI_ALU_nx537)) ;
    inv01 L1_4_L2_4_G5_MINI_ALU_ix19 (.Y (L1_4_L2_4_G5_MINI_ALU_nx18), .A (
          L1_4_L2_4_G5_MINI_ALU_nx544)) ;
    inv01 L1_4_L2_4_G5_MINI_ALU_ix13 (.Y (L1_4_L2_4_G5_MINI_ALU_nx12), .A (
          L1_4_L2_4_G5_MINI_ALU_nx551)) ;
    inv01 L1_4_L2_4_G5_MINI_ALU_ix7 (.Y (L1_4_L2_4_G5_MINI_ALU_nx6), .A (
          L1_4_L2_4_G5_MINI_ALU_nx558)) ;
    inv01 L1_4_L2_4_G5_MINI_ALU_ix1 (.Y (L1_4_L2_4_G5_MINI_ALU_nx0), .A (
          L1_4_L2_4_G5_MINI_ALU_nx565)) ;
    fake_gnd L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix216 (.Y (
             L1_4_L2_4_G5_MINI_ALU_WindowCellShiftedLeft_16)) ;
    nor02ii L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix81 (.Y (
            L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_nx80), .A0 (Instr), .A1 (Start)) ;
    aoi21 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix77 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_10), .A0 (
          FilterDin_4__4__1), .A1 (FilterDin_4__4__0), .B0 (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_nx4)) ;
    nor02_2x L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix5 (.Y (
             L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_nx4), .A0 (FilterDin_4__4__0), .A1 (
             FilterDin_4__4__1)) ;
    aoi21 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix67 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_11), .A0 (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_nx328), .A1 (FilterDin_4__4__2), .B0 (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_nx8)) ;
    nor03_2x L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix9 (.Y (
             L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_nx8), .A0 (FilterDin_4__4__2), .A1 (
             FilterDin_4__4__0), .A2 (FilterDin_4__4__1)) ;
    xnor2 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix59 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_12), .A0 (
          FilterDin_4__4__3), .A1 (L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_nx8)) ;
    xnor2 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix51 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_13), .A0 (
          FilterDin_4__4__4), .A1 (L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_nx12)) ;
    nor04 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix13 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_nx12), .A0 (FilterDin_4__4__3), .A1 (
          FilterDin_4__4__2), .A2 (FilterDin_4__4__0), .A3 (FilterDin_4__4__1)
          ) ;
    xnor2 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix43 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_14), .A0 (
          FilterDin_4__4__5), .A1 (L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_nx16)) ;
    nor02ii L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix17 (.Y (
            L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_nx16), .A0 (FilterDin_4__4__4), .A1 (
            L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_nx12)) ;
    xnor2 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix35 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_15), .A0 (
          FilterDin_4__4__6), .A1 (L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_nx20)) ;
    nor02ii L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix21 (.Y (
            L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_nx20), .A0 (FilterDin_4__4__5), .A1 (
            L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_nx16)) ;
    xnor2 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix27 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_16), .A0 (
          FilterDin_4__4__7), .A1 (L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_nx24)) ;
    nor02ii L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix25 (.Y (
            L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_nx24), .A0 (FilterDin_4__4__6), .A1 (
            L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_nx20)) ;
    inv01 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix329 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_nx328), .A (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_nx4)) ;
    inv02 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix383 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_nx384), .A (
          L1_4_L2_4_G5_MINI_ALU_BoothP_0)) ;
    dff L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_0 (.Q (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_0), .QB (\$dummy [1228])
        , .D (L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .CLK (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    nor02_2x L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix567 (.Y (
             L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566), .A0 (RST), .A1 (
             L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644)) ;
    dff L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_1 (.Q (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_1), .QB (\$dummy [1229])
        , .D (L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .CLK (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_2 (.Q (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_2), .QB (\$dummy [1230])
        , .D (L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .CLK (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_3 (.Q (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_3), .QB (\$dummy [1231])
        , .D (L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .CLK (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_4 (.Q (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_4), .QB (\$dummy [1232])
        , .D (L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .CLK (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_5 (.Q (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_5), .QB (\$dummy [1233])
        , .D (L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .CLK (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_6 (.Q (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_6), .QB (\$dummy [1234])
        , .D (L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .CLK (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624)) ;
    dff L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_7 (.Q (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_7), .QB (\$dummy [1235])
        , .D (L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .CLK (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_8 (.Q (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_8), .QB (\$dummy [1236])
        , .D (L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .CLK (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_9 (.Q (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_9), .QB (\$dummy [1237])
        , .D (L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .CLK (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_10 (.Q (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_10), .QB (\$dummy [1238])
        , .D (L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .CLK (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_11 (.Q (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_11), .QB (\$dummy [1239])
        , .D (L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .CLK (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_12 (.Q (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_12), .QB (\$dummy [1240])
        , .D (L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .CLK (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_13 (.Q (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_13), .QB (\$dummy [1241])
        , .D (L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .CLK (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626)) ;
    dff L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_14 (.Q (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_14), .QB (\$dummy [1242])
        , .D (L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .CLK (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_15 (.Q (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_15), .QB (\$dummy [1243])
        , .D (L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .CLK (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    dff L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_reg_Dout_16 (.Q (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_16), .QB (\$dummy [1244])
        , .D (L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .CLK (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628)) ;
    inv02 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix623 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx624), .A (CLK)) ;
    inv02 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix625 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx626), .A (CLK)) ;
    inv02 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix627 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx628), .A (CLK)) ;
    inv02 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix643 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx644), .A (nx8578)) ;
    dff L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_0 (.Q (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_0), .QB (\$dummy [1245])
        , .D (L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .CLK (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    nor02_2x L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix567 (.Y (
             L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566), .A0 (RST), .A1 (
             L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644)) ;
    dff L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_1 (.Q (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_1), .QB (\$dummy [1246])
        , .D (L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .CLK (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_2 (.Q (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_2), .QB (\$dummy [1247])
        , .D (L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .CLK (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_3 (.Q (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_3), .QB (\$dummy [1248])
        , .D (L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .CLK (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_4 (.Q (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_4), .QB (\$dummy [1249])
        , .D (L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .CLK (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_5 (.Q (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_5), .QB (\$dummy [1250])
        , .D (L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .CLK (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_6 (.Q (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_6), .QB (\$dummy [1251])
        , .D (L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .CLK (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624)) ;
    dff L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_7 (.Q (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_7), .QB (\$dummy [1252])
        , .D (L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .CLK (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_8 (.Q (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_8), .QB (\$dummy [1253])
        , .D (L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .CLK (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_9 (.Q (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_9), .QB (\$dummy [1254])
        , .D (L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .CLK (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_10 (.Q (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_10), .QB (\$dummy [1255])
        , .D (L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .CLK (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_11 (.Q (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_11), .QB (\$dummy [1256])
        , .D (L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .CLK (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_12 (.Q (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_12), .QB (\$dummy [1257])
        , .D (L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .CLK (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_13 (.Q (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_13), .QB (\$dummy [1258])
        , .D (L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .CLK (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626)) ;
    dff L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_14 (.Q (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_14), .QB (\$dummy [1259])
        , .D (L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .CLK (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_15 (.Q (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_15), .QB (\$dummy [1260])
        , .D (L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .CLK (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    dff L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_reg_Dout_16 (.Q (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_16), .QB (\$dummy [1261])
        , .D (L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .CLK (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628)) ;
    inv02 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix623 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx624), .A (CLK)) ;
    inv02 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix625 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx626), .A (CLK)) ;
    inv02 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix627 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx628), .A (CLK)) ;
    inv02 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix643 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx644), .A (nx8584)) ;
    dff L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_0 (.Q (
        L1_4_L2_4_G5_MINI_ALU_BoothP_0), .QB (\$dummy [1262]), .D (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .CLK (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    nor02_2x L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix567 (.Y (
             L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566), .A0 (RST), .A1 (
             L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    dff L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_1 (.Q (
        L1_4_L2_4_G5_MINI_ALU_BoothP_1), .QB (\$dummy [1263]), .D (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .CLK (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_2 (.Q (
        L1_4_L2_4_G5_MINI_ALU_BoothP_2), .QB (\$dummy [1264]), .D (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .CLK (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_3 (.Q (
        L1_4_L2_4_G5_MINI_ALU_BoothP_3), .QB (\$dummy [1265]), .D (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .CLK (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_4 (.Q (
        L1_4_L2_4_G5_MINI_ALU_BoothP_4), .QB (\$dummy [1266]), .D (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .CLK (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_5 (.Q (
        L1_4_L2_4_G5_MINI_ALU_BoothP_5), .QB (\$dummy [1267]), .D (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .CLK (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_6 (.Q (
        L1_4_L2_4_G5_MINI_ALU_BoothP_6), .QB (\$dummy [1268]), .D (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .CLK (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624)) ;
    dff L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_7 (.Q (
        L1_4_L2_4_G5_MINI_ALU_BoothP_7), .QB (\$dummy [1269]), .D (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .CLK (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_8 (.Q (
        L1_4_L2_4_G5_MINI_ALU_BoothP_8), .QB (\$dummy [1270]), .D (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .CLK (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_9 (.Q (
        L1_4_L2_4_G5_MINI_ALU_BoothP_9), .QB (\$dummy [1271]), .D (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .CLK (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_10 (.Q (
        L1_4_L2_4_G5_MINI_ALU_BoothP_10), .QB (\$dummy [1272]), .D (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .CLK (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_11 (.Q (
        L1_4_L2_4_G5_MINI_ALU_BoothP_11), .QB (\$dummy [1273]), .D (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .CLK (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_12 (.Q (
        L1_4_L2_4_G5_MINI_ALU_BoothP_12), .QB (\$dummy [1274]), .D (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .CLK (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_13 (.Q (
        L1_4_L2_4_G5_MINI_ALU_BoothP_13), .QB (\$dummy [1275]), .D (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .CLK (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626)) ;
    dff L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_14 (.Q (
        L1_4_L2_4_G5_MINI_ALU_BoothP_14), .QB (\$dummy [1276]), .D (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .CLK (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_15 (.Q (
        L1_4_L2_4_G5_MINI_ALU_BoothP_15), .QB (\$dummy [1277]), .D (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .CLK (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    dff L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_reg_Dout_16 (.Q (
        L1_4_L2_4_G5_MINI_ALU_BoothP_16), .QB (\$dummy [1278]), .D (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .CLK (
        L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628)) ;
    inv02 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix623 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx624), .A (CLK)) ;
    inv02 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix625 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx626), .A (CLK)) ;
    inv02 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix627 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx628), .A (CLK)) ;
    inv02 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix643 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644), .A (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642)) ;
    oai22 ix61 (.Y (Result[3]), .A0 (nx1336), .A1 (nx1338), .B0 (nx1340), .B1 (
          Instr)) ;
    inv01 ix1335 (.Y (nx1336), .A (L5Results_1__6)) ;
    inv01 ix1337 (.Y (nx1338), .A (nx22)) ;
    inv01 ix1339 (.Y (nx1340), .A (L5Results_1__3)) ;
    oai22 ix69 (.Y (Result[4]), .A0 (nx1342), .A1 (nx1338), .B0 (nx1344), .B1 (
          Instr)) ;
    inv01 ix1341 (.Y (nx1342), .A (L5Results_1__7)) ;
    inv01 ix1343 (.Y (nx1344), .A (L5Results_1__4)) ;
    mux21 ACCELERATOR_COUNTER_ix92 (.Y (ACCELERATOR_COUNTER_nx91), .A0 (nx1346)
          , .A1 (nx993), .S0 (Done)) ;
    inv01 ix1345 (.Y (nx1346), .A (ACCELERATOR_COUNTER_nx6)) ;
    mux21 ACCELERATOR_COUNTER_ix102 (.Y (ACCELERATOR_COUNTER_nx101), .A0 (nx1348
          ), .A1 (nx995), .S0 (Done)) ;
    inv01 ix1347 (.Y (nx1348), .A (ACCELERATOR_COUNTER_nx12)) ;
    mux21 ACCELERATOR_COUNTER_ix112 (.Y (ACCELERATOR_COUNTER_nx111), .A0 (nx1350
          ), .A1 (nx1352), .S0 (Done)) ;
    inv01 ix1349 (.Y (nx1350), .A (ACCELERATOR_COUNTER_nx18)) ;
    inv01 ix1351 (.Y (nx1352), .A (CounterOut_3)) ;
    xnor2 ACCELERATOR_COUNTER_ix82 (.Y (ACCELERATOR_COUNTER_nx81), .A0 (
          CounterOut_0), .A1 (Done)) ;
    mux21 L1_0_L2_0_G1_MINI_ALU_ix404 (.Y (L1_0_L2_0_G1_MINI_ALU_nx403), .A0 (
          nx1354), .A1 (L1_0_L2_0_G1_MINI_ALU_BoothP_2), .S0 (
          L1_0_L2_0_G1_MINI_ALU_nx395)) ;
    inv01 ix1353 (.Y (nx1354), .A (L1_0_L2_0_G1_MINI_ALU_nx391)) ;
    mux21 L1_0_L2_0_G1_MINI_ALU_ix414 (.Y (L1_0_L2_0_G1_MINI_ALU_nx413), .A0 (
          nx1356), .A1 (L1_0_L2_0_G1_MINI_ALU_BoothP_3), .S0 (
          L1_0_L2_0_G1_MINI_ALU_nx405)) ;
    inv01 ix1355 (.Y (nx1356), .A (L1_0_L2_0_G1_MINI_ALU_nx403)) ;
    mux21 L1_0_L2_0_G1_MINI_ALU_ix424 (.Y (L1_0_L2_0_G1_MINI_ALU_nx423), .A0 (
          nx1358), .A1 (L1_0_L2_0_G1_MINI_ALU_BoothP_4), .S0 (
          L1_0_L2_0_G1_MINI_ALU_nx415)) ;
    inv01 ix1357 (.Y (nx1358), .A (L1_0_L2_0_G1_MINI_ALU_nx413)) ;
    mux21 L1_0_L2_0_G1_MINI_ALU_ix434 (.Y (L1_0_L2_0_G1_MINI_ALU_nx433), .A0 (
          nx1360), .A1 (L1_0_L2_0_G1_MINI_ALU_BoothP_5), .S0 (
          L1_0_L2_0_G1_MINI_ALU_nx425)) ;
    inv01 ix1359 (.Y (nx1360), .A (L1_0_L2_0_G1_MINI_ALU_nx423)) ;
    mux21 L1_0_L2_0_G1_MINI_ALU_ix444 (.Y (L1_0_L2_0_G1_MINI_ALU_nx443), .A0 (
          nx1362), .A1 (L1_0_L2_0_G1_MINI_ALU_BoothP_6), .S0 (
          L1_0_L2_0_G1_MINI_ALU_nx435)) ;
    inv01 ix1361 (.Y (nx1362), .A (L1_0_L2_0_G1_MINI_ALU_nx433)) ;
    mux21 L1_0_L2_0_G1_MINI_ALU_ix454 (.Y (L1_0_L2_0_G1_MINI_ALU_nx453), .A0 (
          nx1364), .A1 (L1_0_L2_0_G1_MINI_ALU_BoothP_7), .S0 (
          L1_0_L2_0_G1_MINI_ALU_nx445)) ;
    inv01 ix1363 (.Y (nx1364), .A (L1_0_L2_0_G1_MINI_ALU_nx443)) ;
    mux21 L1_0_L2_0_G1_MINI_ALU_ix462 (.Y (L1_0_L2_0_G1_MINI_ALU_nx461), .A0 (
          nx1366), .A1 (L1_0_L2_0_G1_MINI_ALU_BoothP_8), .S0 (
          L1_0_L2_0_G1_MINI_ALU_nx455)) ;
    inv01 ix1365 (.Y (nx1366), .A (L1_0_L2_0_G1_MINI_ALU_nx453)) ;
    mux21 L1_0_L2_0_G1_MINI_ALU_ix468 (.Y (L1_0_L2_0_G1_MINI_ALU_nx467), .A0 (
          nx1368), .A1 (L1_0_L2_0_G1_MINI_ALU_BoothP_9), .S0 (
          L1_0_L2_0_G1_MINI_ALU_nx463)) ;
    inv01 ix1367 (.Y (nx1368), .A (L1_0_L2_0_G1_MINI_ALU_nx461)) ;
    mux21 L1_0_L2_0_G1_MINI_ALU_ix476 (.Y (L1_0_L2_0_G1_MINI_ALU_nx475), .A0 (
          nx1370), .A1 (L1_0_L2_0_G1_MINI_ALU_BoothP_10), .S0 (
          L1_0_L2_0_G1_MINI_ALU_nx471)) ;
    inv01 ix1369 (.Y (nx1370), .A (L1_0_L2_0_G1_MINI_ALU_nx467)) ;
    mux21 L1_0_L2_0_G1_MINI_ALU_ix484 (.Y (L1_0_L2_0_G1_MINI_ALU_nx483), .A0 (
          nx1372), .A1 (L1_0_L2_0_G1_MINI_ALU_BoothP_11), .S0 (
          L1_0_L2_0_G1_MINI_ALU_nx479)) ;
    inv01 ix1371 (.Y (nx1372), .A (L1_0_L2_0_G1_MINI_ALU_nx475)) ;
    mux21 L1_0_L2_0_G1_MINI_ALU_ix492 (.Y (L1_0_L2_0_G1_MINI_ALU_nx491), .A0 (
          nx1374), .A1 (L1_0_L2_0_G1_MINI_ALU_BoothP_12), .S0 (
          L1_0_L2_0_G1_MINI_ALU_nx487)) ;
    inv01 ix1373 (.Y (nx1374), .A (L1_0_L2_0_G1_MINI_ALU_nx483)) ;
    mux21 L1_0_L2_0_G1_MINI_ALU_ix500 (.Y (L1_0_L2_0_G1_MINI_ALU_nx499), .A0 (
          nx1376), .A1 (L1_0_L2_0_G1_MINI_ALU_BoothP_13), .S0 (
          L1_0_L2_0_G1_MINI_ALU_nx495)) ;
    inv01 ix1375 (.Y (nx1376), .A (L1_0_L2_0_G1_MINI_ALU_nx491)) ;
    mux21 L1_0_L2_0_G1_MINI_ALU_ix508 (.Y (L1_0_L2_0_G1_MINI_ALU_nx507), .A0 (
          nx1378), .A1 (L1_0_L2_0_G1_MINI_ALU_BoothP_14), .S0 (
          L1_0_L2_0_G1_MINI_ALU_nx503)) ;
    inv01 ix1377 (.Y (nx1378), .A (L1_0_L2_0_G1_MINI_ALU_nx499)) ;
    mux21 L1_0_L2_0_G1_MINI_ALU_ix516 (.Y (L1_0_L2_0_G1_MINI_ALU_nx515), .A0 (
          nx1380), .A1 (L1_0_L2_0_G1_MINI_ALU_BoothP_15), .S0 (
          L1_0_L2_0_G1_MINI_ALU_nx511)) ;
    inv01 ix1379 (.Y (nx1380), .A (L1_0_L2_0_G1_MINI_ALU_nx507)) ;
    mux21 L1_0_L2_0_G1_MINI_ALU_ix161 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_1), .A0 (nx1382), .A1 (
          L1_0_L2_0_G1_MINI_ALU_nx379), .S0 (nx7556)) ;
    inv01 ix1381 (.Y (nx1382), .A (L1_0_L2_0_G1_MINI_ALU_BoothP_1)) ;
    mux21 L1_0_L2_0_G1_MINI_ALU_ix181 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_2), .A0 (
          L1_0_L2_0_G1_MINI_ALU_nx387), .A1 (L1_0_L2_0_G1_MINI_ALU_nx389), .S0 (
          nx7556)) ;
    mux21 L1_0_L2_0_G1_MINI_ALU_ix201 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_3), .A0 (
          L1_0_L2_0_G1_MINI_ALU_nx399), .A1 (L1_0_L2_0_G1_MINI_ALU_nx401), .S0 (
          nx7556)) ;
    mux21 L1_0_L2_0_G1_MINI_ALU_ix221 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_4), .A0 (
          L1_0_L2_0_G1_MINI_ALU_nx409), .A1 (L1_0_L2_0_G1_MINI_ALU_nx411), .S0 (
          nx7556)) ;
    mux21 L1_0_L2_0_G1_MINI_ALU_ix241 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_5), .A0 (
          L1_0_L2_0_G1_MINI_ALU_nx419), .A1 (L1_0_L2_0_G1_MINI_ALU_nx421), .S0 (
          nx7556)) ;
    mux21 L1_0_L2_0_G1_MINI_ALU_ix261 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_6), .A0 (
          L1_0_L2_0_G1_MINI_ALU_nx429), .A1 (L1_0_L2_0_G1_MINI_ALU_nx431), .S0 (
          nx7556)) ;
    mux21 L1_0_L2_0_G1_MINI_ALU_ix281 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_7), .A0 (
          L1_0_L2_0_G1_MINI_ALU_nx439), .A1 (L1_0_L2_0_G1_MINI_ALU_nx441), .S0 (
          nx7556)) ;
    mux21 L1_0_L2_0_G1_MINI_ALU_ix301 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_8), .A0 (
          L1_0_L2_0_G1_MINI_ALU_nx449), .A1 (L1_0_L2_0_G1_MINI_ALU_nx451), .S0 (
          nx7558)) ;
    mux21 L1_0_L2_0_G1_MINI_ALU_ix321 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_9), .A0 (
          L1_0_L2_0_G1_MINI_ALU_nx469), .A1 (nx1384), .S0 (nx7558)) ;
    inv01 ix1383 (.Y (nx1384), .A (L1_0_L2_0_G1_MINI_ALU_nx316)) ;
    mux21 L1_0_L2_0_G1_MINI_ALU_ix341 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_10), .A0 (
          L1_0_L2_0_G1_MINI_ALU_nx477), .A1 (nx1386), .S0 (nx7558)) ;
    inv01 ix1385 (.Y (nx1386), .A (L1_0_L2_0_G1_MINI_ALU_nx336)) ;
    mux21 L1_0_L2_0_G1_MINI_ALU_ix361 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_11), .A0 (
          L1_0_L2_0_G1_MINI_ALU_nx485), .A1 (nx1388), .S0 (nx7558)) ;
    inv01 ix1387 (.Y (nx1388), .A (L1_0_L2_0_G1_MINI_ALU_nx356)) ;
    mux21 L1_0_L2_0_G1_MINI_ALU_ix381 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_12), .A0 (
          L1_0_L2_0_G1_MINI_ALU_nx493), .A1 (nx1390), .S0 (nx7558)) ;
    inv01 ix1389 (.Y (nx1390), .A (L1_0_L2_0_G1_MINI_ALU_nx376)) ;
    mux21 L1_0_L2_0_G1_MINI_ALU_ix401 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_13), .A0 (
          L1_0_L2_0_G1_MINI_ALU_nx501), .A1 (nx1392), .S0 (nx7558)) ;
    inv01 ix1391 (.Y (nx1392), .A (L1_0_L2_0_G1_MINI_ALU_nx396)) ;
    mux21 L1_0_L2_0_G1_MINI_ALU_ix421 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_14), .A0 (
          L1_0_L2_0_G1_MINI_ALU_nx509), .A1 (nx1394), .S0 (nx7558)) ;
    inv01 ix1393 (.Y (nx1394), .A (L1_0_L2_0_G1_MINI_ALU_nx416)) ;
    mux21 L1_0_L2_0_G1_MINI_ALU_ix441 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_15), .A0 (
          L1_0_L2_0_G1_MINI_ALU_nx517), .A1 (nx1396), .S0 (nx7560)) ;
    inv01 ix1395 (.Y (nx1396), .A (L1_0_L2_0_G1_MINI_ALU_nx436)) ;
    mux21 L1_0_L2_0_G1_MINI_ALU_ix461 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_16), .A0 (nx1398), .A1 (nx1400
          ), .S0 (nx7560)) ;
    inv01 ix1397 (.Y (nx1398), .A (L1_0_L2_0_G1_MINI_ALU_BoothP_16)) ;
    inv01 ix1399 (.Y (nx1400), .A (L1_0_L2_0_G1_MINI_ALU_nx456)) ;
    nor02_2x L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix319 (.Y (
             L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642), .A0 (Start), .A1 (
             CalculatingBooth_dup_1084)) ;
    nor02_2x L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix85 (.Y (
             L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_0), .A0 (nx7570), .A1 (
             nx1402)) ;
    inv01 ix1401 (.Y (nx1402), .A (L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_1)) ;
    mux21 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix125 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_1), .A0 (nx1404), .A1 (
          nx1406), .S0 (nx7570)) ;
    inv01 ix1403 (.Y (nx1404), .A (L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_2)) ;
    inv01 ix1405 (.Y (nx1406), .A (WindowDin_0__0__0)) ;
    mux21 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix133 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_2), .A0 (nx1408), .A1 (
          nx1410), .S0 (nx7570)) ;
    inv01 ix1407 (.Y (nx1408), .A (L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_3)) ;
    inv01 ix1409 (.Y (nx1410), .A (WindowDin_0__0__1)) ;
    mux21 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix141 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_3), .A0 (nx1412), .A1 (
          nx1414), .S0 (nx7570)) ;
    inv01 ix1411 (.Y (nx1412), .A (L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_4)) ;
    inv01 ix1413 (.Y (nx1414), .A (WindowDin_0__0__2)) ;
    mux21 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix149 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_4), .A0 (nx1416), .A1 (
          nx1418), .S0 (nx7570)) ;
    inv01 ix1415 (.Y (nx1416), .A (L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_5)) ;
    inv01 ix1417 (.Y (nx1418), .A (WindowDin_0__0__3)) ;
    mux21 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix157 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_5), .A0 (nx1420), .A1 (
          nx1422), .S0 (nx7570)) ;
    inv01 ix1419 (.Y (nx1420), .A (L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_6)) ;
    inv01 ix1421 (.Y (nx1422), .A (WindowDin_0__0__4)) ;
    mux21 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix165 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_6), .A0 (nx1424), .A1 (
          nx1426), .S0 (nx7570)) ;
    inv01 ix1423 (.Y (nx1424), .A (L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_7)) ;
    inv01 ix1425 (.Y (nx1426), .A (WindowDin_0__0__5)) ;
    mux21 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix173 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_7), .A0 (nx1428), .A1 (
          nx1430), .S0 (nx7572)) ;
    inv01 ix1427 (.Y (nx1428), .A (L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_8)) ;
    inv01 ix1429 (.Y (nx1430), .A (WindowDin_0__0__6)) ;
    mux21 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix181 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_8), .A0 (nx1432), .A1 (
          nx1434), .S0 (nx7572)) ;
    inv01 ix1431 (.Y (nx1432), .A (L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_9)) ;
    inv01 ix1433 (.Y (nx1434), .A (WindowDin_0__0__7)) ;
    nor02_2x L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix89 (.Y (
             L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_9), .A0 (nx7572), .A1 (
             nx1436)) ;
    inv01 ix1435 (.Y (nx1436), .A (L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_10)
          ) ;
    nor02_2x L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix93 (.Y (
             L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_10), .A0 (nx7572), .A1 (
             nx1438)) ;
    inv01 ix1437 (.Y (nx1438), .A (L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_11)
          ) ;
    nor02_2x L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix97 (.Y (
             L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_11), .A0 (nx7572), .A1 (
             nx1440)) ;
    inv01 ix1439 (.Y (nx1440), .A (L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_12)
          ) ;
    nor02_2x L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix101 (.Y (
             L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_12), .A0 (nx7572), .A1 (
             nx1442)) ;
    inv01 ix1441 (.Y (nx1442), .A (L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_13)
          ) ;
    nor02_2x L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix105 (.Y (
             L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_13), .A0 (nx7572), .A1 (
             nx1444)) ;
    inv01 ix1443 (.Y (nx1444), .A (L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_14)
          ) ;
    nor02_2x L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix109 (.Y (
             L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_14), .A0 (nx7574), .A1 (
             nx1446)) ;
    inv01 ix1445 (.Y (nx1446), .A (L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_15)
          ) ;
    nor02_2x L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix113 (.Y (
             L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_15), .A0 (nx7574), .A1 (
             nx1448)) ;
    inv01 ix1447 (.Y (nx1448), .A (L1_0_L2_0_G1_MINI_ALU_BoothPBeforeShift_16)
          ) ;
    nor02_2x L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix117 (.Y (
             L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_16), .A0 (nx7574), .A1 (
             nx1448)) ;
    mux21 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix189 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BoothOperand_0), .A0 (nx1450), .A1 (nx1452), .S0 (
          nx7562)) ;
    inv01 ix1449 (.Y (nx1450), .A (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_0)) ;
    inv01 ix1451 (.Y (nx1452), .A (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_0)) ;
    mux21 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix197 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BoothOperand_1), .A0 (nx1454), .A1 (nx1456), .S0 (
          nx7562)) ;
    inv01 ix1453 (.Y (nx1454), .A (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_1)) ;
    inv01 ix1455 (.Y (nx1456), .A (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_1)) ;
    mux21 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix205 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BoothOperand_2), .A0 (nx1458), .A1 (nx1460), .S0 (
          nx7562)) ;
    inv01 ix1457 (.Y (nx1458), .A (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_2)) ;
    inv01 ix1459 (.Y (nx1460), .A (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_2)) ;
    mux21 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix213 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BoothOperand_3), .A0 (nx1462), .A1 (nx1464), .S0 (
          nx7562)) ;
    inv01 ix1461 (.Y (nx1462), .A (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_3)) ;
    inv01 ix1463 (.Y (nx1464), .A (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_3)) ;
    mux21 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix221 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BoothOperand_4), .A0 (nx1466), .A1 (nx1468), .S0 (
          nx7562)) ;
    inv01 ix1465 (.Y (nx1466), .A (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_4)) ;
    inv01 ix1467 (.Y (nx1468), .A (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_4)) ;
    mux21 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix229 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BoothOperand_5), .A0 (nx1470), .A1 (nx1472), .S0 (
          nx7564)) ;
    inv01 ix1469 (.Y (nx1470), .A (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_5)) ;
    inv01 ix1471 (.Y (nx1472), .A (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_5)) ;
    mux21 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix237 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BoothOperand_6), .A0 (nx1474), .A1 (nx1476), .S0 (
          nx7564)) ;
    inv01 ix1473 (.Y (nx1474), .A (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_6)) ;
    inv01 ix1475 (.Y (nx1476), .A (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_6)) ;
    mux21 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix245 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BoothOperand_7), .A0 (nx1478), .A1 (nx1480), .S0 (
          nx7564)) ;
    inv01 ix1477 (.Y (nx1478), .A (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_7)) ;
    inv01 ix1479 (.Y (nx1480), .A (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_7)) ;
    mux21 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix253 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BoothOperand_8), .A0 (nx1482), .A1 (nx1484), .S0 (
          nx7564)) ;
    inv01 ix1481 (.Y (nx1482), .A (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_8)) ;
    inv01 ix1483 (.Y (nx1484), .A (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_8)) ;
    mux21 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix261 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BoothOperand_9), .A0 (nx1486), .A1 (nx1488), .S0 (
          nx7564)) ;
    inv01 ix1485 (.Y (nx1486), .A (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_9)) ;
    inv01 ix1487 (.Y (nx1488), .A (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_9)) ;
    mux21 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix269 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BoothOperand_10), .A0 (nx1490), .A1 (nx1492), .S0 (
          nx7564)) ;
    inv01 ix1489 (.Y (nx1490), .A (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_10)) ;
    inv01 ix1491 (.Y (nx1492), .A (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_10)) ;
    mux21 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix277 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BoothOperand_11), .A0 (nx1494), .A1 (nx1496), .S0 (
          nx7564)) ;
    inv01 ix1493 (.Y (nx1494), .A (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_11)) ;
    inv01 ix1495 (.Y (nx1496), .A (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_11)) ;
    mux21 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix285 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BoothOperand_12), .A0 (nx1498), .A1 (nx1500), .S0 (
          nx7566)) ;
    inv01 ix1497 (.Y (nx1498), .A (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_12)) ;
    inv01 ix1499 (.Y (nx1500), .A (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_12)) ;
    mux21 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix293 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BoothOperand_13), .A0 (nx1502), .A1 (nx1504), .S0 (
          nx7566)) ;
    inv01 ix1501 (.Y (nx1502), .A (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_13)) ;
    inv01 ix1503 (.Y (nx1504), .A (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_13)) ;
    mux21 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix301 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BoothOperand_14), .A0 (nx1506), .A1 (nx1508), .S0 (
          nx7566)) ;
    inv01 ix1505 (.Y (nx1506), .A (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_14)) ;
    inv01 ix1507 (.Y (nx1508), .A (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_14)) ;
    mux21 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix309 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BoothOperand_15), .A0 (nx1510), .A1 (nx1512), .S0 (
          nx7566)) ;
    inv01 ix1509 (.Y (nx1510), .A (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_15)) ;
    inv01 ix1511 (.Y (nx1512), .A (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_15)) ;
    mux21 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix317 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BoothOperand_16), .A0 (nx1514), .A1 (nx1516), .S0 (
          nx7566)) ;
    inv01 ix1513 (.Y (nx1514), .A (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_16)) ;
    inv01 ix1515 (.Y (nx1516), .A (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_16)) ;
    xnor2 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix321 (.Y (
          L1_0_L2_0_G1_MINI_ALU_AddPToBoothOperand), .A0 (nx7566), .A1 (nx1382)
          ) ;
    oai32 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix393 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .A0 (nx8596), .A1 (
          RST), .A2 (nx7618), .B0 (nx1452), .B1 (nx1520)) ;
    oai32 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix403 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .A0 (nx8596), .A1 (
          RST), .A2 (nx7618), .B0 (nx1456), .B1 (nx1520)) ;
    oai32 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix413 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .A0 (nx8596), .A1 (
          RST), .A2 (nx7618), .B0 (nx1460), .B1 (nx1520)) ;
    oai32 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix423 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .A0 (nx8596), .A1 (
          RST), .A2 (nx7618), .B0 (nx1464), .B1 (nx1520)) ;
    oai32 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix433 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .A0 (nx8596), .A1 (
          RST), .A2 (nx7618), .B0 (nx1468), .B1 (nx1520)) ;
    oai32 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix443 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .A0 (nx8596), .A1 (
          RST), .A2 (nx7618), .B0 (nx1472), .B1 (nx1520)) ;
    oai32 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix453 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .A0 (nx8596), .A1 (
          RST), .A2 (nx7620), .B0 (nx1476), .B1 (nx1520)) ;
    oai32 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix463 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .A0 (nx8598), .A1 (
          RST), .A2 (nx7620), .B0 (nx1480), .B1 (nx1522)) ;
    oai32 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix473 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .A0 (nx8598), .A1 (
          RST), .A2 (nx7620), .B0 (nx1484), .B1 (nx1522)) ;
    oai32 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix483 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .A0 (nx1524), .A1 (
          RST), .A2 (nx7620), .B0 (nx1488), .B1 (nx1522)) ;
    inv01 ix1523 (.Y (nx1524), .A (FilterDin_0__0__0)) ;
    oai32 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix493 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .A0 (nx1526), .A1 (
          RST), .A2 (nx7620), .B0 (nx1492), .B1 (nx1522)) ;
    inv01 ix1525 (.Y (nx1526), .A (FilterDin_0__0__1)) ;
    oai32 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix503 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .A0 (nx1528), .A1 (
          RST), .A2 (nx7620), .B0 (nx1496), .B1 (nx1522)) ;
    inv01 ix1527 (.Y (nx1528), .A (FilterDin_0__0__2)) ;
    oai32 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix513 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .A0 (nx1530), .A1 (
          RST), .A2 (nx7620), .B0 (nx1500), .B1 (nx1522)) ;
    inv01 ix1529 (.Y (nx1530), .A (FilterDin_0__0__3)) ;
    oai32 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix523 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .A0 (nx1532), .A1 (
          RST), .A2 (nx7622), .B0 (nx1504), .B1 (nx1522)) ;
    inv01 ix1531 (.Y (nx1532), .A (FilterDin_0__0__4)) ;
    oai32 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix533 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .A0 (nx1534), .A1 (
          RST), .A2 (nx7622), .B0 (nx1508), .B1 (nx1536)) ;
    inv01 ix1533 (.Y (nx1534), .A (FilterDin_0__0__5)) ;
    inv01 ix1535 (.Y (nx1536), .A (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566)) ;
    oai32 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix543 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .A0 (nx1538), .A1 (
          RST), .A2 (nx7622), .B0 (nx1512), .B1 (nx1536)) ;
    inv01 ix1537 (.Y (nx1538), .A (FilterDin_0__0__6)) ;
    oai32 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix553 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .A0 (nx1540), .A1 (
          RST), .A2 (nx7622), .B0 (nx1516), .B1 (nx1536)) ;
    inv01 ix1539 (.Y (nx1540), .A (FilterDin_0__0__7)) ;
    nand02_2x L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix633 (.Y (nx1520), .A0 (
              nx7576), .A1 (nx7622)) ;
    nand02_2x L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix635 (.Y (nx1522), .A0 (
              nx7576), .A1 (nx7622)) ;
    oai32 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix393 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .A0 (nx8598), .A1 (
          RST), .A2 (nx7624), .B0 (nx1450), .B1 (nx1542)) ;
    oai32 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix403 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .A0 (nx8598), .A1 (
          RST), .A2 (nx7624), .B0 (nx1454), .B1 (nx1542)) ;
    oai32 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix413 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .A0 (nx8598), .A1 (
          RST), .A2 (nx7624), .B0 (nx1458), .B1 (nx1542)) ;
    oai32 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix423 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .A0 (nx8598), .A1 (
          RST), .A2 (nx7624), .B0 (nx1462), .B1 (nx1542)) ;
    oai32 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix433 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .A0 (nx8598), .A1 (
          RST), .A2 (nx7624), .B0 (nx1466), .B1 (nx1542)) ;
    oai32 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix443 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .A0 (nx8600), .A1 (
          RST), .A2 (nx7624), .B0 (nx1470), .B1 (nx1542)) ;
    oai32 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix453 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .A0 (nx8600), .A1 (
          RST), .A2 (nx7626), .B0 (nx1474), .B1 (nx1542)) ;
    oai32 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix463 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .A0 (nx8600), .A1 (
          RST), .A2 (nx7626), .B0 (nx1478), .B1 (nx1544)) ;
    oai32 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix473 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .A0 (nx8600), .A1 (
          RST), .A2 (nx7626), .B0 (nx1482), .B1 (nx1544)) ;
    oai32 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix483 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .A0 (nx1524), .A1 (
          RST), .A2 (nx7626), .B0 (nx1486), .B1 (nx1544)) ;
    oai32 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix493 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .A0 (nx1546), .A1 (
          RST), .A2 (nx7626), .B0 (nx1490), .B1 (nx1544)) ;
    inv01 ix1545 (.Y (nx1546), .A (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_10)) ;
    oai32 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix503 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .A0 (nx1548), .A1 (
          RST), .A2 (nx7626), .B0 (nx1494), .B1 (nx1544)) ;
    inv01 ix1547 (.Y (nx1548), .A (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_11)) ;
    oai32 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix513 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .A0 (nx1550), .A1 (
          RST), .A2 (nx7626), .B0 (nx1498), .B1 (nx1544)) ;
    inv01 ix1549 (.Y (nx1550), .A (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_12)) ;
    oai32 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix523 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .A0 (nx1552), .A1 (
          RST), .A2 (nx7628), .B0 (nx1502), .B1 (nx1544)) ;
    inv01 ix1551 (.Y (nx1552), .A (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_13)) ;
    oai32 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix533 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .A0 (nx1554), .A1 (
          RST), .A2 (nx7628), .B0 (nx1506), .B1 (nx1556)) ;
    inv01 ix1553 (.Y (nx1554), .A (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_14)) ;
    inv01 ix1555 (.Y (nx1556), .A (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566)) ;
    oai32 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix543 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .A0 (nx1558), .A1 (
          RST), .A2 (nx7628), .B0 (nx1510), .B1 (nx1556)) ;
    inv01 ix1557 (.Y (nx1558), .A (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_15)) ;
    oai32 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix553 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .A0 (nx1560), .A1 (
          RST), .A2 (nx7628), .B0 (nx1514), .B1 (nx1556)) ;
    inv01 ix1559 (.Y (nx1560), .A (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_16)) ;
    nand02_2x L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix633 (.Y (nx1542), .A0 (
              nx7576), .A1 (nx7628)) ;
    nand02_2x L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix635 (.Y (nx1544), .A0 (
              nx7576), .A1 (nx7628)) ;
    oai32 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix393 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .A0 (nx1562), .A1 (
          RST), .A2 (nx7630), .B0 (L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx384), .B1 (
          nx1564)) ;
    inv01 ix1561 (.Y (nx1562), .A (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_0)) ;
    oai32 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix403 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .A0 (nx1566), .A1 (
          RST), .A2 (nx7630), .B0 (nx1382), .B1 (nx1564)) ;
    inv01 ix1565 (.Y (nx1566), .A (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_1)) ;
    oai32 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix413 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .A0 (nx1568), .A1 (
          RST), .A2 (nx7630), .B0 (L1_0_L2_0_G1_MINI_ALU_nx387), .B1 (nx1564)) ;
    inv01 ix1567 (.Y (nx1568), .A (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_2)) ;
    oai32 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix423 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .A0 (nx1570), .A1 (
          RST), .A2 (nx7630), .B0 (L1_0_L2_0_G1_MINI_ALU_nx399), .B1 (nx1564)) ;
    inv01 ix1569 (.Y (nx1570), .A (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_3)) ;
    oai32 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix433 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .A0 (nx1572), .A1 (
          RST), .A2 (nx7630), .B0 (L1_0_L2_0_G1_MINI_ALU_nx409), .B1 (nx1564)) ;
    inv01 ix1571 (.Y (nx1572), .A (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_4)) ;
    oai32 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix443 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .A0 (nx1574), .A1 (
          RST), .A2 (nx7630), .B0 (L1_0_L2_0_G1_MINI_ALU_nx419), .B1 (nx1564)) ;
    inv01 ix1573 (.Y (nx1574), .A (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_5)) ;
    oai32 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix453 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .A0 (nx1576), .A1 (
          RST), .A2 (nx7630), .B0 (L1_0_L2_0_G1_MINI_ALU_nx429), .B1 (nx1564)) ;
    inv01 ix1575 (.Y (nx1576), .A (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_6)) ;
    oai32 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix463 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .A0 (nx1578), .A1 (
          RST), .A2 (nx7632), .B0 (L1_0_L2_0_G1_MINI_ALU_nx439), .B1 (nx1580)) ;
    inv01 ix1577 (.Y (nx1578), .A (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_7)) ;
    oai32 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix473 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .A0 (nx1582), .A1 (
          RST), .A2 (nx7632), .B0 (L1_0_L2_0_G1_MINI_ALU_nx449), .B1 (nx1580)) ;
    inv01 ix1581 (.Y (nx1582), .A (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_8)) ;
    oai32 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix483 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .A0 (nx1584), .A1 (
          RST), .A2 (nx7632), .B0 (L1_0_L2_0_G1_MINI_ALU_nx469), .B1 (nx1580)) ;
    inv01 ix1583 (.Y (nx1584), .A (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_9)) ;
    oai32 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix493 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .A0 (nx1586), .A1 (
          RST), .A2 (nx7632), .B0 (L1_0_L2_0_G1_MINI_ALU_nx477), .B1 (nx1580)) ;
    inv01 ix1585 (.Y (nx1586), .A (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_10)) ;
    oai32 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix503 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .A0 (nx1588), .A1 (
          RST), .A2 (nx7632), .B0 (L1_0_L2_0_G1_MINI_ALU_nx485), .B1 (nx1580)) ;
    inv01 ix1587 (.Y (nx1588), .A (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_11)) ;
    oai32 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix513 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .A0 (nx1590), .A1 (
          RST), .A2 (nx7632), .B0 (L1_0_L2_0_G1_MINI_ALU_nx493), .B1 (nx1580)) ;
    inv01 ix1589 (.Y (nx1590), .A (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_12)) ;
    oai32 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix523 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .A0 (nx1592), .A1 (
          RST), .A2 (nx7632), .B0 (L1_0_L2_0_G1_MINI_ALU_nx501), .B1 (nx1580)) ;
    inv01 ix1591 (.Y (nx1592), .A (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_13)) ;
    oai32 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix533 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .A0 (nx1594), .A1 (
          RST), .A2 (nx7634), .B0 (L1_0_L2_0_G1_MINI_ALU_nx509), .B1 (nx1596)) ;
    inv01 ix1593 (.Y (nx1594), .A (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_14)) ;
    inv01 ix1595 (.Y (nx1596), .A (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566)) ;
    oai32 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix543 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .A0 (nx1598), .A1 (
          RST), .A2 (nx7634), .B0 (L1_0_L2_0_G1_MINI_ALU_nx517), .B1 (nx1596)) ;
    inv01 ix1597 (.Y (nx1598), .A (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_15)) ;
    oai32 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix553 (.Y (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .A0 (nx1600), .A1 (
          RST), .A2 (nx7634), .B0 (nx1398), .B1 (nx1596)) ;
    inv01 ix1599 (.Y (nx1600), .A (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_16)) ;
    nand02_2x L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix633 (.Y (nx1564), .A0 (
              nx7576), .A1 (nx7634)) ;
    nand02_2x L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix635 (.Y (nx1580), .A0 (
              nx7576), .A1 (nx7634)) ;
    mux21 L1_0_L2_1_G1_MINI_ALU_ix404 (.Y (L1_0_L2_1_G1_MINI_ALU_nx403), .A0 (
          nx1602), .A1 (L1_0_L2_1_G1_MINI_ALU_BoothP_2), .S0 (
          L1_0_L2_1_G1_MINI_ALU_nx395)) ;
    inv01 ix1601 (.Y (nx1602), .A (L1_0_L2_1_G1_MINI_ALU_nx391)) ;
    mux21 L1_0_L2_1_G1_MINI_ALU_ix414 (.Y (L1_0_L2_1_G1_MINI_ALU_nx413), .A0 (
          nx1604), .A1 (L1_0_L2_1_G1_MINI_ALU_BoothP_3), .S0 (
          L1_0_L2_1_G1_MINI_ALU_nx405)) ;
    inv01 ix1603 (.Y (nx1604), .A (L1_0_L2_1_G1_MINI_ALU_nx403)) ;
    mux21 L1_0_L2_1_G1_MINI_ALU_ix424 (.Y (L1_0_L2_1_G1_MINI_ALU_nx423), .A0 (
          nx1606), .A1 (L1_0_L2_1_G1_MINI_ALU_BoothP_4), .S0 (
          L1_0_L2_1_G1_MINI_ALU_nx415)) ;
    inv01 ix1605 (.Y (nx1606), .A (L1_0_L2_1_G1_MINI_ALU_nx413)) ;
    mux21 L1_0_L2_1_G1_MINI_ALU_ix434 (.Y (L1_0_L2_1_G1_MINI_ALU_nx433), .A0 (
          nx1608), .A1 (L1_0_L2_1_G1_MINI_ALU_BoothP_5), .S0 (
          L1_0_L2_1_G1_MINI_ALU_nx425)) ;
    inv01 ix1607 (.Y (nx1608), .A (L1_0_L2_1_G1_MINI_ALU_nx423)) ;
    mux21 L1_0_L2_1_G1_MINI_ALU_ix444 (.Y (L1_0_L2_1_G1_MINI_ALU_nx443), .A0 (
          nx1610), .A1 (L1_0_L2_1_G1_MINI_ALU_BoothP_6), .S0 (
          L1_0_L2_1_G1_MINI_ALU_nx435)) ;
    inv01 ix1609 (.Y (nx1610), .A (L1_0_L2_1_G1_MINI_ALU_nx433)) ;
    mux21 L1_0_L2_1_G1_MINI_ALU_ix454 (.Y (L1_0_L2_1_G1_MINI_ALU_nx453), .A0 (
          nx1612), .A1 (L1_0_L2_1_G1_MINI_ALU_BoothP_7), .S0 (
          L1_0_L2_1_G1_MINI_ALU_nx445)) ;
    inv01 ix1611 (.Y (nx1612), .A (L1_0_L2_1_G1_MINI_ALU_nx443)) ;
    mux21 L1_0_L2_1_G1_MINI_ALU_ix462 (.Y (L1_0_L2_1_G1_MINI_ALU_nx461), .A0 (
          nx1614), .A1 (L1_0_L2_1_G1_MINI_ALU_BoothP_8), .S0 (
          L1_0_L2_1_G1_MINI_ALU_nx455)) ;
    inv01 ix1613 (.Y (nx1614), .A (L1_0_L2_1_G1_MINI_ALU_nx453)) ;
    mux21 L1_0_L2_1_G1_MINI_ALU_ix468 (.Y (L1_0_L2_1_G1_MINI_ALU_nx467), .A0 (
          nx1616), .A1 (L1_0_L2_1_G1_MINI_ALU_BoothP_9), .S0 (
          L1_0_L2_1_G1_MINI_ALU_nx463)) ;
    inv01 ix1615 (.Y (nx1616), .A (L1_0_L2_1_G1_MINI_ALU_nx461)) ;
    mux21 L1_0_L2_1_G1_MINI_ALU_ix476 (.Y (L1_0_L2_1_G1_MINI_ALU_nx475), .A0 (
          nx1618), .A1 (L1_0_L2_1_G1_MINI_ALU_BoothP_10), .S0 (
          L1_0_L2_1_G1_MINI_ALU_nx471)) ;
    inv01 ix1617 (.Y (nx1618), .A (L1_0_L2_1_G1_MINI_ALU_nx467)) ;
    mux21 L1_0_L2_1_G1_MINI_ALU_ix484 (.Y (L1_0_L2_1_G1_MINI_ALU_nx483), .A0 (
          nx1620), .A1 (L1_0_L2_1_G1_MINI_ALU_BoothP_11), .S0 (
          L1_0_L2_1_G1_MINI_ALU_nx479)) ;
    inv01 ix1619 (.Y (nx1620), .A (L1_0_L2_1_G1_MINI_ALU_nx475)) ;
    mux21 L1_0_L2_1_G1_MINI_ALU_ix492 (.Y (L1_0_L2_1_G1_MINI_ALU_nx491), .A0 (
          nx1622), .A1 (L1_0_L2_1_G1_MINI_ALU_BoothP_12), .S0 (
          L1_0_L2_1_G1_MINI_ALU_nx487)) ;
    inv01 ix1621 (.Y (nx1622), .A (L1_0_L2_1_G1_MINI_ALU_nx483)) ;
    mux21 L1_0_L2_1_G1_MINI_ALU_ix500 (.Y (L1_0_L2_1_G1_MINI_ALU_nx499), .A0 (
          nx1624), .A1 (L1_0_L2_1_G1_MINI_ALU_BoothP_13), .S0 (
          L1_0_L2_1_G1_MINI_ALU_nx495)) ;
    inv01 ix1623 (.Y (nx1624), .A (L1_0_L2_1_G1_MINI_ALU_nx491)) ;
    mux21 L1_0_L2_1_G1_MINI_ALU_ix508 (.Y (L1_0_L2_1_G1_MINI_ALU_nx507), .A0 (
          nx1626), .A1 (L1_0_L2_1_G1_MINI_ALU_BoothP_14), .S0 (
          L1_0_L2_1_G1_MINI_ALU_nx503)) ;
    inv01 ix1625 (.Y (nx1626), .A (L1_0_L2_1_G1_MINI_ALU_nx499)) ;
    mux21 L1_0_L2_1_G1_MINI_ALU_ix516 (.Y (L1_0_L2_1_G1_MINI_ALU_nx515), .A0 (
          nx1628), .A1 (L1_0_L2_1_G1_MINI_ALU_BoothP_15), .S0 (
          L1_0_L2_1_G1_MINI_ALU_nx511)) ;
    inv01 ix1627 (.Y (nx1628), .A (L1_0_L2_1_G1_MINI_ALU_nx507)) ;
    mux21 L1_0_L2_1_G1_MINI_ALU_ix161 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_1), .A0 (nx1630), .A1 (
          L1_0_L2_1_G1_MINI_ALU_nx379), .S0 (nx7638)) ;
    inv01 ix1629 (.Y (nx1630), .A (L1_0_L2_1_G1_MINI_ALU_BoothP_1)) ;
    mux21 L1_0_L2_1_G1_MINI_ALU_ix181 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_2), .A0 (
          L1_0_L2_1_G1_MINI_ALU_nx387), .A1 (L1_0_L2_1_G1_MINI_ALU_nx389), .S0 (
          nx7638)) ;
    mux21 L1_0_L2_1_G1_MINI_ALU_ix201 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_3), .A0 (
          L1_0_L2_1_G1_MINI_ALU_nx399), .A1 (L1_0_L2_1_G1_MINI_ALU_nx401), .S0 (
          nx7638)) ;
    mux21 L1_0_L2_1_G1_MINI_ALU_ix221 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_4), .A0 (
          L1_0_L2_1_G1_MINI_ALU_nx409), .A1 (L1_0_L2_1_G1_MINI_ALU_nx411), .S0 (
          nx7638)) ;
    mux21 L1_0_L2_1_G1_MINI_ALU_ix241 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_5), .A0 (
          L1_0_L2_1_G1_MINI_ALU_nx419), .A1 (L1_0_L2_1_G1_MINI_ALU_nx421), .S0 (
          nx7638)) ;
    mux21 L1_0_L2_1_G1_MINI_ALU_ix261 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_6), .A0 (
          L1_0_L2_1_G1_MINI_ALU_nx429), .A1 (L1_0_L2_1_G1_MINI_ALU_nx431), .S0 (
          nx7638)) ;
    mux21 L1_0_L2_1_G1_MINI_ALU_ix281 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_7), .A0 (
          L1_0_L2_1_G1_MINI_ALU_nx439), .A1 (L1_0_L2_1_G1_MINI_ALU_nx441), .S0 (
          nx7638)) ;
    mux21 L1_0_L2_1_G1_MINI_ALU_ix301 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_8), .A0 (
          L1_0_L2_1_G1_MINI_ALU_nx449), .A1 (L1_0_L2_1_G1_MINI_ALU_nx451), .S0 (
          nx7640)) ;
    mux21 L1_0_L2_1_G1_MINI_ALU_ix321 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_9), .A0 (
          L1_0_L2_1_G1_MINI_ALU_nx469), .A1 (nx1632), .S0 (nx7640)) ;
    inv01 ix1631 (.Y (nx1632), .A (L1_0_L2_1_G1_MINI_ALU_nx316)) ;
    mux21 L1_0_L2_1_G1_MINI_ALU_ix341 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_10), .A0 (
          L1_0_L2_1_G1_MINI_ALU_nx477), .A1 (nx1634), .S0 (nx7640)) ;
    inv01 ix1633 (.Y (nx1634), .A (L1_0_L2_1_G1_MINI_ALU_nx336)) ;
    mux21 L1_0_L2_1_G1_MINI_ALU_ix361 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_11), .A0 (
          L1_0_L2_1_G1_MINI_ALU_nx485), .A1 (nx1636), .S0 (nx7640)) ;
    inv01 ix1635 (.Y (nx1636), .A (L1_0_L2_1_G1_MINI_ALU_nx356)) ;
    mux21 L1_0_L2_1_G1_MINI_ALU_ix381 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_12), .A0 (
          L1_0_L2_1_G1_MINI_ALU_nx493), .A1 (nx1638), .S0 (nx7640)) ;
    inv01 ix1637 (.Y (nx1638), .A (L1_0_L2_1_G1_MINI_ALU_nx376)) ;
    mux21 L1_0_L2_1_G1_MINI_ALU_ix401 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_13), .A0 (
          L1_0_L2_1_G1_MINI_ALU_nx501), .A1 (nx1640), .S0 (nx7640)) ;
    inv01 ix1639 (.Y (nx1640), .A (L1_0_L2_1_G1_MINI_ALU_nx396)) ;
    mux21 L1_0_L2_1_G1_MINI_ALU_ix421 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_14), .A0 (
          L1_0_L2_1_G1_MINI_ALU_nx509), .A1 (nx1642), .S0 (nx7640)) ;
    inv01 ix1641 (.Y (nx1642), .A (L1_0_L2_1_G1_MINI_ALU_nx416)) ;
    mux21 L1_0_L2_1_G1_MINI_ALU_ix441 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_15), .A0 (
          L1_0_L2_1_G1_MINI_ALU_nx517), .A1 (nx1644), .S0 (nx7642)) ;
    inv01 ix1643 (.Y (nx1644), .A (L1_0_L2_1_G1_MINI_ALU_nx436)) ;
    mux21 L1_0_L2_1_G1_MINI_ALU_ix461 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_16), .A0 (nx1646), .A1 (nx1648
          ), .S0 (nx7642)) ;
    inv01 ix1645 (.Y (nx1646), .A (L1_0_L2_1_G1_MINI_ALU_BoothP_16)) ;
    inv01 ix1647 (.Y (nx1648), .A (L1_0_L2_1_G1_MINI_ALU_nx456)) ;
    nor02_2x L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix319 (.Y (
             L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642), .A0 (Start), .A1 (
             CalculatingBooth_dup_1084)) ;
    nor02_2x L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix85 (.Y (
             L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_0), .A0 (nx7652), .A1 (
             nx1650)) ;
    inv01 ix1649 (.Y (nx1650), .A (L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_1)) ;
    mux21 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix125 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_1), .A0 (nx1652), .A1 (
          nx1654), .S0 (nx7652)) ;
    inv01 ix1651 (.Y (nx1652), .A (L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_2)) ;
    inv01 ix1653 (.Y (nx1654), .A (WindowDin_0__1__0)) ;
    mux21 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix133 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_2), .A0 (nx1656), .A1 (
          nx1658), .S0 (nx7652)) ;
    inv01 ix1655 (.Y (nx1656), .A (L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_3)) ;
    inv01 ix1657 (.Y (nx1658), .A (WindowDin_0__1__1)) ;
    mux21 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix141 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_3), .A0 (nx1660), .A1 (
          nx1662), .S0 (nx7652)) ;
    inv01 ix1659 (.Y (nx1660), .A (L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_4)) ;
    inv01 ix1661 (.Y (nx1662), .A (WindowDin_0__1__2)) ;
    mux21 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix149 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_4), .A0 (nx1664), .A1 (
          nx1666), .S0 (nx7652)) ;
    inv01 ix1663 (.Y (nx1664), .A (L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_5)) ;
    inv01 ix1665 (.Y (nx1666), .A (WindowDin_0__1__3)) ;
    mux21 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix157 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_5), .A0 (nx1668), .A1 (
          nx1670), .S0 (nx7652)) ;
    inv01 ix1667 (.Y (nx1668), .A (L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_6)) ;
    inv01 ix1669 (.Y (nx1670), .A (WindowDin_0__1__4)) ;
    mux21 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix165 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_6), .A0 (nx1672), .A1 (
          nx1674), .S0 (nx7652)) ;
    inv01 ix1671 (.Y (nx1672), .A (L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_7)) ;
    inv01 ix1673 (.Y (nx1674), .A (WindowDin_0__1__5)) ;
    mux21 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix173 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_7), .A0 (nx1676), .A1 (
          nx1678), .S0 (nx7654)) ;
    inv01 ix1675 (.Y (nx1676), .A (L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_8)) ;
    inv01 ix1677 (.Y (nx1678), .A (WindowDin_0__1__6)) ;
    mux21 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix181 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_8), .A0 (nx1680), .A1 (
          nx1682), .S0 (nx7654)) ;
    inv01 ix1679 (.Y (nx1680), .A (L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_9)) ;
    inv01 ix1681 (.Y (nx1682), .A (WindowDin_0__1__7)) ;
    nor02_2x L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix89 (.Y (
             L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_9), .A0 (nx7654), .A1 (
             nx1684)) ;
    inv01 ix1683 (.Y (nx1684), .A (L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_10)
          ) ;
    nor02_2x L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix93 (.Y (
             L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_10), .A0 (nx7654), .A1 (
             nx1686)) ;
    inv01 ix1685 (.Y (nx1686), .A (L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_11)
          ) ;
    nor02_2x L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix97 (.Y (
             L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_11), .A0 (nx7654), .A1 (
             nx1688)) ;
    inv01 ix1687 (.Y (nx1688), .A (L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_12)
          ) ;
    nor02_2x L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix101 (.Y (
             L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_12), .A0 (nx7654), .A1 (
             nx1690)) ;
    inv01 ix1689 (.Y (nx1690), .A (L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_13)
          ) ;
    nor02_2x L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix105 (.Y (
             L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_13), .A0 (nx7654), .A1 (
             nx1692)) ;
    inv01 ix1691 (.Y (nx1692), .A (L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_14)
          ) ;
    nor02_2x L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix109 (.Y (
             L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_14), .A0 (nx7656), .A1 (
             nx1694)) ;
    inv01 ix1693 (.Y (nx1694), .A (L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_15)
          ) ;
    nor02_2x L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix113 (.Y (
             L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_15), .A0 (nx7656), .A1 (
             nx1696)) ;
    inv01 ix1695 (.Y (nx1696), .A (L1_0_L2_1_G1_MINI_ALU_BoothPBeforeShift_16)
          ) ;
    nor02_2x L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix117 (.Y (
             L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_16), .A0 (nx7656), .A1 (
             nx1696)) ;
    mux21 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix189 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BoothOperand_0), .A0 (nx1698), .A1 (nx1700), .S0 (
          nx7644)) ;
    inv01 ix1697 (.Y (nx1698), .A (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_0)) ;
    inv01 ix1699 (.Y (nx1700), .A (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_0)) ;
    mux21 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix197 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BoothOperand_1), .A0 (nx1702), .A1 (nx1704), .S0 (
          nx7644)) ;
    inv01 ix1701 (.Y (nx1702), .A (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_1)) ;
    inv01 ix1703 (.Y (nx1704), .A (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_1)) ;
    mux21 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix205 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BoothOperand_2), .A0 (nx1706), .A1 (nx1708), .S0 (
          nx7644)) ;
    inv01 ix1705 (.Y (nx1706), .A (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_2)) ;
    inv01 ix1707 (.Y (nx1708), .A (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_2)) ;
    mux21 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix213 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BoothOperand_3), .A0 (nx1710), .A1 (nx1712), .S0 (
          nx7644)) ;
    inv01 ix1709 (.Y (nx1710), .A (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_3)) ;
    inv01 ix1711 (.Y (nx1712), .A (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_3)) ;
    mux21 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix221 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BoothOperand_4), .A0 (nx1714), .A1 (nx1716), .S0 (
          nx7644)) ;
    inv01 ix1713 (.Y (nx1714), .A (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_4)) ;
    inv01 ix1715 (.Y (nx1716), .A (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_4)) ;
    mux21 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix229 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BoothOperand_5), .A0 (nx1718), .A1 (nx1720), .S0 (
          nx7646)) ;
    inv01 ix1717 (.Y (nx1718), .A (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_5)) ;
    inv01 ix1719 (.Y (nx1720), .A (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_5)) ;
    mux21 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix237 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BoothOperand_6), .A0 (nx1722), .A1 (nx1724), .S0 (
          nx7646)) ;
    inv01 ix1721 (.Y (nx1722), .A (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_6)) ;
    inv01 ix1723 (.Y (nx1724), .A (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_6)) ;
    mux21 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix245 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BoothOperand_7), .A0 (nx1726), .A1 (nx1728), .S0 (
          nx7646)) ;
    inv01 ix1725 (.Y (nx1726), .A (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_7)) ;
    inv01 ix1727 (.Y (nx1728), .A (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_7)) ;
    mux21 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix253 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BoothOperand_8), .A0 (nx1730), .A1 (nx1732), .S0 (
          nx7646)) ;
    inv01 ix1729 (.Y (nx1730), .A (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_8)) ;
    inv01 ix1731 (.Y (nx1732), .A (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_8)) ;
    mux21 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix261 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BoothOperand_9), .A0 (nx1734), .A1 (nx1736), .S0 (
          nx7646)) ;
    inv01 ix1733 (.Y (nx1734), .A (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_9)) ;
    inv01 ix1735 (.Y (nx1736), .A (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_9)) ;
    mux21 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix269 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BoothOperand_10), .A0 (nx1738), .A1 (nx1740), .S0 (
          nx7646)) ;
    inv01 ix1737 (.Y (nx1738), .A (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_10)) ;
    inv01 ix1739 (.Y (nx1740), .A (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_10)) ;
    mux21 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix277 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BoothOperand_11), .A0 (nx1742), .A1 (nx1744), .S0 (
          nx7646)) ;
    inv01 ix1741 (.Y (nx1742), .A (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_11)) ;
    inv01 ix1743 (.Y (nx1744), .A (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_11)) ;
    mux21 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix285 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BoothOperand_12), .A0 (nx1746), .A1 (nx1748), .S0 (
          nx7648)) ;
    inv01 ix1745 (.Y (nx1746), .A (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_12)) ;
    inv01 ix1747 (.Y (nx1748), .A (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_12)) ;
    mux21 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix293 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BoothOperand_13), .A0 (nx1750), .A1 (nx1752), .S0 (
          nx7648)) ;
    inv01 ix1749 (.Y (nx1750), .A (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_13)) ;
    inv01 ix1751 (.Y (nx1752), .A (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_13)) ;
    mux21 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix301 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BoothOperand_14), .A0 (nx1754), .A1 (nx1756), .S0 (
          nx7648)) ;
    inv01 ix1753 (.Y (nx1754), .A (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_14)) ;
    inv01 ix1755 (.Y (nx1756), .A (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_14)) ;
    mux21 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix309 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BoothOperand_15), .A0 (nx1758), .A1 (nx1760), .S0 (
          nx7648)) ;
    inv01 ix1757 (.Y (nx1758), .A (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_15)) ;
    inv01 ix1759 (.Y (nx1760), .A (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_15)) ;
    mux21 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix317 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BoothOperand_16), .A0 (nx1762), .A1 (nx1764), .S0 (
          nx7648)) ;
    inv01 ix1761 (.Y (nx1762), .A (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_16)) ;
    inv01 ix1763 (.Y (nx1764), .A (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_16)) ;
    xnor2 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix321 (.Y (
          L1_0_L2_1_G1_MINI_ALU_AddPToBoothOperand), .A0 (nx7648), .A1 (nx1630)
          ) ;
    oai32 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix393 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .A0 (nx8602), .A1 (
          RST), .A2 (nx7658), .B0 (nx1700), .B1 (nx1768)) ;
    oai32 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix403 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .A0 (nx8602), .A1 (
          RST), .A2 (nx7658), .B0 (nx1704), .B1 (nx1768)) ;
    oai32 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix413 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .A0 (nx8602), .A1 (
          RST), .A2 (nx7658), .B0 (nx1708), .B1 (nx1768)) ;
    oai32 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix423 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .A0 (nx8602), .A1 (
          RST), .A2 (nx7658), .B0 (nx1712), .B1 (nx1768)) ;
    oai32 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix433 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .A0 (nx8602), .A1 (
          RST), .A2 (nx7658), .B0 (nx1716), .B1 (nx1768)) ;
    oai32 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix443 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .A0 (nx8602), .A1 (
          RST), .A2 (nx7658), .B0 (nx1720), .B1 (nx1768)) ;
    oai32 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix453 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .A0 (nx8602), .A1 (
          RST), .A2 (nx7660), .B0 (nx1724), .B1 (nx1768)) ;
    oai32 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix463 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .A0 (nx8604), .A1 (
          RST), .A2 (nx7660), .B0 (nx1728), .B1 (nx1770)) ;
    oai32 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix473 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .A0 (nx8604), .A1 (
          RST), .A2 (nx7660), .B0 (nx1732), .B1 (nx1770)) ;
    oai32 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix483 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .A0 (nx1772), .A1 (
          RST), .A2 (nx7660), .B0 (nx1736), .B1 (nx1770)) ;
    inv01 ix1771 (.Y (nx1772), .A (FilterDin_0__1__0)) ;
    oai32 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix493 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .A0 (nx1774), .A1 (
          RST), .A2 (nx7660), .B0 (nx1740), .B1 (nx1770)) ;
    inv01 ix1773 (.Y (nx1774), .A (FilterDin_0__1__1)) ;
    oai32 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix503 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .A0 (nx1776), .A1 (
          RST), .A2 (nx7660), .B0 (nx1744), .B1 (nx1770)) ;
    inv01 ix1775 (.Y (nx1776), .A (FilterDin_0__1__2)) ;
    oai32 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix513 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .A0 (nx1778), .A1 (
          RST), .A2 (nx7660), .B0 (nx1748), .B1 (nx1770)) ;
    inv01 ix1777 (.Y (nx1778), .A (FilterDin_0__1__3)) ;
    oai32 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix523 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .A0 (nx1780), .A1 (
          RST), .A2 (nx7662), .B0 (nx1752), .B1 (nx1770)) ;
    inv01 ix1779 (.Y (nx1780), .A (FilterDin_0__1__4)) ;
    oai32 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix533 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .A0 (nx1782), .A1 (
          RST), .A2 (nx7662), .B0 (nx1756), .B1 (nx1784)) ;
    inv01 ix1781 (.Y (nx1782), .A (FilterDin_0__1__5)) ;
    inv01 ix1783 (.Y (nx1784), .A (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566)) ;
    oai32 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix543 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .A0 (nx1786), .A1 (
          RST), .A2 (nx7662), .B0 (nx1760), .B1 (nx1784)) ;
    inv01 ix1785 (.Y (nx1786), .A (FilterDin_0__1__6)) ;
    oai32 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix553 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .A0 (nx1788), .A1 (
          RST), .A2 (nx7662), .B0 (nx1764), .B1 (nx1784)) ;
    inv01 ix1787 (.Y (nx1788), .A (FilterDin_0__1__7)) ;
    nand02_2x L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix633 (.Y (nx1768), .A0 (
              nx7576), .A1 (nx7662)) ;
    nand02_2x L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix635 (.Y (nx1770), .A0 (
              nx7578), .A1 (nx7662)) ;
    oai32 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix393 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .A0 (nx8604), .A1 (
          RST), .A2 (nx7664), .B0 (nx1698), .B1 (nx1790)) ;
    oai32 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix403 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .A0 (nx8604), .A1 (
          RST), .A2 (nx7664), .B0 (nx1702), .B1 (nx1790)) ;
    oai32 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix413 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .A0 (nx8604), .A1 (
          RST), .A2 (nx7664), .B0 (nx1706), .B1 (nx1790)) ;
    oai32 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix423 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .A0 (nx8604), .A1 (
          RST), .A2 (nx7664), .B0 (nx1710), .B1 (nx1790)) ;
    oai32 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix433 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .A0 (nx8604), .A1 (
          RST), .A2 (nx7664), .B0 (nx1714), .B1 (nx1790)) ;
    oai32 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix443 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .A0 (nx8606), .A1 (
          RST), .A2 (nx7664), .B0 (nx1718), .B1 (nx1790)) ;
    oai32 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix453 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .A0 (nx8606), .A1 (
          RST), .A2 (nx7666), .B0 (nx1722), .B1 (nx1790)) ;
    oai32 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix463 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .A0 (nx8606), .A1 (
          RST), .A2 (nx7666), .B0 (nx1726), .B1 (nx1792)) ;
    oai32 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix473 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .A0 (nx8606), .A1 (
          RST), .A2 (nx7666), .B0 (nx1730), .B1 (nx1792)) ;
    oai32 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix483 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .A0 (nx1772), .A1 (
          RST), .A2 (nx7666), .B0 (nx1734), .B1 (nx1792)) ;
    oai32 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix493 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .A0 (nx1794), .A1 (
          RST), .A2 (nx7666), .B0 (nx1738), .B1 (nx1792)) ;
    inv01 ix1793 (.Y (nx1794), .A (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_10)) ;
    oai32 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix503 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .A0 (nx1796), .A1 (
          RST), .A2 (nx7666), .B0 (nx1742), .B1 (nx1792)) ;
    inv01 ix1795 (.Y (nx1796), .A (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_11)) ;
    oai32 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix513 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .A0 (nx1798), .A1 (
          RST), .A2 (nx7666), .B0 (nx1746), .B1 (nx1792)) ;
    inv01 ix1797 (.Y (nx1798), .A (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_12)) ;
    oai32 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix523 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .A0 (nx1800), .A1 (
          RST), .A2 (nx7668), .B0 (nx1750), .B1 (nx1792)) ;
    inv01 ix1799 (.Y (nx1800), .A (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_13)) ;
    oai32 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix533 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .A0 (nx1802), .A1 (
          RST), .A2 (nx7668), .B0 (nx1754), .B1 (nx1804)) ;
    inv01 ix1801 (.Y (nx1802), .A (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_14)) ;
    inv01 ix1803 (.Y (nx1804), .A (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566)) ;
    oai32 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix543 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .A0 (nx1806), .A1 (
          RST), .A2 (nx7668), .B0 (nx1758), .B1 (nx1804)) ;
    inv01 ix1805 (.Y (nx1806), .A (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_15)) ;
    oai32 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix553 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .A0 (nx1808), .A1 (
          RST), .A2 (nx7668), .B0 (nx1762), .B1 (nx1804)) ;
    inv01 ix1807 (.Y (nx1808), .A (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_16)) ;
    nand02_2x L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix633 (.Y (nx1790), .A0 (
              nx7578), .A1 (nx7668)) ;
    nand02_2x L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix635 (.Y (nx1792), .A0 (
              nx7578), .A1 (nx7668)) ;
    oai32 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix393 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .A0 (nx1810), .A1 (
          RST), .A2 (nx7670), .B0 (L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx384), .B1 (
          nx1812)) ;
    inv01 ix1809 (.Y (nx1810), .A (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_0)) ;
    oai32 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix403 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .A0 (nx1814), .A1 (
          RST), .A2 (nx7670), .B0 (nx1630), .B1 (nx1812)) ;
    inv01 ix1813 (.Y (nx1814), .A (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_1)) ;
    oai32 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix413 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .A0 (nx1816), .A1 (
          RST), .A2 (nx7670), .B0 (L1_0_L2_1_G1_MINI_ALU_nx387), .B1 (nx1812)) ;
    inv01 ix1815 (.Y (nx1816), .A (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_2)) ;
    oai32 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix423 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .A0 (nx1818), .A1 (
          RST), .A2 (nx7670), .B0 (L1_0_L2_1_G1_MINI_ALU_nx399), .B1 (nx1812)) ;
    inv01 ix1817 (.Y (nx1818), .A (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_3)) ;
    oai32 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix433 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .A0 (nx1820), .A1 (
          RST), .A2 (nx7670), .B0 (L1_0_L2_1_G1_MINI_ALU_nx409), .B1 (nx1812)) ;
    inv01 ix1819 (.Y (nx1820), .A (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_4)) ;
    oai32 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix443 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .A0 (nx1822), .A1 (
          RST), .A2 (nx7670), .B0 (L1_0_L2_1_G1_MINI_ALU_nx419), .B1 (nx1812)) ;
    inv01 ix1821 (.Y (nx1822), .A (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_5)) ;
    oai32 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix453 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .A0 (nx1824), .A1 (
          RST), .A2 (nx7670), .B0 (L1_0_L2_1_G1_MINI_ALU_nx429), .B1 (nx1812)) ;
    inv01 ix1823 (.Y (nx1824), .A (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_6)) ;
    oai32 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix463 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .A0 (nx1826), .A1 (
          RST), .A2 (nx7672), .B0 (L1_0_L2_1_G1_MINI_ALU_nx439), .B1 (nx1828)) ;
    inv01 ix1825 (.Y (nx1826), .A (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_7)) ;
    oai32 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix473 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .A0 (nx1830), .A1 (
          RST), .A2 (nx7672), .B0 (L1_0_L2_1_G1_MINI_ALU_nx449), .B1 (nx1828)) ;
    inv01 ix1829 (.Y (nx1830), .A (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_8)) ;
    oai32 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix483 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .A0 (nx1832), .A1 (
          RST), .A2 (nx7672), .B0 (L1_0_L2_1_G1_MINI_ALU_nx469), .B1 (nx1828)) ;
    inv01 ix1831 (.Y (nx1832), .A (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_9)) ;
    oai32 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix493 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .A0 (nx1834), .A1 (
          RST), .A2 (nx7672), .B0 (L1_0_L2_1_G1_MINI_ALU_nx477), .B1 (nx1828)) ;
    inv01 ix1833 (.Y (nx1834), .A (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_10)) ;
    oai32 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix503 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .A0 (nx1836), .A1 (
          RST), .A2 (nx7672), .B0 (L1_0_L2_1_G1_MINI_ALU_nx485), .B1 (nx1828)) ;
    inv01 ix1835 (.Y (nx1836), .A (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_11)) ;
    oai32 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix513 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .A0 (nx1838), .A1 (
          RST), .A2 (nx7672), .B0 (L1_0_L2_1_G1_MINI_ALU_nx493), .B1 (nx1828)) ;
    inv01 ix1837 (.Y (nx1838), .A (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_12)) ;
    oai32 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix523 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .A0 (nx1840), .A1 (
          RST), .A2 (nx7672), .B0 (L1_0_L2_1_G1_MINI_ALU_nx501), .B1 (nx1828)) ;
    inv01 ix1839 (.Y (nx1840), .A (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_13)) ;
    oai32 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix533 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .A0 (nx1842), .A1 (
          RST), .A2 (nx7674), .B0 (L1_0_L2_1_G1_MINI_ALU_nx509), .B1 (nx1844)) ;
    inv01 ix1841 (.Y (nx1842), .A (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_14)) ;
    inv01 ix1843 (.Y (nx1844), .A (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566)) ;
    oai32 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix543 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .A0 (nx1846), .A1 (
          RST), .A2 (nx7674), .B0 (L1_0_L2_1_G1_MINI_ALU_nx517), .B1 (nx1844)) ;
    inv01 ix1845 (.Y (nx1846), .A (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_15)) ;
    oai32 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix553 (.Y (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .A0 (nx1848), .A1 (
          RST), .A2 (nx7674), .B0 (nx1646), .B1 (nx1844)) ;
    inv01 ix1847 (.Y (nx1848), .A (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_16)) ;
    nand02_2x L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix633 (.Y (nx1812), .A0 (
              nx7578), .A1 (nx7674)) ;
    nand02_2x L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix635 (.Y (nx1828), .A0 (
              nx7578), .A1 (nx7674)) ;
    mux21 L1_0_L2_2_G1_MINI_ALU_ix404 (.Y (L1_0_L2_2_G1_MINI_ALU_nx403), .A0 (
          nx1850), .A1 (L1_0_L2_2_G1_MINI_ALU_BoothP_2), .S0 (
          L1_0_L2_2_G1_MINI_ALU_nx395)) ;
    inv01 ix1849 (.Y (nx1850), .A (L1_0_L2_2_G1_MINI_ALU_nx391)) ;
    mux21 L1_0_L2_2_G1_MINI_ALU_ix414 (.Y (L1_0_L2_2_G1_MINI_ALU_nx413), .A0 (
          nx1852), .A1 (L1_0_L2_2_G1_MINI_ALU_BoothP_3), .S0 (
          L1_0_L2_2_G1_MINI_ALU_nx405)) ;
    inv01 ix1851 (.Y (nx1852), .A (L1_0_L2_2_G1_MINI_ALU_nx403)) ;
    mux21 L1_0_L2_2_G1_MINI_ALU_ix424 (.Y (L1_0_L2_2_G1_MINI_ALU_nx423), .A0 (
          nx1854), .A1 (L1_0_L2_2_G1_MINI_ALU_BoothP_4), .S0 (
          L1_0_L2_2_G1_MINI_ALU_nx415)) ;
    inv01 ix1853 (.Y (nx1854), .A (L1_0_L2_2_G1_MINI_ALU_nx413)) ;
    mux21 L1_0_L2_2_G1_MINI_ALU_ix434 (.Y (L1_0_L2_2_G1_MINI_ALU_nx433), .A0 (
          nx1856), .A1 (L1_0_L2_2_G1_MINI_ALU_BoothP_5), .S0 (
          L1_0_L2_2_G1_MINI_ALU_nx425)) ;
    inv01 ix1855 (.Y (nx1856), .A (L1_0_L2_2_G1_MINI_ALU_nx423)) ;
    mux21 L1_0_L2_2_G1_MINI_ALU_ix444 (.Y (L1_0_L2_2_G1_MINI_ALU_nx443), .A0 (
          nx1858), .A1 (L1_0_L2_2_G1_MINI_ALU_BoothP_6), .S0 (
          L1_0_L2_2_G1_MINI_ALU_nx435)) ;
    inv01 ix1857 (.Y (nx1858), .A (L1_0_L2_2_G1_MINI_ALU_nx433)) ;
    mux21 L1_0_L2_2_G1_MINI_ALU_ix454 (.Y (L1_0_L2_2_G1_MINI_ALU_nx453), .A0 (
          nx1860), .A1 (L1_0_L2_2_G1_MINI_ALU_BoothP_7), .S0 (
          L1_0_L2_2_G1_MINI_ALU_nx445)) ;
    inv01 ix1859 (.Y (nx1860), .A (L1_0_L2_2_G1_MINI_ALU_nx443)) ;
    mux21 L1_0_L2_2_G1_MINI_ALU_ix462 (.Y (L1_0_L2_2_G1_MINI_ALU_nx461), .A0 (
          nx1862), .A1 (L1_0_L2_2_G1_MINI_ALU_BoothP_8), .S0 (
          L1_0_L2_2_G1_MINI_ALU_nx455)) ;
    inv01 ix1861 (.Y (nx1862), .A (L1_0_L2_2_G1_MINI_ALU_nx453)) ;
    mux21 L1_0_L2_2_G1_MINI_ALU_ix468 (.Y (L1_0_L2_2_G1_MINI_ALU_nx467), .A0 (
          nx1864), .A1 (L1_0_L2_2_G1_MINI_ALU_BoothP_9), .S0 (
          L1_0_L2_2_G1_MINI_ALU_nx463)) ;
    inv01 ix1863 (.Y (nx1864), .A (L1_0_L2_2_G1_MINI_ALU_nx461)) ;
    mux21 L1_0_L2_2_G1_MINI_ALU_ix476 (.Y (L1_0_L2_2_G1_MINI_ALU_nx475), .A0 (
          nx1866), .A1 (L1_0_L2_2_G1_MINI_ALU_BoothP_10), .S0 (
          L1_0_L2_2_G1_MINI_ALU_nx471)) ;
    inv01 ix1865 (.Y (nx1866), .A (L1_0_L2_2_G1_MINI_ALU_nx467)) ;
    mux21 L1_0_L2_2_G1_MINI_ALU_ix484 (.Y (L1_0_L2_2_G1_MINI_ALU_nx483), .A0 (
          nx1868), .A1 (L1_0_L2_2_G1_MINI_ALU_BoothP_11), .S0 (
          L1_0_L2_2_G1_MINI_ALU_nx479)) ;
    inv01 ix1867 (.Y (nx1868), .A (L1_0_L2_2_G1_MINI_ALU_nx475)) ;
    mux21 L1_0_L2_2_G1_MINI_ALU_ix492 (.Y (L1_0_L2_2_G1_MINI_ALU_nx491), .A0 (
          nx1870), .A1 (L1_0_L2_2_G1_MINI_ALU_BoothP_12), .S0 (
          L1_0_L2_2_G1_MINI_ALU_nx487)) ;
    inv01 ix1869 (.Y (nx1870), .A (L1_0_L2_2_G1_MINI_ALU_nx483)) ;
    mux21 L1_0_L2_2_G1_MINI_ALU_ix500 (.Y (L1_0_L2_2_G1_MINI_ALU_nx499), .A0 (
          nx1872), .A1 (L1_0_L2_2_G1_MINI_ALU_BoothP_13), .S0 (
          L1_0_L2_2_G1_MINI_ALU_nx495)) ;
    inv01 ix1871 (.Y (nx1872), .A (L1_0_L2_2_G1_MINI_ALU_nx491)) ;
    mux21 L1_0_L2_2_G1_MINI_ALU_ix508 (.Y (L1_0_L2_2_G1_MINI_ALU_nx507), .A0 (
          nx1874), .A1 (L1_0_L2_2_G1_MINI_ALU_BoothP_14), .S0 (
          L1_0_L2_2_G1_MINI_ALU_nx503)) ;
    inv01 ix1873 (.Y (nx1874), .A (L1_0_L2_2_G1_MINI_ALU_nx499)) ;
    mux21 L1_0_L2_2_G1_MINI_ALU_ix516 (.Y (L1_0_L2_2_G1_MINI_ALU_nx515), .A0 (
          nx1876), .A1 (L1_0_L2_2_G1_MINI_ALU_BoothP_15), .S0 (
          L1_0_L2_2_G1_MINI_ALU_nx511)) ;
    inv01 ix1875 (.Y (nx1876), .A (L1_0_L2_2_G1_MINI_ALU_nx507)) ;
    mux21 L1_0_L2_2_G1_MINI_ALU_ix161 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_1), .A0 (nx1878), .A1 (
          L1_0_L2_2_G1_MINI_ALU_nx379), .S0 (nx7678)) ;
    inv01 ix1877 (.Y (nx1878), .A (L1_0_L2_2_G1_MINI_ALU_BoothP_1)) ;
    mux21 L1_0_L2_2_G1_MINI_ALU_ix181 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_2), .A0 (
          L1_0_L2_2_G1_MINI_ALU_nx387), .A1 (L1_0_L2_2_G1_MINI_ALU_nx389), .S0 (
          nx7678)) ;
    mux21 L1_0_L2_2_G1_MINI_ALU_ix201 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_3), .A0 (
          L1_0_L2_2_G1_MINI_ALU_nx399), .A1 (L1_0_L2_2_G1_MINI_ALU_nx401), .S0 (
          nx7678)) ;
    mux21 L1_0_L2_2_G1_MINI_ALU_ix221 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_4), .A0 (
          L1_0_L2_2_G1_MINI_ALU_nx409), .A1 (L1_0_L2_2_G1_MINI_ALU_nx411), .S0 (
          nx7678)) ;
    mux21 L1_0_L2_2_G1_MINI_ALU_ix241 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_5), .A0 (
          L1_0_L2_2_G1_MINI_ALU_nx419), .A1 (L1_0_L2_2_G1_MINI_ALU_nx421), .S0 (
          nx7678)) ;
    mux21 L1_0_L2_2_G1_MINI_ALU_ix261 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_6), .A0 (
          L1_0_L2_2_G1_MINI_ALU_nx429), .A1 (L1_0_L2_2_G1_MINI_ALU_nx431), .S0 (
          nx7678)) ;
    mux21 L1_0_L2_2_G1_MINI_ALU_ix281 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_7), .A0 (
          L1_0_L2_2_G1_MINI_ALU_nx439), .A1 (L1_0_L2_2_G1_MINI_ALU_nx441), .S0 (
          nx7678)) ;
    mux21 L1_0_L2_2_G1_MINI_ALU_ix301 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_8), .A0 (
          L1_0_L2_2_G1_MINI_ALU_nx449), .A1 (L1_0_L2_2_G1_MINI_ALU_nx451), .S0 (
          nx7680)) ;
    mux21 L1_0_L2_2_G1_MINI_ALU_ix321 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_9), .A0 (
          L1_0_L2_2_G1_MINI_ALU_nx469), .A1 (nx1880), .S0 (nx7680)) ;
    inv01 ix1879 (.Y (nx1880), .A (L1_0_L2_2_G1_MINI_ALU_nx316)) ;
    mux21 L1_0_L2_2_G1_MINI_ALU_ix341 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_10), .A0 (
          L1_0_L2_2_G1_MINI_ALU_nx477), .A1 (nx1882), .S0 (nx7680)) ;
    inv01 ix1881 (.Y (nx1882), .A (L1_0_L2_2_G1_MINI_ALU_nx336)) ;
    mux21 L1_0_L2_2_G1_MINI_ALU_ix361 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_11), .A0 (
          L1_0_L2_2_G1_MINI_ALU_nx485), .A1 (nx1884), .S0 (nx7680)) ;
    inv01 ix1883 (.Y (nx1884), .A (L1_0_L2_2_G1_MINI_ALU_nx356)) ;
    mux21 L1_0_L2_2_G1_MINI_ALU_ix381 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_12), .A0 (
          L1_0_L2_2_G1_MINI_ALU_nx493), .A1 (nx1886), .S0 (nx7680)) ;
    inv01 ix1885 (.Y (nx1886), .A (L1_0_L2_2_G1_MINI_ALU_nx376)) ;
    mux21 L1_0_L2_2_G1_MINI_ALU_ix401 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_13), .A0 (
          L1_0_L2_2_G1_MINI_ALU_nx501), .A1 (nx1888), .S0 (nx7680)) ;
    inv01 ix1887 (.Y (nx1888), .A (L1_0_L2_2_G1_MINI_ALU_nx396)) ;
    mux21 L1_0_L2_2_G1_MINI_ALU_ix421 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_14), .A0 (
          L1_0_L2_2_G1_MINI_ALU_nx509), .A1 (nx1890), .S0 (nx7680)) ;
    inv01 ix1889 (.Y (nx1890), .A (L1_0_L2_2_G1_MINI_ALU_nx416)) ;
    mux21 L1_0_L2_2_G1_MINI_ALU_ix441 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_15), .A0 (
          L1_0_L2_2_G1_MINI_ALU_nx517), .A1 (nx1892), .S0 (nx7682)) ;
    inv01 ix1891 (.Y (nx1892), .A (L1_0_L2_2_G1_MINI_ALU_nx436)) ;
    mux21 L1_0_L2_2_G1_MINI_ALU_ix461 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_16), .A0 (nx1894), .A1 (nx1896
          ), .S0 (nx7682)) ;
    inv01 ix1893 (.Y (nx1894), .A (L1_0_L2_2_G1_MINI_ALU_BoothP_16)) ;
    inv01 ix1895 (.Y (nx1896), .A (L1_0_L2_2_G1_MINI_ALU_nx456)) ;
    nor02_2x L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix319 (.Y (
             L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642), .A0 (Start), .A1 (
             CalculatingBooth_dup_1084)) ;
    nor02_2x L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix85 (.Y (
             L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_0), .A0 (nx7692), .A1 (
             nx1898)) ;
    inv01 ix1897 (.Y (nx1898), .A (L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_1)) ;
    mux21 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix125 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_1), .A0 (nx1900), .A1 (
          nx1902), .S0 (nx7692)) ;
    inv01 ix1899 (.Y (nx1900), .A (L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_2)) ;
    inv01 ix1901 (.Y (nx1902), .A (WindowDin_0__2__0)) ;
    mux21 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix133 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_2), .A0 (nx1904), .A1 (
          nx1906), .S0 (nx7692)) ;
    inv01 ix1903 (.Y (nx1904), .A (L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_3)) ;
    inv01 ix1905 (.Y (nx1906), .A (WindowDin_0__2__1)) ;
    mux21 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix141 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_3), .A0 (nx1908), .A1 (
          nx1910), .S0 (nx7692)) ;
    inv01 ix1907 (.Y (nx1908), .A (L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_4)) ;
    inv01 ix1909 (.Y (nx1910), .A (WindowDin_0__2__2)) ;
    mux21 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix149 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_4), .A0 (nx1912), .A1 (
          nx1914), .S0 (nx7692)) ;
    inv01 ix1911 (.Y (nx1912), .A (L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_5)) ;
    inv01 ix1913 (.Y (nx1914), .A (WindowDin_0__2__3)) ;
    mux21 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix157 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_5), .A0 (nx1916), .A1 (
          nx1918), .S0 (nx7692)) ;
    inv01 ix1915 (.Y (nx1916), .A (L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_6)) ;
    inv01 ix1917 (.Y (nx1918), .A (WindowDin_0__2__4)) ;
    mux21 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix165 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_6), .A0 (nx1920), .A1 (
          nx1922), .S0 (nx7692)) ;
    inv01 ix1919 (.Y (nx1920), .A (L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_7)) ;
    inv01 ix1921 (.Y (nx1922), .A (WindowDin_0__2__5)) ;
    mux21 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix173 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_7), .A0 (nx1924), .A1 (
          nx1926), .S0 (nx7694)) ;
    inv01 ix1923 (.Y (nx1924), .A (L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_8)) ;
    inv01 ix1925 (.Y (nx1926), .A (WindowDin_0__2__6)) ;
    mux21 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix181 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_8), .A0 (nx1928), .A1 (
          nx1930), .S0 (nx7694)) ;
    inv01 ix1927 (.Y (nx1928), .A (L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_9)) ;
    inv01 ix1929 (.Y (nx1930), .A (WindowDin_0__2__7)) ;
    nor02_2x L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix89 (.Y (
             L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_9), .A0 (nx7694), .A1 (
             nx1932)) ;
    inv01 ix1931 (.Y (nx1932), .A (L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_10)
          ) ;
    nor02_2x L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix93 (.Y (
             L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_10), .A0 (nx7694), .A1 (
             nx1934)) ;
    inv01 ix1933 (.Y (nx1934), .A (L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_11)
          ) ;
    nor02_2x L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix97 (.Y (
             L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_11), .A0 (nx7694), .A1 (
             nx1936)) ;
    inv01 ix1935 (.Y (nx1936), .A (L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_12)
          ) ;
    nor02_2x L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix101 (.Y (
             L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_12), .A0 (nx7694), .A1 (
             nx1938)) ;
    inv01 ix1937 (.Y (nx1938), .A (L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_13)
          ) ;
    nor02_2x L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix105 (.Y (
             L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_13), .A0 (nx7694), .A1 (
             nx1940)) ;
    inv01 ix1939 (.Y (nx1940), .A (L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_14)
          ) ;
    nor02_2x L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix109 (.Y (
             L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_14), .A0 (nx7696), .A1 (
             nx1942)) ;
    inv01 ix1941 (.Y (nx1942), .A (L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_15)
          ) ;
    nor02_2x L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix113 (.Y (
             L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_15), .A0 (nx7696), .A1 (
             nx1944)) ;
    inv01 ix1943 (.Y (nx1944), .A (L1_0_L2_2_G1_MINI_ALU_BoothPBeforeShift_16)
          ) ;
    nor02_2x L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix117 (.Y (
             L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_16), .A0 (nx7696), .A1 (
             nx1944)) ;
    mux21 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix189 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BoothOperand_0), .A0 (nx1946), .A1 (nx1948), .S0 (
          nx7684)) ;
    inv01 ix1945 (.Y (nx1946), .A (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_0)) ;
    inv01 ix1947 (.Y (nx1948), .A (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_0)) ;
    mux21 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix197 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BoothOperand_1), .A0 (nx1950), .A1 (nx1952), .S0 (
          nx7684)) ;
    inv01 ix1949 (.Y (nx1950), .A (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_1)) ;
    inv01 ix1951 (.Y (nx1952), .A (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_1)) ;
    mux21 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix205 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BoothOperand_2), .A0 (nx1954), .A1 (nx1956), .S0 (
          nx7684)) ;
    inv01 ix1953 (.Y (nx1954), .A (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_2)) ;
    inv01 ix1955 (.Y (nx1956), .A (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_2)) ;
    mux21 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix213 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BoothOperand_3), .A0 (nx1958), .A1 (nx1960), .S0 (
          nx7684)) ;
    inv01 ix1957 (.Y (nx1958), .A (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_3)) ;
    inv01 ix1959 (.Y (nx1960), .A (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_3)) ;
    mux21 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix221 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BoothOperand_4), .A0 (nx1962), .A1 (nx1964), .S0 (
          nx7684)) ;
    inv01 ix1961 (.Y (nx1962), .A (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_4)) ;
    inv01 ix1963 (.Y (nx1964), .A (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_4)) ;
    mux21 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix229 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BoothOperand_5), .A0 (nx1966), .A1 (nx1968), .S0 (
          nx7686)) ;
    inv01 ix1965 (.Y (nx1966), .A (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_5)) ;
    inv01 ix1967 (.Y (nx1968), .A (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_5)) ;
    mux21 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix237 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BoothOperand_6), .A0 (nx1970), .A1 (nx1972), .S0 (
          nx7686)) ;
    inv01 ix1969 (.Y (nx1970), .A (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_6)) ;
    inv01 ix1971 (.Y (nx1972), .A (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_6)) ;
    mux21 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix245 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BoothOperand_7), .A0 (nx1974), .A1 (nx1976), .S0 (
          nx7686)) ;
    inv01 ix1973 (.Y (nx1974), .A (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_7)) ;
    inv01 ix1975 (.Y (nx1976), .A (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_7)) ;
    mux21 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix253 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BoothOperand_8), .A0 (nx1978), .A1 (nx1980), .S0 (
          nx7686)) ;
    inv01 ix1977 (.Y (nx1978), .A (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_8)) ;
    inv01 ix1979 (.Y (nx1980), .A (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_8)) ;
    mux21 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix261 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BoothOperand_9), .A0 (nx1982), .A1 (nx1984), .S0 (
          nx7686)) ;
    inv01 ix1981 (.Y (nx1982), .A (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_9)) ;
    inv01 ix1983 (.Y (nx1984), .A (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_9)) ;
    mux21 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix269 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BoothOperand_10), .A0 (nx1986), .A1 (nx1988), .S0 (
          nx7686)) ;
    inv01 ix1985 (.Y (nx1986), .A (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_10)) ;
    inv01 ix1987 (.Y (nx1988), .A (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_10)) ;
    mux21 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix277 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BoothOperand_11), .A0 (nx1990), .A1 (nx1992), .S0 (
          nx7686)) ;
    inv01 ix1989 (.Y (nx1990), .A (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_11)) ;
    inv01 ix1991 (.Y (nx1992), .A (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_11)) ;
    mux21 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix285 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BoothOperand_12), .A0 (nx1994), .A1 (nx1996), .S0 (
          nx7688)) ;
    inv01 ix1993 (.Y (nx1994), .A (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_12)) ;
    inv01 ix1995 (.Y (nx1996), .A (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_12)) ;
    mux21 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix293 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BoothOperand_13), .A0 (nx1998), .A1 (nx2000), .S0 (
          nx7688)) ;
    inv01 ix1997 (.Y (nx1998), .A (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_13)) ;
    inv01 ix1999 (.Y (nx2000), .A (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_13)) ;
    mux21 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix301 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BoothOperand_14), .A0 (nx2002), .A1 (nx2004), .S0 (
          nx7688)) ;
    inv01 ix2001 (.Y (nx2002), .A (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_14)) ;
    inv01 ix2003 (.Y (nx2004), .A (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_14)) ;
    mux21 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix309 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BoothOperand_15), .A0 (nx2006), .A1 (nx2008), .S0 (
          nx7688)) ;
    inv01 ix2005 (.Y (nx2006), .A (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_15)) ;
    inv01 ix2007 (.Y (nx2008), .A (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_15)) ;
    mux21 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix317 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BoothOperand_16), .A0 (nx2010), .A1 (nx2012), .S0 (
          nx7688)) ;
    inv01 ix2009 (.Y (nx2010), .A (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_16)) ;
    inv01 ix2011 (.Y (nx2012), .A (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_16)) ;
    xnor2 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix321 (.Y (
          L1_0_L2_2_G1_MINI_ALU_AddPToBoothOperand), .A0 (nx7688), .A1 (nx1878)
          ) ;
    oai32 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix393 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .A0 (nx8608), .A1 (
          RST), .A2 (nx7698), .B0 (nx1948), .B1 (nx2016)) ;
    oai32 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix403 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .A0 (nx8608), .A1 (
          RST), .A2 (nx7698), .B0 (nx1952), .B1 (nx2016)) ;
    oai32 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix413 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .A0 (nx8608), .A1 (
          RST), .A2 (nx7698), .B0 (nx1956), .B1 (nx2016)) ;
    oai32 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix423 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .A0 (nx8608), .A1 (
          RST), .A2 (nx7698), .B0 (nx1960), .B1 (nx2016)) ;
    oai32 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix433 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .A0 (nx8608), .A1 (
          RST), .A2 (nx7698), .B0 (nx1964), .B1 (nx2016)) ;
    oai32 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix443 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .A0 (nx8608), .A1 (
          RST), .A2 (nx7698), .B0 (nx1968), .B1 (nx2016)) ;
    oai32 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix453 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .A0 (nx8608), .A1 (
          RST), .A2 (nx7700), .B0 (nx1972), .B1 (nx2016)) ;
    oai32 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix463 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .A0 (nx8610), .A1 (
          RST), .A2 (nx7700), .B0 (nx1976), .B1 (nx2018)) ;
    oai32 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix473 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .A0 (nx8610), .A1 (
          RST), .A2 (nx7700), .B0 (nx1980), .B1 (nx2018)) ;
    oai32 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix483 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .A0 (nx2020), .A1 (
          RST), .A2 (nx7700), .B0 (nx1984), .B1 (nx2018)) ;
    inv01 ix2019 (.Y (nx2020), .A (FilterDin_0__2__0)) ;
    oai32 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix493 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .A0 (nx2022), .A1 (
          RST), .A2 (nx7700), .B0 (nx1988), .B1 (nx2018)) ;
    inv01 ix2021 (.Y (nx2022), .A (FilterDin_0__2__1)) ;
    oai32 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix503 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .A0 (nx2024), .A1 (
          RST), .A2 (nx7700), .B0 (nx1992), .B1 (nx2018)) ;
    inv01 ix2023 (.Y (nx2024), .A (FilterDin_0__2__2)) ;
    oai32 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix513 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .A0 (nx2026), .A1 (
          RST), .A2 (nx7700), .B0 (nx1996), .B1 (nx2018)) ;
    inv01 ix2025 (.Y (nx2026), .A (FilterDin_0__2__3)) ;
    oai32 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix523 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .A0 (nx2028), .A1 (
          RST), .A2 (nx7702), .B0 (nx2000), .B1 (nx2018)) ;
    inv01 ix2027 (.Y (nx2028), .A (FilterDin_0__2__4)) ;
    oai32 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix533 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .A0 (nx2030), .A1 (
          RST), .A2 (nx7702), .B0 (nx2004), .B1 (nx2032)) ;
    inv01 ix2029 (.Y (nx2030), .A (FilterDin_0__2__5)) ;
    inv01 ix2031 (.Y (nx2032), .A (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566)) ;
    oai32 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix543 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .A0 (nx2034), .A1 (
          RST), .A2 (nx7702), .B0 (nx2008), .B1 (nx2032)) ;
    inv01 ix2033 (.Y (nx2034), .A (FilterDin_0__2__6)) ;
    oai32 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix553 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .A0 (nx2036), .A1 (
          RST), .A2 (nx7702), .B0 (nx2012), .B1 (nx2032)) ;
    inv01 ix2035 (.Y (nx2036), .A (FilterDin_0__2__7)) ;
    nand02_2x L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix633 (.Y (nx2016), .A0 (
              nx7578), .A1 (nx7702)) ;
    nand02_2x L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix635 (.Y (nx2018), .A0 (
              nx7578), .A1 (nx7702)) ;
    oai32 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix393 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .A0 (nx8610), .A1 (
          RST), .A2 (nx7704), .B0 (nx1946), .B1 (nx2038)) ;
    oai32 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix403 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .A0 (nx8610), .A1 (
          RST), .A2 (nx7704), .B0 (nx1950), .B1 (nx2038)) ;
    oai32 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix413 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .A0 (nx8610), .A1 (
          RST), .A2 (nx7704), .B0 (nx1954), .B1 (nx2038)) ;
    oai32 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix423 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .A0 (nx8610), .A1 (
          RST), .A2 (nx7704), .B0 (nx1958), .B1 (nx2038)) ;
    oai32 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix433 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .A0 (nx8610), .A1 (
          RST), .A2 (nx7704), .B0 (nx1962), .B1 (nx2038)) ;
    oai32 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix443 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .A0 (nx8612), .A1 (
          RST), .A2 (nx7704), .B0 (nx1966), .B1 (nx2038)) ;
    oai32 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix453 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .A0 (nx8612), .A1 (
          RST), .A2 (nx7706), .B0 (nx1970), .B1 (nx2038)) ;
    oai32 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix463 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .A0 (nx8612), .A1 (
          RST), .A2 (nx7706), .B0 (nx1974), .B1 (nx2040)) ;
    oai32 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix473 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .A0 (nx8612), .A1 (
          RST), .A2 (nx7706), .B0 (nx1978), .B1 (nx2040)) ;
    oai32 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix483 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .A0 (nx2020), .A1 (
          RST), .A2 (nx7706), .B0 (nx1982), .B1 (nx2040)) ;
    oai32 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix493 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .A0 (nx2042), .A1 (
          RST), .A2 (nx7706), .B0 (nx1986), .B1 (nx2040)) ;
    inv01 ix2041 (.Y (nx2042), .A (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_10)) ;
    oai32 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix503 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .A0 (nx2044), .A1 (
          RST), .A2 (nx7706), .B0 (nx1990), .B1 (nx2040)) ;
    inv01 ix2043 (.Y (nx2044), .A (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_11)) ;
    oai32 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix513 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .A0 (nx2046), .A1 (
          RST), .A2 (nx7706), .B0 (nx1994), .B1 (nx2040)) ;
    inv01 ix2045 (.Y (nx2046), .A (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_12)) ;
    oai32 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix523 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .A0 (nx2048), .A1 (
          RST), .A2 (nx7708), .B0 (nx1998), .B1 (nx2040)) ;
    inv01 ix2047 (.Y (nx2048), .A (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_13)) ;
    oai32 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix533 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .A0 (nx2050), .A1 (
          RST), .A2 (nx7708), .B0 (nx2002), .B1 (nx2052)) ;
    inv01 ix2049 (.Y (nx2050), .A (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_14)) ;
    inv01 ix2051 (.Y (nx2052), .A (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566)) ;
    oai32 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix543 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .A0 (nx2054), .A1 (
          RST), .A2 (nx7708), .B0 (nx2006), .B1 (nx2052)) ;
    inv01 ix2053 (.Y (nx2054), .A (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_15)) ;
    oai32 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix553 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .A0 (nx2056), .A1 (
          RST), .A2 (nx7708), .B0 (nx2010), .B1 (nx2052)) ;
    inv01 ix2055 (.Y (nx2056), .A (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_16)) ;
    nand02_2x L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix633 (.Y (nx2038), .A0 (
              nx7580), .A1 (nx7708)) ;
    nand02_2x L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix635 (.Y (nx2040), .A0 (
              nx7580), .A1 (nx7708)) ;
    oai32 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix393 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .A0 (nx2058), .A1 (
          RST), .A2 (nx7710), .B0 (L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx384), .B1 (
          nx2060)) ;
    inv01 ix2057 (.Y (nx2058), .A (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_0)) ;
    oai32 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix403 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .A0 (nx2062), .A1 (
          RST), .A2 (nx7710), .B0 (nx1878), .B1 (nx2060)) ;
    inv01 ix2061 (.Y (nx2062), .A (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_1)) ;
    oai32 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix413 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .A0 (nx2064), .A1 (
          RST), .A2 (nx7710), .B0 (L1_0_L2_2_G1_MINI_ALU_nx387), .B1 (nx2060)) ;
    inv01 ix2063 (.Y (nx2064), .A (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_2)) ;
    oai32 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix423 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .A0 (nx2066), .A1 (
          RST), .A2 (nx7710), .B0 (L1_0_L2_2_G1_MINI_ALU_nx399), .B1 (nx2060)) ;
    inv01 ix2065 (.Y (nx2066), .A (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_3)) ;
    oai32 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix433 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .A0 (nx2068), .A1 (
          RST), .A2 (nx7710), .B0 (L1_0_L2_2_G1_MINI_ALU_nx409), .B1 (nx2060)) ;
    inv01 ix2067 (.Y (nx2068), .A (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_4)) ;
    oai32 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix443 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .A0 (nx2070), .A1 (
          RST), .A2 (nx7710), .B0 (L1_0_L2_2_G1_MINI_ALU_nx419), .B1 (nx2060)) ;
    inv01 ix2069 (.Y (nx2070), .A (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_5)) ;
    oai32 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix453 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .A0 (nx2072), .A1 (
          RST), .A2 (nx7710), .B0 (L1_0_L2_2_G1_MINI_ALU_nx429), .B1 (nx2060)) ;
    inv01 ix2071 (.Y (nx2072), .A (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_6)) ;
    oai32 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix463 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .A0 (nx2074), .A1 (
          RST), .A2 (nx7712), .B0 (L1_0_L2_2_G1_MINI_ALU_nx439), .B1 (nx2076)) ;
    inv01 ix2073 (.Y (nx2074), .A (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_7)) ;
    oai32 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix473 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .A0 (nx2078), .A1 (
          RST), .A2 (nx7712), .B0 (L1_0_L2_2_G1_MINI_ALU_nx449), .B1 (nx2076)) ;
    inv01 ix2077 (.Y (nx2078), .A (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_8)) ;
    oai32 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix483 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .A0 (nx2080), .A1 (
          RST), .A2 (nx7712), .B0 (L1_0_L2_2_G1_MINI_ALU_nx469), .B1 (nx2076)) ;
    inv01 ix2079 (.Y (nx2080), .A (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_9)) ;
    oai32 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix493 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .A0 (nx2082), .A1 (
          RST), .A2 (nx7712), .B0 (L1_0_L2_2_G1_MINI_ALU_nx477), .B1 (nx2076)) ;
    inv01 ix2081 (.Y (nx2082), .A (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_10)) ;
    oai32 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix503 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .A0 (nx2084), .A1 (
          RST), .A2 (nx7712), .B0 (L1_0_L2_2_G1_MINI_ALU_nx485), .B1 (nx2076)) ;
    inv01 ix2083 (.Y (nx2084), .A (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_11)) ;
    oai32 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix513 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .A0 (nx2086), .A1 (
          RST), .A2 (nx7712), .B0 (L1_0_L2_2_G1_MINI_ALU_nx493), .B1 (nx2076)) ;
    inv01 ix2085 (.Y (nx2086), .A (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_12)) ;
    oai32 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix523 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .A0 (nx2088), .A1 (
          RST), .A2 (nx7712), .B0 (L1_0_L2_2_G1_MINI_ALU_nx501), .B1 (nx2076)) ;
    inv01 ix2087 (.Y (nx2088), .A (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_13)) ;
    oai32 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix533 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .A0 (nx2090), .A1 (
          RST), .A2 (nx7714), .B0 (L1_0_L2_2_G1_MINI_ALU_nx509), .B1 (nx2092)) ;
    inv01 ix2089 (.Y (nx2090), .A (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_14)) ;
    inv01 ix2091 (.Y (nx2092), .A (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566)) ;
    oai32 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix543 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .A0 (nx2094), .A1 (
          RST), .A2 (nx7714), .B0 (L1_0_L2_2_G1_MINI_ALU_nx517), .B1 (nx2092)) ;
    inv01 ix2093 (.Y (nx2094), .A (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_15)) ;
    oai32 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix553 (.Y (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .A0 (nx2096), .A1 (
          RST), .A2 (nx7714), .B0 (nx1894), .B1 (nx2092)) ;
    inv01 ix2095 (.Y (nx2096), .A (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_16)) ;
    nand02_2x L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix633 (.Y (nx2060), .A0 (
              nx7580), .A1 (nx7714)) ;
    nand02_2x L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix635 (.Y (nx2076), .A0 (
              nx7580), .A1 (nx7714)) ;
    mux21 L1_0_L2_3_G1_MINI_ALU_ix404 (.Y (L1_0_L2_3_G1_MINI_ALU_nx403), .A0 (
          nx2098), .A1 (L1_0_L2_3_G1_MINI_ALU_BoothP_2), .S0 (
          L1_0_L2_3_G1_MINI_ALU_nx395)) ;
    inv01 ix2097 (.Y (nx2098), .A (L1_0_L2_3_G1_MINI_ALU_nx391)) ;
    mux21 L1_0_L2_3_G1_MINI_ALU_ix414 (.Y (L1_0_L2_3_G1_MINI_ALU_nx413), .A0 (
          nx2100), .A1 (L1_0_L2_3_G1_MINI_ALU_BoothP_3), .S0 (
          L1_0_L2_3_G1_MINI_ALU_nx405)) ;
    inv01 ix2099 (.Y (nx2100), .A (L1_0_L2_3_G1_MINI_ALU_nx403)) ;
    mux21 L1_0_L2_3_G1_MINI_ALU_ix424 (.Y (L1_0_L2_3_G1_MINI_ALU_nx423), .A0 (
          nx2102), .A1 (L1_0_L2_3_G1_MINI_ALU_BoothP_4), .S0 (
          L1_0_L2_3_G1_MINI_ALU_nx415)) ;
    inv01 ix2101 (.Y (nx2102), .A (L1_0_L2_3_G1_MINI_ALU_nx413)) ;
    mux21 L1_0_L2_3_G1_MINI_ALU_ix434 (.Y (L1_0_L2_3_G1_MINI_ALU_nx433), .A0 (
          nx2104), .A1 (L1_0_L2_3_G1_MINI_ALU_BoothP_5), .S0 (
          L1_0_L2_3_G1_MINI_ALU_nx425)) ;
    inv01 ix2103 (.Y (nx2104), .A (L1_0_L2_3_G1_MINI_ALU_nx423)) ;
    mux21 L1_0_L2_3_G1_MINI_ALU_ix444 (.Y (L1_0_L2_3_G1_MINI_ALU_nx443), .A0 (
          nx2106), .A1 (L1_0_L2_3_G1_MINI_ALU_BoothP_6), .S0 (
          L1_0_L2_3_G1_MINI_ALU_nx435)) ;
    inv01 ix2105 (.Y (nx2106), .A (L1_0_L2_3_G1_MINI_ALU_nx433)) ;
    mux21 L1_0_L2_3_G1_MINI_ALU_ix454 (.Y (L1_0_L2_3_G1_MINI_ALU_nx453), .A0 (
          nx2108), .A1 (L1_0_L2_3_G1_MINI_ALU_BoothP_7), .S0 (
          L1_0_L2_3_G1_MINI_ALU_nx445)) ;
    inv01 ix2107 (.Y (nx2108), .A (L1_0_L2_3_G1_MINI_ALU_nx443)) ;
    mux21 L1_0_L2_3_G1_MINI_ALU_ix462 (.Y (L1_0_L2_3_G1_MINI_ALU_nx461), .A0 (
          nx2110), .A1 (L1_0_L2_3_G1_MINI_ALU_BoothP_8), .S0 (
          L1_0_L2_3_G1_MINI_ALU_nx455)) ;
    inv01 ix2109 (.Y (nx2110), .A (L1_0_L2_3_G1_MINI_ALU_nx453)) ;
    mux21 L1_0_L2_3_G1_MINI_ALU_ix468 (.Y (L1_0_L2_3_G1_MINI_ALU_nx467), .A0 (
          nx2112), .A1 (L1_0_L2_3_G1_MINI_ALU_BoothP_9), .S0 (
          L1_0_L2_3_G1_MINI_ALU_nx463)) ;
    inv01 ix2111 (.Y (nx2112), .A (L1_0_L2_3_G1_MINI_ALU_nx461)) ;
    mux21 L1_0_L2_3_G1_MINI_ALU_ix476 (.Y (L1_0_L2_3_G1_MINI_ALU_nx475), .A0 (
          nx2114), .A1 (L1_0_L2_3_G1_MINI_ALU_BoothP_10), .S0 (
          L1_0_L2_3_G1_MINI_ALU_nx471)) ;
    inv01 ix2113 (.Y (nx2114), .A (L1_0_L2_3_G1_MINI_ALU_nx467)) ;
    mux21 L1_0_L2_3_G1_MINI_ALU_ix484 (.Y (L1_0_L2_3_G1_MINI_ALU_nx483), .A0 (
          nx2116), .A1 (L1_0_L2_3_G1_MINI_ALU_BoothP_11), .S0 (
          L1_0_L2_3_G1_MINI_ALU_nx479)) ;
    inv01 ix2115 (.Y (nx2116), .A (L1_0_L2_3_G1_MINI_ALU_nx475)) ;
    mux21 L1_0_L2_3_G1_MINI_ALU_ix492 (.Y (L1_0_L2_3_G1_MINI_ALU_nx491), .A0 (
          nx2118), .A1 (L1_0_L2_3_G1_MINI_ALU_BoothP_12), .S0 (
          L1_0_L2_3_G1_MINI_ALU_nx487)) ;
    inv01 ix2117 (.Y (nx2118), .A (L1_0_L2_3_G1_MINI_ALU_nx483)) ;
    mux21 L1_0_L2_3_G1_MINI_ALU_ix500 (.Y (L1_0_L2_3_G1_MINI_ALU_nx499), .A0 (
          nx2120), .A1 (L1_0_L2_3_G1_MINI_ALU_BoothP_13), .S0 (
          L1_0_L2_3_G1_MINI_ALU_nx495)) ;
    inv01 ix2119 (.Y (nx2120), .A (L1_0_L2_3_G1_MINI_ALU_nx491)) ;
    mux21 L1_0_L2_3_G1_MINI_ALU_ix508 (.Y (L1_0_L2_3_G1_MINI_ALU_nx507), .A0 (
          nx2122), .A1 (L1_0_L2_3_G1_MINI_ALU_BoothP_14), .S0 (
          L1_0_L2_3_G1_MINI_ALU_nx503)) ;
    inv01 ix2121 (.Y (nx2122), .A (L1_0_L2_3_G1_MINI_ALU_nx499)) ;
    mux21 L1_0_L2_3_G1_MINI_ALU_ix516 (.Y (L1_0_L2_3_G1_MINI_ALU_nx515), .A0 (
          nx2124), .A1 (L1_0_L2_3_G1_MINI_ALU_BoothP_15), .S0 (
          L1_0_L2_3_G1_MINI_ALU_nx511)) ;
    inv01 ix2123 (.Y (nx2124), .A (L1_0_L2_3_G1_MINI_ALU_nx507)) ;
    mux21 L1_0_L2_3_G1_MINI_ALU_ix161 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_1), .A0 (nx2126), .A1 (
          L1_0_L2_3_G1_MINI_ALU_nx379), .S0 (nx7718)) ;
    inv01 ix2125 (.Y (nx2126), .A (L1_0_L2_3_G1_MINI_ALU_BoothP_1)) ;
    mux21 L1_0_L2_3_G1_MINI_ALU_ix181 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_2), .A0 (
          L1_0_L2_3_G1_MINI_ALU_nx387), .A1 (L1_0_L2_3_G1_MINI_ALU_nx389), .S0 (
          nx7718)) ;
    mux21 L1_0_L2_3_G1_MINI_ALU_ix201 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_3), .A0 (
          L1_0_L2_3_G1_MINI_ALU_nx399), .A1 (L1_0_L2_3_G1_MINI_ALU_nx401), .S0 (
          nx7718)) ;
    mux21 L1_0_L2_3_G1_MINI_ALU_ix221 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_4), .A0 (
          L1_0_L2_3_G1_MINI_ALU_nx409), .A1 (L1_0_L2_3_G1_MINI_ALU_nx411), .S0 (
          nx7718)) ;
    mux21 L1_0_L2_3_G1_MINI_ALU_ix241 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_5), .A0 (
          L1_0_L2_3_G1_MINI_ALU_nx419), .A1 (L1_0_L2_3_G1_MINI_ALU_nx421), .S0 (
          nx7718)) ;
    mux21 L1_0_L2_3_G1_MINI_ALU_ix261 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_6), .A0 (
          L1_0_L2_3_G1_MINI_ALU_nx429), .A1 (L1_0_L2_3_G1_MINI_ALU_nx431), .S0 (
          nx7718)) ;
    mux21 L1_0_L2_3_G1_MINI_ALU_ix281 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_7), .A0 (
          L1_0_L2_3_G1_MINI_ALU_nx439), .A1 (L1_0_L2_3_G1_MINI_ALU_nx441), .S0 (
          nx7718)) ;
    mux21 L1_0_L2_3_G1_MINI_ALU_ix301 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_8), .A0 (
          L1_0_L2_3_G1_MINI_ALU_nx449), .A1 (L1_0_L2_3_G1_MINI_ALU_nx451), .S0 (
          nx7720)) ;
    mux21 L1_0_L2_3_G1_MINI_ALU_ix321 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_9), .A0 (
          L1_0_L2_3_G1_MINI_ALU_nx469), .A1 (nx2128), .S0 (nx7720)) ;
    inv01 ix2127 (.Y (nx2128), .A (L1_0_L2_3_G1_MINI_ALU_nx316)) ;
    mux21 L1_0_L2_3_G1_MINI_ALU_ix341 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_10), .A0 (
          L1_0_L2_3_G1_MINI_ALU_nx477), .A1 (nx2130), .S0 (nx7720)) ;
    inv01 ix2129 (.Y (nx2130), .A (L1_0_L2_3_G1_MINI_ALU_nx336)) ;
    mux21 L1_0_L2_3_G1_MINI_ALU_ix361 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_11), .A0 (
          L1_0_L2_3_G1_MINI_ALU_nx485), .A1 (nx2132), .S0 (nx7720)) ;
    inv01 ix2131 (.Y (nx2132), .A (L1_0_L2_3_G1_MINI_ALU_nx356)) ;
    mux21 L1_0_L2_3_G1_MINI_ALU_ix381 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_12), .A0 (
          L1_0_L2_3_G1_MINI_ALU_nx493), .A1 (nx2134), .S0 (nx7720)) ;
    inv01 ix2133 (.Y (nx2134), .A (L1_0_L2_3_G1_MINI_ALU_nx376)) ;
    mux21 L1_0_L2_3_G1_MINI_ALU_ix401 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_13), .A0 (
          L1_0_L2_3_G1_MINI_ALU_nx501), .A1 (nx2136), .S0 (nx7720)) ;
    inv01 ix2135 (.Y (nx2136), .A (L1_0_L2_3_G1_MINI_ALU_nx396)) ;
    mux21 L1_0_L2_3_G1_MINI_ALU_ix421 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_14), .A0 (
          L1_0_L2_3_G1_MINI_ALU_nx509), .A1 (nx2138), .S0 (nx7720)) ;
    inv01 ix2137 (.Y (nx2138), .A (L1_0_L2_3_G1_MINI_ALU_nx416)) ;
    mux21 L1_0_L2_3_G1_MINI_ALU_ix441 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_15), .A0 (
          L1_0_L2_3_G1_MINI_ALU_nx517), .A1 (nx2140), .S0 (nx7722)) ;
    inv01 ix2139 (.Y (nx2140), .A (L1_0_L2_3_G1_MINI_ALU_nx436)) ;
    mux21 L1_0_L2_3_G1_MINI_ALU_ix461 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_16), .A0 (nx2142), .A1 (nx2144
          ), .S0 (nx7722)) ;
    inv01 ix2141 (.Y (nx2142), .A (L1_0_L2_3_G1_MINI_ALU_BoothP_16)) ;
    inv01 ix2143 (.Y (nx2144), .A (L1_0_L2_3_G1_MINI_ALU_nx456)) ;
    nor02_2x L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix319 (.Y (
             L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642), .A0 (Start), .A1 (
             CalculatingBooth_dup_1084)) ;
    nor02_2x L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix85 (.Y (
             L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_0), .A0 (nx7732), .A1 (
             nx2146)) ;
    inv01 ix2145 (.Y (nx2146), .A (L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_1)) ;
    mux21 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix125 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_1), .A0 (nx2148), .A1 (
          nx2150), .S0 (nx7732)) ;
    inv01 ix2147 (.Y (nx2148), .A (L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_2)) ;
    inv01 ix2149 (.Y (nx2150), .A (WindowDin_0__3__0)) ;
    mux21 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix133 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_2), .A0 (nx2152), .A1 (
          nx2154), .S0 (nx7732)) ;
    inv01 ix2151 (.Y (nx2152), .A (L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_3)) ;
    inv01 ix2153 (.Y (nx2154), .A (WindowDin_0__3__1)) ;
    mux21 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix141 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_3), .A0 (nx2156), .A1 (
          nx2158), .S0 (nx7732)) ;
    inv01 ix2155 (.Y (nx2156), .A (L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_4)) ;
    inv01 ix2157 (.Y (nx2158), .A (WindowDin_0__3__2)) ;
    mux21 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix149 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_4), .A0 (nx2160), .A1 (
          nx2162), .S0 (nx7732)) ;
    inv01 ix2159 (.Y (nx2160), .A (L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_5)) ;
    inv01 ix2161 (.Y (nx2162), .A (WindowDin_0__3__3)) ;
    mux21 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix157 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_5), .A0 (nx2164), .A1 (
          nx2166), .S0 (nx7732)) ;
    inv01 ix2163 (.Y (nx2164), .A (L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_6)) ;
    inv01 ix2165 (.Y (nx2166), .A (WindowDin_0__3__4)) ;
    mux21 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix165 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_6), .A0 (nx2168), .A1 (
          nx2170), .S0 (nx7732)) ;
    inv01 ix2167 (.Y (nx2168), .A (L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_7)) ;
    inv01 ix2169 (.Y (nx2170), .A (WindowDin_0__3__5)) ;
    mux21 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix173 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_7), .A0 (nx2172), .A1 (
          nx2174), .S0 (nx7734)) ;
    inv01 ix2171 (.Y (nx2172), .A (L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_8)) ;
    inv01 ix2173 (.Y (nx2174), .A (WindowDin_0__3__6)) ;
    mux21 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix181 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_8), .A0 (nx2176), .A1 (
          nx2178), .S0 (nx7734)) ;
    inv01 ix2175 (.Y (nx2176), .A (L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_9)) ;
    inv01 ix2177 (.Y (nx2178), .A (WindowDin_0__3__7)) ;
    nor02_2x L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix89 (.Y (
             L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_9), .A0 (nx7734), .A1 (
             nx2180)) ;
    inv01 ix2179 (.Y (nx2180), .A (L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_10)
          ) ;
    nor02_2x L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix93 (.Y (
             L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_10), .A0 (nx7734), .A1 (
             nx2182)) ;
    inv01 ix2181 (.Y (nx2182), .A (L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_11)
          ) ;
    nor02_2x L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix97 (.Y (
             L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_11), .A0 (nx7734), .A1 (
             nx2184)) ;
    inv01 ix2183 (.Y (nx2184), .A (L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_12)
          ) ;
    nor02_2x L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix101 (.Y (
             L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_12), .A0 (nx7734), .A1 (
             nx2186)) ;
    inv01 ix2185 (.Y (nx2186), .A (L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_13)
          ) ;
    nor02_2x L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix105 (.Y (
             L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_13), .A0 (nx7734), .A1 (
             nx2188)) ;
    inv01 ix2187 (.Y (nx2188), .A (L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_14)
          ) ;
    nor02_2x L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix109 (.Y (
             L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_14), .A0 (nx7736), .A1 (
             nx2190)) ;
    inv01 ix2189 (.Y (nx2190), .A (L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_15)
          ) ;
    nor02_2x L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix113 (.Y (
             L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_15), .A0 (nx7736), .A1 (
             nx2192)) ;
    inv01 ix2191 (.Y (nx2192), .A (L1_0_L2_3_G1_MINI_ALU_BoothPBeforeShift_16)
          ) ;
    nor02_2x L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix117 (.Y (
             L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_16), .A0 (nx7736), .A1 (
             nx2192)) ;
    mux21 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix189 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BoothOperand_0), .A0 (nx2194), .A1 (nx2196), .S0 (
          nx7724)) ;
    inv01 ix2193 (.Y (nx2194), .A (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_0)) ;
    inv01 ix2195 (.Y (nx2196), .A (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_0)) ;
    mux21 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix197 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BoothOperand_1), .A0 (nx2198), .A1 (nx2200), .S0 (
          nx7724)) ;
    inv01 ix2197 (.Y (nx2198), .A (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_1)) ;
    inv01 ix2199 (.Y (nx2200), .A (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_1)) ;
    mux21 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix205 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BoothOperand_2), .A0 (nx2202), .A1 (nx2204), .S0 (
          nx7724)) ;
    inv01 ix2201 (.Y (nx2202), .A (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_2)) ;
    inv01 ix2203 (.Y (nx2204), .A (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_2)) ;
    mux21 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix213 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BoothOperand_3), .A0 (nx2206), .A1 (nx2208), .S0 (
          nx7724)) ;
    inv01 ix2205 (.Y (nx2206), .A (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_3)) ;
    inv01 ix2207 (.Y (nx2208), .A (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_3)) ;
    mux21 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix221 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BoothOperand_4), .A0 (nx2210), .A1 (nx2212), .S0 (
          nx7724)) ;
    inv01 ix2209 (.Y (nx2210), .A (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_4)) ;
    inv01 ix2211 (.Y (nx2212), .A (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_4)) ;
    mux21 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix229 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BoothOperand_5), .A0 (nx2214), .A1 (nx2216), .S0 (
          nx7726)) ;
    inv01 ix2213 (.Y (nx2214), .A (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_5)) ;
    inv01 ix2215 (.Y (nx2216), .A (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_5)) ;
    mux21 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix237 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BoothOperand_6), .A0 (nx2218), .A1 (nx2220), .S0 (
          nx7726)) ;
    inv01 ix2217 (.Y (nx2218), .A (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_6)) ;
    inv01 ix2219 (.Y (nx2220), .A (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_6)) ;
    mux21 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix245 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BoothOperand_7), .A0 (nx2222), .A1 (nx2224), .S0 (
          nx7726)) ;
    inv01 ix2221 (.Y (nx2222), .A (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_7)) ;
    inv01 ix2223 (.Y (nx2224), .A (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_7)) ;
    mux21 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix253 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BoothOperand_8), .A0 (nx2226), .A1 (nx2228), .S0 (
          nx7726)) ;
    inv01 ix2225 (.Y (nx2226), .A (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_8)) ;
    inv01 ix2227 (.Y (nx2228), .A (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_8)) ;
    mux21 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix261 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BoothOperand_9), .A0 (nx2230), .A1 (nx2232), .S0 (
          nx7726)) ;
    inv01 ix2229 (.Y (nx2230), .A (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_9)) ;
    inv01 ix2231 (.Y (nx2232), .A (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_9)) ;
    mux21 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix269 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BoothOperand_10), .A0 (nx2234), .A1 (nx2236), .S0 (
          nx7726)) ;
    inv01 ix2233 (.Y (nx2234), .A (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_10)) ;
    inv01 ix2235 (.Y (nx2236), .A (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_10)) ;
    mux21 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix277 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BoothOperand_11), .A0 (nx2238), .A1 (nx2240), .S0 (
          nx7726)) ;
    inv01 ix2237 (.Y (nx2238), .A (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_11)) ;
    inv01 ix2239 (.Y (nx2240), .A (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_11)) ;
    mux21 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix285 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BoothOperand_12), .A0 (nx2242), .A1 (nx2244), .S0 (
          nx7728)) ;
    inv01 ix2241 (.Y (nx2242), .A (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_12)) ;
    inv01 ix2243 (.Y (nx2244), .A (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_12)) ;
    mux21 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix293 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BoothOperand_13), .A0 (nx2246), .A1 (nx2248), .S0 (
          nx7728)) ;
    inv01 ix2245 (.Y (nx2246), .A (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_13)) ;
    inv01 ix2247 (.Y (nx2248), .A (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_13)) ;
    mux21 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix301 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BoothOperand_14), .A0 (nx2250), .A1 (nx2252), .S0 (
          nx7728)) ;
    inv01 ix2249 (.Y (nx2250), .A (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_14)) ;
    inv01 ix2251 (.Y (nx2252), .A (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_14)) ;
    mux21 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix309 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BoothOperand_15), .A0 (nx2254), .A1 (nx2256), .S0 (
          nx7728)) ;
    inv01 ix2253 (.Y (nx2254), .A (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_15)) ;
    inv01 ix2255 (.Y (nx2256), .A (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_15)) ;
    mux21 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix317 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BoothOperand_16), .A0 (nx2258), .A1 (nx2260), .S0 (
          nx7728)) ;
    inv01 ix2257 (.Y (nx2258), .A (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_16)) ;
    inv01 ix2259 (.Y (nx2260), .A (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_16)) ;
    xnor2 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix321 (.Y (
          L1_0_L2_3_G1_MINI_ALU_AddPToBoothOperand), .A0 (nx7728), .A1 (nx2126)
          ) ;
    oai32 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix393 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .A0 (nx8614), .A1 (
          RST), .A2 (nx7738), .B0 (nx2196), .B1 (nx2264)) ;
    oai32 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix403 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .A0 (nx8614), .A1 (
          RST), .A2 (nx7738), .B0 (nx2200), .B1 (nx2264)) ;
    oai32 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix413 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .A0 (nx8614), .A1 (
          RST), .A2 (nx7738), .B0 (nx2204), .B1 (nx2264)) ;
    oai32 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix423 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .A0 (nx8614), .A1 (
          RST), .A2 (nx7738), .B0 (nx2208), .B1 (nx2264)) ;
    oai32 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix433 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .A0 (nx8614), .A1 (
          RST), .A2 (nx7738), .B0 (nx2212), .B1 (nx2264)) ;
    oai32 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix443 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .A0 (nx8614), .A1 (
          RST), .A2 (nx7738), .B0 (nx2216), .B1 (nx2264)) ;
    oai32 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix453 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .A0 (nx8614), .A1 (
          RST), .A2 (nx7740), .B0 (nx2220), .B1 (nx2264)) ;
    oai32 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix463 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .A0 (nx8616), .A1 (
          RST), .A2 (nx7740), .B0 (nx2224), .B1 (nx2266)) ;
    oai32 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix473 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .A0 (nx8616), .A1 (
          RST), .A2 (nx7740), .B0 (nx2228), .B1 (nx2266)) ;
    oai32 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix483 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .A0 (nx2268), .A1 (
          RST), .A2 (nx7740), .B0 (nx2232), .B1 (nx2266)) ;
    inv01 ix2267 (.Y (nx2268), .A (FilterDin_0__3__0)) ;
    oai32 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix493 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .A0 (nx2270), .A1 (
          RST), .A2 (nx7740), .B0 (nx2236), .B1 (nx2266)) ;
    inv01 ix2269 (.Y (nx2270), .A (FilterDin_0__3__1)) ;
    oai32 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix503 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .A0 (nx2272), .A1 (
          RST), .A2 (nx7740), .B0 (nx2240), .B1 (nx2266)) ;
    inv01 ix2271 (.Y (nx2272), .A (FilterDin_0__3__2)) ;
    oai32 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix513 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .A0 (nx2274), .A1 (
          RST), .A2 (nx7740), .B0 (nx2244), .B1 (nx2266)) ;
    inv01 ix2273 (.Y (nx2274), .A (FilterDin_0__3__3)) ;
    oai32 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix523 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .A0 (nx2276), .A1 (
          RST), .A2 (nx7742), .B0 (nx2248), .B1 (nx2266)) ;
    inv01 ix2275 (.Y (nx2276), .A (FilterDin_0__3__4)) ;
    oai32 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix533 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .A0 (nx2278), .A1 (
          RST), .A2 (nx7742), .B0 (nx2252), .B1 (nx2280)) ;
    inv01 ix2277 (.Y (nx2278), .A (FilterDin_0__3__5)) ;
    inv01 ix2279 (.Y (nx2280), .A (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566)) ;
    oai32 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix543 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .A0 (nx2282), .A1 (
          RST), .A2 (nx7742), .B0 (nx2256), .B1 (nx2280)) ;
    inv01 ix2281 (.Y (nx2282), .A (FilterDin_0__3__6)) ;
    oai32 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix553 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .A0 (nx2284), .A1 (
          RST), .A2 (nx7742), .B0 (nx2260), .B1 (nx2280)) ;
    inv01 ix2283 (.Y (nx2284), .A (FilterDin_0__3__7)) ;
    nand02_2x L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix633 (.Y (nx2264), .A0 (
              nx7580), .A1 (nx7742)) ;
    nand02_2x L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix635 (.Y (nx2266), .A0 (
              nx7580), .A1 (nx7742)) ;
    oai32 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix393 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .A0 (nx8616), .A1 (
          RST), .A2 (nx7744), .B0 (nx2194), .B1 (nx2286)) ;
    oai32 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix403 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .A0 (nx8616), .A1 (
          RST), .A2 (nx7744), .B0 (nx2198), .B1 (nx2286)) ;
    oai32 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix413 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .A0 (nx8616), .A1 (
          RST), .A2 (nx7744), .B0 (nx2202), .B1 (nx2286)) ;
    oai32 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix423 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .A0 (nx8616), .A1 (
          RST), .A2 (nx7744), .B0 (nx2206), .B1 (nx2286)) ;
    oai32 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix433 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .A0 (nx8616), .A1 (
          RST), .A2 (nx7744), .B0 (nx2210), .B1 (nx2286)) ;
    oai32 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix443 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .A0 (nx8618), .A1 (
          RST), .A2 (nx7744), .B0 (nx2214), .B1 (nx2286)) ;
    oai32 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix453 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .A0 (nx8618), .A1 (
          RST), .A2 (nx7746), .B0 (nx2218), .B1 (nx2286)) ;
    oai32 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix463 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .A0 (nx8618), .A1 (
          RST), .A2 (nx7746), .B0 (nx2222), .B1 (nx2288)) ;
    oai32 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix473 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .A0 (nx8618), .A1 (
          RST), .A2 (nx7746), .B0 (nx2226), .B1 (nx2288)) ;
    oai32 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix483 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .A0 (nx2268), .A1 (
          RST), .A2 (nx7746), .B0 (nx2230), .B1 (nx2288)) ;
    oai32 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix493 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .A0 (nx2290), .A1 (
          RST), .A2 (nx7746), .B0 (nx2234), .B1 (nx2288)) ;
    inv01 ix2289 (.Y (nx2290), .A (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_10)) ;
    oai32 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix503 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .A0 (nx2292), .A1 (
          RST), .A2 (nx7746), .B0 (nx2238), .B1 (nx2288)) ;
    inv01 ix2291 (.Y (nx2292), .A (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_11)) ;
    oai32 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix513 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .A0 (nx2294), .A1 (
          RST), .A2 (nx7746), .B0 (nx2242), .B1 (nx2288)) ;
    inv01 ix2293 (.Y (nx2294), .A (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_12)) ;
    oai32 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix523 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .A0 (nx2296), .A1 (
          RST), .A2 (nx7748), .B0 (nx2246), .B1 (nx2288)) ;
    inv01 ix2295 (.Y (nx2296), .A (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_13)) ;
    oai32 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix533 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .A0 (nx2298), .A1 (
          RST), .A2 (nx7748), .B0 (nx2250), .B1 (nx2300)) ;
    inv01 ix2297 (.Y (nx2298), .A (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_14)) ;
    inv01 ix2299 (.Y (nx2300), .A (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566)) ;
    oai32 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix543 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .A0 (nx2302), .A1 (
          RST), .A2 (nx7748), .B0 (nx2254), .B1 (nx2300)) ;
    inv01 ix2301 (.Y (nx2302), .A (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_15)) ;
    oai32 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix553 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .A0 (nx2304), .A1 (
          RST), .A2 (nx7748), .B0 (nx2258), .B1 (nx2300)) ;
    inv01 ix2303 (.Y (nx2304), .A (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_16)) ;
    nand02_2x L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix633 (.Y (nx2286), .A0 (
              nx7580), .A1 (nx7748)) ;
    nand02_2x L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix635 (.Y (nx2288), .A0 (
              nx7582), .A1 (nx7748)) ;
    oai32 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix393 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .A0 (nx2306), .A1 (
          RST), .A2 (nx7750), .B0 (L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx384), .B1 (
          nx2308)) ;
    inv01 ix2305 (.Y (nx2306), .A (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_0)) ;
    oai32 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix403 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .A0 (nx2310), .A1 (
          RST), .A2 (nx7750), .B0 (nx2126), .B1 (nx2308)) ;
    inv01 ix2309 (.Y (nx2310), .A (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_1)) ;
    oai32 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix413 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .A0 (nx2312), .A1 (
          RST), .A2 (nx7750), .B0 (L1_0_L2_3_G1_MINI_ALU_nx387), .B1 (nx2308)) ;
    inv01 ix2311 (.Y (nx2312), .A (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_2)) ;
    oai32 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix423 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .A0 (nx2314), .A1 (
          RST), .A2 (nx7750), .B0 (L1_0_L2_3_G1_MINI_ALU_nx399), .B1 (nx2308)) ;
    inv01 ix2313 (.Y (nx2314), .A (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_3)) ;
    oai32 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix433 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .A0 (nx2316), .A1 (
          RST), .A2 (nx7750), .B0 (L1_0_L2_3_G1_MINI_ALU_nx409), .B1 (nx2308)) ;
    inv01 ix2315 (.Y (nx2316), .A (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_4)) ;
    oai32 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix443 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .A0 (nx2318), .A1 (
          RST), .A2 (nx7750), .B0 (L1_0_L2_3_G1_MINI_ALU_nx419), .B1 (nx2308)) ;
    inv01 ix2317 (.Y (nx2318), .A (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_5)) ;
    oai32 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix453 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .A0 (nx2320), .A1 (
          RST), .A2 (nx7750), .B0 (L1_0_L2_3_G1_MINI_ALU_nx429), .B1 (nx2308)) ;
    inv01 ix2319 (.Y (nx2320), .A (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_6)) ;
    oai32 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix463 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .A0 (nx2322), .A1 (
          RST), .A2 (nx7752), .B0 (L1_0_L2_3_G1_MINI_ALU_nx439), .B1 (nx2324)) ;
    inv01 ix2321 (.Y (nx2322), .A (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_7)) ;
    oai32 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix473 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .A0 (nx2326), .A1 (
          RST), .A2 (nx7752), .B0 (L1_0_L2_3_G1_MINI_ALU_nx449), .B1 (nx2324)) ;
    inv01 ix2325 (.Y (nx2326), .A (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_8)) ;
    oai32 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix483 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .A0 (nx2328), .A1 (
          RST), .A2 (nx7752), .B0 (L1_0_L2_3_G1_MINI_ALU_nx469), .B1 (nx2324)) ;
    inv01 ix2327 (.Y (nx2328), .A (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_9)) ;
    oai32 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix493 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .A0 (nx2330), .A1 (
          RST), .A2 (nx7752), .B0 (L1_0_L2_3_G1_MINI_ALU_nx477), .B1 (nx2324)) ;
    inv01 ix2329 (.Y (nx2330), .A (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_10)) ;
    oai32 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix503 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .A0 (nx2332), .A1 (
          RST), .A2 (nx7752), .B0 (L1_0_L2_3_G1_MINI_ALU_nx485), .B1 (nx2324)) ;
    inv01 ix2331 (.Y (nx2332), .A (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_11)) ;
    oai32 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix513 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .A0 (nx2334), .A1 (
          RST), .A2 (nx7752), .B0 (L1_0_L2_3_G1_MINI_ALU_nx493), .B1 (nx2324)) ;
    inv01 ix2333 (.Y (nx2334), .A (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_12)) ;
    oai32 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix523 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .A0 (nx2336), .A1 (
          RST), .A2 (nx7752), .B0 (L1_0_L2_3_G1_MINI_ALU_nx501), .B1 (nx2324)) ;
    inv01 ix2335 (.Y (nx2336), .A (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_13)) ;
    oai32 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix533 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .A0 (nx2338), .A1 (
          RST), .A2 (nx7754), .B0 (L1_0_L2_3_G1_MINI_ALU_nx509), .B1 (nx2340)) ;
    inv01 ix2337 (.Y (nx2338), .A (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_14)) ;
    inv01 ix2339 (.Y (nx2340), .A (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566)) ;
    oai32 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix543 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .A0 (nx2342), .A1 (
          RST), .A2 (nx7754), .B0 (L1_0_L2_3_G1_MINI_ALU_nx517), .B1 (nx2340)) ;
    inv01 ix2341 (.Y (nx2342), .A (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_15)) ;
    oai32 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix553 (.Y (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .A0 (nx2344), .A1 (
          RST), .A2 (nx7754), .B0 (nx2142), .B1 (nx2340)) ;
    inv01 ix2343 (.Y (nx2344), .A (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_16)) ;
    nand02_2x L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix633 (.Y (nx2308), .A0 (
              nx7582), .A1 (nx7754)) ;
    nand02_2x L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix635 (.Y (nx2324), .A0 (
              nx7582), .A1 (nx7754)) ;
    mux21 L1_0_L2_4_G1_MINI_ALU_ix404 (.Y (L1_0_L2_4_G1_MINI_ALU_nx403), .A0 (
          nx2346), .A1 (L1_0_L2_4_G1_MINI_ALU_BoothP_2), .S0 (
          L1_0_L2_4_G1_MINI_ALU_nx395)) ;
    inv01 ix2345 (.Y (nx2346), .A (L1_0_L2_4_G1_MINI_ALU_nx391)) ;
    mux21 L1_0_L2_4_G1_MINI_ALU_ix414 (.Y (L1_0_L2_4_G1_MINI_ALU_nx413), .A0 (
          nx2348), .A1 (L1_0_L2_4_G1_MINI_ALU_BoothP_3), .S0 (
          L1_0_L2_4_G1_MINI_ALU_nx405)) ;
    inv01 ix2347 (.Y (nx2348), .A (L1_0_L2_4_G1_MINI_ALU_nx403)) ;
    mux21 L1_0_L2_4_G1_MINI_ALU_ix424 (.Y (L1_0_L2_4_G1_MINI_ALU_nx423), .A0 (
          nx2350), .A1 (L1_0_L2_4_G1_MINI_ALU_BoothP_4), .S0 (
          L1_0_L2_4_G1_MINI_ALU_nx415)) ;
    inv01 ix2349 (.Y (nx2350), .A (L1_0_L2_4_G1_MINI_ALU_nx413)) ;
    mux21 L1_0_L2_4_G1_MINI_ALU_ix434 (.Y (L1_0_L2_4_G1_MINI_ALU_nx433), .A0 (
          nx2352), .A1 (L1_0_L2_4_G1_MINI_ALU_BoothP_5), .S0 (
          L1_0_L2_4_G1_MINI_ALU_nx425)) ;
    inv01 ix2351 (.Y (nx2352), .A (L1_0_L2_4_G1_MINI_ALU_nx423)) ;
    mux21 L1_0_L2_4_G1_MINI_ALU_ix444 (.Y (L1_0_L2_4_G1_MINI_ALU_nx443), .A0 (
          nx2354), .A1 (L1_0_L2_4_G1_MINI_ALU_BoothP_6), .S0 (
          L1_0_L2_4_G1_MINI_ALU_nx435)) ;
    inv01 ix2353 (.Y (nx2354), .A (L1_0_L2_4_G1_MINI_ALU_nx433)) ;
    mux21 L1_0_L2_4_G1_MINI_ALU_ix454 (.Y (L1_0_L2_4_G1_MINI_ALU_nx453), .A0 (
          nx2356), .A1 (L1_0_L2_4_G1_MINI_ALU_BoothP_7), .S0 (
          L1_0_L2_4_G1_MINI_ALU_nx445)) ;
    inv01 ix2355 (.Y (nx2356), .A (L1_0_L2_4_G1_MINI_ALU_nx443)) ;
    mux21 L1_0_L2_4_G1_MINI_ALU_ix462 (.Y (L1_0_L2_4_G1_MINI_ALU_nx461), .A0 (
          nx2358), .A1 (L1_0_L2_4_G1_MINI_ALU_BoothP_8), .S0 (
          L1_0_L2_4_G1_MINI_ALU_nx455)) ;
    inv01 ix2357 (.Y (nx2358), .A (L1_0_L2_4_G1_MINI_ALU_nx453)) ;
    mux21 L1_0_L2_4_G1_MINI_ALU_ix468 (.Y (L1_0_L2_4_G1_MINI_ALU_nx467), .A0 (
          nx2360), .A1 (L1_0_L2_4_G1_MINI_ALU_BoothP_9), .S0 (
          L1_0_L2_4_G1_MINI_ALU_nx463)) ;
    inv01 ix2359 (.Y (nx2360), .A (L1_0_L2_4_G1_MINI_ALU_nx461)) ;
    mux21 L1_0_L2_4_G1_MINI_ALU_ix476 (.Y (L1_0_L2_4_G1_MINI_ALU_nx475), .A0 (
          nx2362), .A1 (L1_0_L2_4_G1_MINI_ALU_BoothP_10), .S0 (
          L1_0_L2_4_G1_MINI_ALU_nx471)) ;
    inv01 ix2361 (.Y (nx2362), .A (L1_0_L2_4_G1_MINI_ALU_nx467)) ;
    mux21 L1_0_L2_4_G1_MINI_ALU_ix484 (.Y (L1_0_L2_4_G1_MINI_ALU_nx483), .A0 (
          nx2364), .A1 (L1_0_L2_4_G1_MINI_ALU_BoothP_11), .S0 (
          L1_0_L2_4_G1_MINI_ALU_nx479)) ;
    inv01 ix2363 (.Y (nx2364), .A (L1_0_L2_4_G1_MINI_ALU_nx475)) ;
    mux21 L1_0_L2_4_G1_MINI_ALU_ix492 (.Y (L1_0_L2_4_G1_MINI_ALU_nx491), .A0 (
          nx2366), .A1 (L1_0_L2_4_G1_MINI_ALU_BoothP_12), .S0 (
          L1_0_L2_4_G1_MINI_ALU_nx487)) ;
    inv01 ix2365 (.Y (nx2366), .A (L1_0_L2_4_G1_MINI_ALU_nx483)) ;
    mux21 L1_0_L2_4_G1_MINI_ALU_ix500 (.Y (L1_0_L2_4_G1_MINI_ALU_nx499), .A0 (
          nx2368), .A1 (L1_0_L2_4_G1_MINI_ALU_BoothP_13), .S0 (
          L1_0_L2_4_G1_MINI_ALU_nx495)) ;
    inv01 ix2367 (.Y (nx2368), .A (L1_0_L2_4_G1_MINI_ALU_nx491)) ;
    mux21 L1_0_L2_4_G1_MINI_ALU_ix508 (.Y (L1_0_L2_4_G1_MINI_ALU_nx507), .A0 (
          nx2370), .A1 (L1_0_L2_4_G1_MINI_ALU_BoothP_14), .S0 (
          L1_0_L2_4_G1_MINI_ALU_nx503)) ;
    inv01 ix2369 (.Y (nx2370), .A (L1_0_L2_4_G1_MINI_ALU_nx499)) ;
    mux21 L1_0_L2_4_G1_MINI_ALU_ix516 (.Y (L1_0_L2_4_G1_MINI_ALU_nx515), .A0 (
          nx2372), .A1 (L1_0_L2_4_G1_MINI_ALU_BoothP_15), .S0 (
          L1_0_L2_4_G1_MINI_ALU_nx511)) ;
    inv01 ix2371 (.Y (nx2372), .A (L1_0_L2_4_G1_MINI_ALU_nx507)) ;
    mux21 L1_0_L2_4_G1_MINI_ALU_ix161 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_1), .A0 (nx2374), .A1 (
          L1_0_L2_4_G1_MINI_ALU_nx379), .S0 (nx7758)) ;
    inv01 ix2373 (.Y (nx2374), .A (L1_0_L2_4_G1_MINI_ALU_BoothP_1)) ;
    mux21 L1_0_L2_4_G1_MINI_ALU_ix181 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_2), .A0 (
          L1_0_L2_4_G1_MINI_ALU_nx387), .A1 (L1_0_L2_4_G1_MINI_ALU_nx389), .S0 (
          nx7758)) ;
    mux21 L1_0_L2_4_G1_MINI_ALU_ix201 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_3), .A0 (
          L1_0_L2_4_G1_MINI_ALU_nx399), .A1 (L1_0_L2_4_G1_MINI_ALU_nx401), .S0 (
          nx7758)) ;
    mux21 L1_0_L2_4_G1_MINI_ALU_ix221 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_4), .A0 (
          L1_0_L2_4_G1_MINI_ALU_nx409), .A1 (L1_0_L2_4_G1_MINI_ALU_nx411), .S0 (
          nx7758)) ;
    mux21 L1_0_L2_4_G1_MINI_ALU_ix241 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_5), .A0 (
          L1_0_L2_4_G1_MINI_ALU_nx419), .A1 (L1_0_L2_4_G1_MINI_ALU_nx421), .S0 (
          nx7758)) ;
    mux21 L1_0_L2_4_G1_MINI_ALU_ix261 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_6), .A0 (
          L1_0_L2_4_G1_MINI_ALU_nx429), .A1 (L1_0_L2_4_G1_MINI_ALU_nx431), .S0 (
          nx7758)) ;
    mux21 L1_0_L2_4_G1_MINI_ALU_ix281 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_7), .A0 (
          L1_0_L2_4_G1_MINI_ALU_nx439), .A1 (L1_0_L2_4_G1_MINI_ALU_nx441), .S0 (
          nx7758)) ;
    mux21 L1_0_L2_4_G1_MINI_ALU_ix301 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_8), .A0 (
          L1_0_L2_4_G1_MINI_ALU_nx449), .A1 (L1_0_L2_4_G1_MINI_ALU_nx451), .S0 (
          nx7760)) ;
    mux21 L1_0_L2_4_G1_MINI_ALU_ix321 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_9), .A0 (
          L1_0_L2_4_G1_MINI_ALU_nx469), .A1 (nx2376), .S0 (nx7760)) ;
    inv01 ix2375 (.Y (nx2376), .A (L1_0_L2_4_G1_MINI_ALU_nx316)) ;
    mux21 L1_0_L2_4_G1_MINI_ALU_ix341 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_10), .A0 (
          L1_0_L2_4_G1_MINI_ALU_nx477), .A1 (nx2378), .S0 (nx7760)) ;
    inv01 ix2377 (.Y (nx2378), .A (L1_0_L2_4_G1_MINI_ALU_nx336)) ;
    mux21 L1_0_L2_4_G1_MINI_ALU_ix361 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_11), .A0 (
          L1_0_L2_4_G1_MINI_ALU_nx485), .A1 (nx2380), .S0 (nx7760)) ;
    inv01 ix2379 (.Y (nx2380), .A (L1_0_L2_4_G1_MINI_ALU_nx356)) ;
    mux21 L1_0_L2_4_G1_MINI_ALU_ix381 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_12), .A0 (
          L1_0_L2_4_G1_MINI_ALU_nx493), .A1 (nx2382), .S0 (nx7760)) ;
    inv01 ix2381 (.Y (nx2382), .A (L1_0_L2_4_G1_MINI_ALU_nx376)) ;
    mux21 L1_0_L2_4_G1_MINI_ALU_ix401 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_13), .A0 (
          L1_0_L2_4_G1_MINI_ALU_nx501), .A1 (nx2384), .S0 (nx7760)) ;
    inv01 ix2383 (.Y (nx2384), .A (L1_0_L2_4_G1_MINI_ALU_nx396)) ;
    mux21 L1_0_L2_4_G1_MINI_ALU_ix421 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_14), .A0 (
          L1_0_L2_4_G1_MINI_ALU_nx509), .A1 (nx2386), .S0 (nx7760)) ;
    inv01 ix2385 (.Y (nx2386), .A (L1_0_L2_4_G1_MINI_ALU_nx416)) ;
    mux21 L1_0_L2_4_G1_MINI_ALU_ix441 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_15), .A0 (
          L1_0_L2_4_G1_MINI_ALU_nx517), .A1 (nx2388), .S0 (nx7762)) ;
    inv01 ix2387 (.Y (nx2388), .A (L1_0_L2_4_G1_MINI_ALU_nx436)) ;
    mux21 L1_0_L2_4_G1_MINI_ALU_ix461 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_16), .A0 (nx2390), .A1 (nx2392
          ), .S0 (nx7762)) ;
    inv01 ix2389 (.Y (nx2390), .A (L1_0_L2_4_G1_MINI_ALU_BoothP_16)) ;
    inv01 ix2391 (.Y (nx2392), .A (L1_0_L2_4_G1_MINI_ALU_nx456)) ;
    nor02_2x L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix319 (.Y (
             L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642), .A0 (Start), .A1 (
             CalculatingBooth_dup_1084)) ;
    nor02_2x L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix85 (.Y (
             L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_0), .A0 (nx7772), .A1 (
             nx2394)) ;
    inv01 ix2393 (.Y (nx2394), .A (L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_1)) ;
    mux21 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix125 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_1), .A0 (nx2396), .A1 (
          nx2398), .S0 (nx7772)) ;
    inv01 ix2395 (.Y (nx2396), .A (L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_2)) ;
    inv01 ix2397 (.Y (nx2398), .A (WindowDin_0__4__0)) ;
    mux21 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix133 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_2), .A0 (nx2400), .A1 (
          nx2402), .S0 (nx7772)) ;
    inv01 ix2399 (.Y (nx2400), .A (L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_3)) ;
    inv01 ix2401 (.Y (nx2402), .A (WindowDin_0__4__1)) ;
    mux21 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix141 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_3), .A0 (nx2404), .A1 (
          nx2406), .S0 (nx7772)) ;
    inv01 ix2403 (.Y (nx2404), .A (L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_4)) ;
    inv01 ix2405 (.Y (nx2406), .A (WindowDin_0__4__2)) ;
    mux21 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix149 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_4), .A0 (nx2408), .A1 (
          nx2410), .S0 (nx7772)) ;
    inv01 ix2407 (.Y (nx2408), .A (L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_5)) ;
    inv01 ix2409 (.Y (nx2410), .A (WindowDin_0__4__3)) ;
    mux21 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix157 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_5), .A0 (nx2412), .A1 (
          nx2414), .S0 (nx7772)) ;
    inv01 ix2411 (.Y (nx2412), .A (L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_6)) ;
    inv01 ix2413 (.Y (nx2414), .A (WindowDin_0__4__4)) ;
    mux21 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix165 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_6), .A0 (nx2416), .A1 (
          nx2418), .S0 (nx7772)) ;
    inv01 ix2415 (.Y (nx2416), .A (L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_7)) ;
    inv01 ix2417 (.Y (nx2418), .A (WindowDin_0__4__5)) ;
    mux21 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix173 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_7), .A0 (nx2420), .A1 (
          nx2422), .S0 (nx7774)) ;
    inv01 ix2419 (.Y (nx2420), .A (L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_8)) ;
    inv01 ix2421 (.Y (nx2422), .A (WindowDin_0__4__6)) ;
    mux21 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix181 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_8), .A0 (nx2424), .A1 (
          nx2426), .S0 (nx7774)) ;
    inv01 ix2423 (.Y (nx2424), .A (L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_9)) ;
    inv01 ix2425 (.Y (nx2426), .A (WindowDin_0__4__7)) ;
    nor02_2x L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix89 (.Y (
             L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_9), .A0 (nx7774), .A1 (
             nx2428)) ;
    inv01 ix2427 (.Y (nx2428), .A (L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_10)
          ) ;
    nor02_2x L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix93 (.Y (
             L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_10), .A0 (nx7774), .A1 (
             nx2430)) ;
    inv01 ix2429 (.Y (nx2430), .A (L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_11)
          ) ;
    nor02_2x L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix97 (.Y (
             L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_11), .A0 (nx7774), .A1 (
             nx2432)) ;
    inv01 ix2431 (.Y (nx2432), .A (L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_12)
          ) ;
    nor02_2x L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix101 (.Y (
             L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_12), .A0 (nx7774), .A1 (
             nx2434)) ;
    inv01 ix2433 (.Y (nx2434), .A (L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_13)
          ) ;
    nor02_2x L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix105 (.Y (
             L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_13), .A0 (nx7774), .A1 (
             nx2436)) ;
    inv01 ix2435 (.Y (nx2436), .A (L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_14)
          ) ;
    nor02_2x L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix109 (.Y (
             L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_14), .A0 (nx7776), .A1 (
             nx2438)) ;
    inv01 ix2437 (.Y (nx2438), .A (L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_15)
          ) ;
    nor02_2x L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix113 (.Y (
             L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_15), .A0 (nx7776), .A1 (
             nx2440)) ;
    inv01 ix2439 (.Y (nx2440), .A (L1_0_L2_4_G1_MINI_ALU_BoothPBeforeShift_16)
          ) ;
    nor02_2x L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix117 (.Y (
             L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_16), .A0 (nx7776), .A1 (
             nx2440)) ;
    mux21 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix189 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BoothOperand_0), .A0 (nx2442), .A1 (nx2444), .S0 (
          nx7764)) ;
    inv01 ix2441 (.Y (nx2442), .A (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_0)) ;
    inv01 ix2443 (.Y (nx2444), .A (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_0)) ;
    mux21 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix197 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BoothOperand_1), .A0 (nx2446), .A1 (nx2448), .S0 (
          nx7764)) ;
    inv01 ix2445 (.Y (nx2446), .A (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_1)) ;
    inv01 ix2447 (.Y (nx2448), .A (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_1)) ;
    mux21 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix205 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BoothOperand_2), .A0 (nx2450), .A1 (nx2452), .S0 (
          nx7764)) ;
    inv01 ix2449 (.Y (nx2450), .A (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_2)) ;
    inv01 ix2451 (.Y (nx2452), .A (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_2)) ;
    mux21 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix213 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BoothOperand_3), .A0 (nx2454), .A1 (nx2456), .S0 (
          nx7764)) ;
    inv01 ix2453 (.Y (nx2454), .A (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_3)) ;
    inv01 ix2455 (.Y (nx2456), .A (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_3)) ;
    mux21 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix221 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BoothOperand_4), .A0 (nx2458), .A1 (nx2460), .S0 (
          nx7764)) ;
    inv01 ix2457 (.Y (nx2458), .A (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_4)) ;
    inv01 ix2459 (.Y (nx2460), .A (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_4)) ;
    mux21 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix229 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BoothOperand_5), .A0 (nx2462), .A1 (nx2464), .S0 (
          nx7766)) ;
    inv01 ix2461 (.Y (nx2462), .A (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_5)) ;
    inv01 ix2463 (.Y (nx2464), .A (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_5)) ;
    mux21 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix237 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BoothOperand_6), .A0 (nx2466), .A1 (nx2468), .S0 (
          nx7766)) ;
    inv01 ix2465 (.Y (nx2466), .A (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_6)) ;
    inv01 ix2467 (.Y (nx2468), .A (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_6)) ;
    mux21 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix245 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BoothOperand_7), .A0 (nx2470), .A1 (nx2472), .S0 (
          nx7766)) ;
    inv01 ix2469 (.Y (nx2470), .A (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_7)) ;
    inv01 ix2471 (.Y (nx2472), .A (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_7)) ;
    mux21 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix253 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BoothOperand_8), .A0 (nx2474), .A1 (nx2476), .S0 (
          nx7766)) ;
    inv01 ix2473 (.Y (nx2474), .A (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_8)) ;
    inv01 ix2475 (.Y (nx2476), .A (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_8)) ;
    mux21 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix261 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BoothOperand_9), .A0 (nx2478), .A1 (nx2480), .S0 (
          nx7766)) ;
    inv01 ix2477 (.Y (nx2478), .A (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_9)) ;
    inv01 ix2479 (.Y (nx2480), .A (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_9)) ;
    mux21 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix269 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BoothOperand_10), .A0 (nx2482), .A1 (nx2484), .S0 (
          nx7766)) ;
    inv01 ix2481 (.Y (nx2482), .A (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_10)) ;
    inv01 ix2483 (.Y (nx2484), .A (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_10)) ;
    mux21 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix277 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BoothOperand_11), .A0 (nx2486), .A1 (nx2488), .S0 (
          nx7766)) ;
    inv01 ix2485 (.Y (nx2486), .A (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_11)) ;
    inv01 ix2487 (.Y (nx2488), .A (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_11)) ;
    mux21 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix285 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BoothOperand_12), .A0 (nx2490), .A1 (nx2492), .S0 (
          nx7768)) ;
    inv01 ix2489 (.Y (nx2490), .A (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_12)) ;
    inv01 ix2491 (.Y (nx2492), .A (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_12)) ;
    mux21 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix293 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BoothOperand_13), .A0 (nx2494), .A1 (nx2496), .S0 (
          nx7768)) ;
    inv01 ix2493 (.Y (nx2494), .A (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_13)) ;
    inv01 ix2495 (.Y (nx2496), .A (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_13)) ;
    mux21 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix301 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BoothOperand_14), .A0 (nx2498), .A1 (nx2500), .S0 (
          nx7768)) ;
    inv01 ix2497 (.Y (nx2498), .A (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_14)) ;
    inv01 ix2499 (.Y (nx2500), .A (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_14)) ;
    mux21 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix309 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BoothOperand_15), .A0 (nx2502), .A1 (nx2504), .S0 (
          nx7768)) ;
    inv01 ix2501 (.Y (nx2502), .A (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_15)) ;
    inv01 ix2503 (.Y (nx2504), .A (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_15)) ;
    mux21 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix317 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BoothOperand_16), .A0 (nx2506), .A1 (nx2508), .S0 (
          nx7768)) ;
    inv01 ix2505 (.Y (nx2506), .A (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_16)) ;
    inv01 ix2507 (.Y (nx2508), .A (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_16)) ;
    xnor2 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix321 (.Y (
          L1_0_L2_4_G1_MINI_ALU_AddPToBoothOperand), .A0 (nx7768), .A1 (nx2374)
          ) ;
    oai32 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix393 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .A0 (nx8620), .A1 (
          RST), .A2 (nx7778), .B0 (nx2444), .B1 (nx2512)) ;
    oai32 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix403 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .A0 (nx8620), .A1 (
          RST), .A2 (nx7778), .B0 (nx2448), .B1 (nx2512)) ;
    oai32 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix413 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .A0 (nx8620), .A1 (
          RST), .A2 (nx7778), .B0 (nx2452), .B1 (nx2512)) ;
    oai32 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix423 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .A0 (nx8620), .A1 (
          RST), .A2 (nx7778), .B0 (nx2456), .B1 (nx2512)) ;
    oai32 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix433 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .A0 (nx8620), .A1 (
          RST), .A2 (nx7778), .B0 (nx2460), .B1 (nx2512)) ;
    oai32 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix443 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .A0 (nx8620), .A1 (
          RST), .A2 (nx7778), .B0 (nx2464), .B1 (nx2512)) ;
    oai32 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix453 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .A0 (nx8620), .A1 (
          RST), .A2 (nx7780), .B0 (nx2468), .B1 (nx2512)) ;
    oai32 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix463 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .A0 (nx8622), .A1 (
          RST), .A2 (nx7780), .B0 (nx2472), .B1 (nx2514)) ;
    oai32 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix473 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .A0 (nx8622), .A1 (
          RST), .A2 (nx7780), .B0 (nx2476), .B1 (nx2514)) ;
    oai32 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix483 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .A0 (nx2516), .A1 (
          RST), .A2 (nx7780), .B0 (nx2480), .B1 (nx2514)) ;
    inv01 ix2515 (.Y (nx2516), .A (FilterDin_0__4__0)) ;
    oai32 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix493 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .A0 (nx2518), .A1 (
          RST), .A2 (nx7780), .B0 (nx2484), .B1 (nx2514)) ;
    inv01 ix2517 (.Y (nx2518), .A (FilterDin_0__4__1)) ;
    oai32 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix503 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .A0 (nx2520), .A1 (
          RST), .A2 (nx7780), .B0 (nx2488), .B1 (nx2514)) ;
    inv01 ix2519 (.Y (nx2520), .A (FilterDin_0__4__2)) ;
    oai32 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix513 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .A0 (nx2522), .A1 (
          RST), .A2 (nx7780), .B0 (nx2492), .B1 (nx2514)) ;
    inv01 ix2521 (.Y (nx2522), .A (FilterDin_0__4__3)) ;
    oai32 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix523 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .A0 (nx2524), .A1 (
          RST), .A2 (nx7782), .B0 (nx2496), .B1 (nx2514)) ;
    inv01 ix2523 (.Y (nx2524), .A (FilterDin_0__4__4)) ;
    oai32 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix533 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .A0 (nx2526), .A1 (
          RST), .A2 (nx7782), .B0 (nx2500), .B1 (nx2528)) ;
    inv01 ix2525 (.Y (nx2526), .A (FilterDin_0__4__5)) ;
    inv01 ix2527 (.Y (nx2528), .A (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566)) ;
    oai32 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix543 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .A0 (nx2530), .A1 (
          RST), .A2 (nx7782), .B0 (nx2504), .B1 (nx2528)) ;
    inv01 ix2529 (.Y (nx2530), .A (FilterDin_0__4__6)) ;
    oai32 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix553 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .A0 (nx2532), .A1 (
          RST), .A2 (nx7782), .B0 (nx2508), .B1 (nx2528)) ;
    inv01 ix2531 (.Y (nx2532), .A (FilterDin_0__4__7)) ;
    nand02_2x L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix633 (.Y (nx2512), .A0 (
              nx7582), .A1 (nx7782)) ;
    nand02_2x L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix635 (.Y (nx2514), .A0 (
              nx7582), .A1 (nx7782)) ;
    oai32 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix393 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .A0 (nx8622), .A1 (
          RST), .A2 (nx7784), .B0 (nx2442), .B1 (nx2534)) ;
    oai32 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix403 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .A0 (nx8622), .A1 (
          RST), .A2 (nx7784), .B0 (nx2446), .B1 (nx2534)) ;
    oai32 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix413 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .A0 (nx8622), .A1 (
          RST), .A2 (nx7784), .B0 (nx2450), .B1 (nx2534)) ;
    oai32 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix423 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .A0 (nx8622), .A1 (
          RST), .A2 (nx7784), .B0 (nx2454), .B1 (nx2534)) ;
    oai32 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix433 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .A0 (nx8622), .A1 (
          RST), .A2 (nx7784), .B0 (nx2458), .B1 (nx2534)) ;
    oai32 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix443 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .A0 (nx8624), .A1 (
          RST), .A2 (nx7784), .B0 (nx2462), .B1 (nx2534)) ;
    oai32 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix453 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .A0 (nx8624), .A1 (
          RST), .A2 (nx7786), .B0 (nx2466), .B1 (nx2534)) ;
    oai32 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix463 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .A0 (nx8624), .A1 (
          RST), .A2 (nx7786), .B0 (nx2470), .B1 (nx2536)) ;
    oai32 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix473 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .A0 (nx8624), .A1 (
          RST), .A2 (nx7786), .B0 (nx2474), .B1 (nx2536)) ;
    oai32 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix483 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .A0 (nx2516), .A1 (
          RST), .A2 (nx7786), .B0 (nx2478), .B1 (nx2536)) ;
    oai32 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix493 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .A0 (nx2538), .A1 (
          RST), .A2 (nx7786), .B0 (nx2482), .B1 (nx2536)) ;
    inv01 ix2537 (.Y (nx2538), .A (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_10)) ;
    oai32 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix503 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .A0 (nx2540), .A1 (
          RST), .A2 (nx7786), .B0 (nx2486), .B1 (nx2536)) ;
    inv01 ix2539 (.Y (nx2540), .A (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_11)) ;
    oai32 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix513 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .A0 (nx2542), .A1 (
          RST), .A2 (nx7786), .B0 (nx2490), .B1 (nx2536)) ;
    inv01 ix2541 (.Y (nx2542), .A (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_12)) ;
    oai32 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix523 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .A0 (nx2544), .A1 (
          RST), .A2 (nx7788), .B0 (nx2494), .B1 (nx2536)) ;
    inv01 ix2543 (.Y (nx2544), .A (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_13)) ;
    oai32 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix533 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .A0 (nx2546), .A1 (
          RST), .A2 (nx7788), .B0 (nx2498), .B1 (nx2548)) ;
    inv01 ix2545 (.Y (nx2546), .A (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_14)) ;
    inv01 ix2547 (.Y (nx2548), .A (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566)) ;
    oai32 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix543 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .A0 (nx2550), .A1 (
          RST), .A2 (nx7788), .B0 (nx2502), .B1 (nx2548)) ;
    inv01 ix2549 (.Y (nx2550), .A (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_15)) ;
    oai32 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix553 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .A0 (nx2552), .A1 (
          RST), .A2 (nx7788), .B0 (nx2506), .B1 (nx2548)) ;
    inv01 ix2551 (.Y (nx2552), .A (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_16)) ;
    nand02_2x L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix633 (.Y (nx2534), .A0 (
              nx7582), .A1 (nx7788)) ;
    nand02_2x L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix635 (.Y (nx2536), .A0 (
              nx7582), .A1 (nx7788)) ;
    oai32 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix393 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .A0 (nx2554), .A1 (
          RST), .A2 (nx7790), .B0 (L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx384), .B1 (
          nx2556)) ;
    inv01 ix2553 (.Y (nx2554), .A (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_0)) ;
    oai32 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix403 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .A0 (nx2558), .A1 (
          RST), .A2 (nx7790), .B0 (nx2374), .B1 (nx2556)) ;
    inv01 ix2557 (.Y (nx2558), .A (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_1)) ;
    oai32 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix413 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .A0 (nx2560), .A1 (
          RST), .A2 (nx7790), .B0 (L1_0_L2_4_G1_MINI_ALU_nx387), .B1 (nx2556)) ;
    inv01 ix2559 (.Y (nx2560), .A (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_2)) ;
    oai32 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix423 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .A0 (nx2562), .A1 (
          RST), .A2 (nx7790), .B0 (L1_0_L2_4_G1_MINI_ALU_nx399), .B1 (nx2556)) ;
    inv01 ix2561 (.Y (nx2562), .A (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_3)) ;
    oai32 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix433 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .A0 (nx2564), .A1 (
          RST), .A2 (nx7790), .B0 (L1_0_L2_4_G1_MINI_ALU_nx409), .B1 (nx2556)) ;
    inv01 ix2563 (.Y (nx2564), .A (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_4)) ;
    oai32 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix443 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .A0 (nx2566), .A1 (
          RST), .A2 (nx7790), .B0 (L1_0_L2_4_G1_MINI_ALU_nx419), .B1 (nx2556)) ;
    inv01 ix2565 (.Y (nx2566), .A (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_5)) ;
    oai32 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix453 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .A0 (nx2568), .A1 (
          RST), .A2 (nx7790), .B0 (L1_0_L2_4_G1_MINI_ALU_nx429), .B1 (nx2556)) ;
    inv01 ix2567 (.Y (nx2568), .A (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_6)) ;
    oai32 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix463 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .A0 (nx2570), .A1 (
          RST), .A2 (nx7792), .B0 (L1_0_L2_4_G1_MINI_ALU_nx439), .B1 (nx2572)) ;
    inv01 ix2569 (.Y (nx2570), .A (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_7)) ;
    oai32 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix473 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .A0 (nx2574), .A1 (
          RST), .A2 (nx7792), .B0 (L1_0_L2_4_G1_MINI_ALU_nx449), .B1 (nx2572)) ;
    inv01 ix2573 (.Y (nx2574), .A (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_8)) ;
    oai32 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix483 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .A0 (nx2576), .A1 (
          RST), .A2 (nx7792), .B0 (L1_0_L2_4_G1_MINI_ALU_nx469), .B1 (nx2572)) ;
    inv01 ix2575 (.Y (nx2576), .A (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_9)) ;
    oai32 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix493 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .A0 (nx2578), .A1 (
          RST), .A2 (nx7792), .B0 (L1_0_L2_4_G1_MINI_ALU_nx477), .B1 (nx2572)) ;
    inv01 ix2577 (.Y (nx2578), .A (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_10)) ;
    oai32 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix503 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .A0 (nx2580), .A1 (
          RST), .A2 (nx7792), .B0 (L1_0_L2_4_G1_MINI_ALU_nx485), .B1 (nx2572)) ;
    inv01 ix2579 (.Y (nx2580), .A (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_11)) ;
    oai32 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix513 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .A0 (nx2582), .A1 (
          RST), .A2 (nx7792), .B0 (L1_0_L2_4_G1_MINI_ALU_nx493), .B1 (nx2572)) ;
    inv01 ix2581 (.Y (nx2582), .A (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_12)) ;
    oai32 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix523 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .A0 (nx2584), .A1 (
          RST), .A2 (nx7792), .B0 (L1_0_L2_4_G1_MINI_ALU_nx501), .B1 (nx2572)) ;
    inv01 ix2583 (.Y (nx2584), .A (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_13)) ;
    oai32 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix533 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .A0 (nx2586), .A1 (
          RST), .A2 (nx7794), .B0 (L1_0_L2_4_G1_MINI_ALU_nx509), .B1 (nx2588)) ;
    inv01 ix2585 (.Y (nx2586), .A (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_14)) ;
    inv01 ix2587 (.Y (nx2588), .A (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566)) ;
    oai32 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix543 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .A0 (nx2590), .A1 (
          RST), .A2 (nx7794), .B0 (L1_0_L2_4_G1_MINI_ALU_nx517), .B1 (nx2588)) ;
    inv01 ix2589 (.Y (nx2590), .A (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_15)) ;
    oai32 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix553 (.Y (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .A0 (nx2592), .A1 (
          RST), .A2 (nx7794), .B0 (nx2390), .B1 (nx2588)) ;
    inv01 ix2591 (.Y (nx2592), .A (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_16)) ;
    nand02_2x L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix633 (.Y (nx2556), .A0 (
              nx7584), .A1 (nx7794)) ;
    nand02_2x L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix635 (.Y (nx2572), .A0 (
              nx7584), .A1 (nx7794)) ;
    mux21 L1_1_L2_0_G1_MINI_ALU_ix404 (.Y (L1_1_L2_0_G1_MINI_ALU_nx403), .A0 (
          nx2594), .A1 (L1_1_L2_0_G1_MINI_ALU_BoothP_2), .S0 (
          L1_1_L2_0_G1_MINI_ALU_nx395)) ;
    inv01 ix2593 (.Y (nx2594), .A (L1_1_L2_0_G1_MINI_ALU_nx391)) ;
    mux21 L1_1_L2_0_G1_MINI_ALU_ix414 (.Y (L1_1_L2_0_G1_MINI_ALU_nx413), .A0 (
          nx2596), .A1 (L1_1_L2_0_G1_MINI_ALU_BoothP_3), .S0 (
          L1_1_L2_0_G1_MINI_ALU_nx405)) ;
    inv01 ix2595 (.Y (nx2596), .A (L1_1_L2_0_G1_MINI_ALU_nx403)) ;
    mux21 L1_1_L2_0_G1_MINI_ALU_ix424 (.Y (L1_1_L2_0_G1_MINI_ALU_nx423), .A0 (
          nx2598), .A1 (L1_1_L2_0_G1_MINI_ALU_BoothP_4), .S0 (
          L1_1_L2_0_G1_MINI_ALU_nx415)) ;
    inv01 ix2597 (.Y (nx2598), .A (L1_1_L2_0_G1_MINI_ALU_nx413)) ;
    mux21 L1_1_L2_0_G1_MINI_ALU_ix434 (.Y (L1_1_L2_0_G1_MINI_ALU_nx433), .A0 (
          nx2600), .A1 (L1_1_L2_0_G1_MINI_ALU_BoothP_5), .S0 (
          L1_1_L2_0_G1_MINI_ALU_nx425)) ;
    inv01 ix2599 (.Y (nx2600), .A (L1_1_L2_0_G1_MINI_ALU_nx423)) ;
    mux21 L1_1_L2_0_G1_MINI_ALU_ix444 (.Y (L1_1_L2_0_G1_MINI_ALU_nx443), .A0 (
          nx2602), .A1 (L1_1_L2_0_G1_MINI_ALU_BoothP_6), .S0 (
          L1_1_L2_0_G1_MINI_ALU_nx435)) ;
    inv01 ix2601 (.Y (nx2602), .A (L1_1_L2_0_G1_MINI_ALU_nx433)) ;
    mux21 L1_1_L2_0_G1_MINI_ALU_ix454 (.Y (L1_1_L2_0_G1_MINI_ALU_nx453), .A0 (
          nx2604), .A1 (L1_1_L2_0_G1_MINI_ALU_BoothP_7), .S0 (
          L1_1_L2_0_G1_MINI_ALU_nx445)) ;
    inv01 ix2603 (.Y (nx2604), .A (L1_1_L2_0_G1_MINI_ALU_nx443)) ;
    mux21 L1_1_L2_0_G1_MINI_ALU_ix462 (.Y (L1_1_L2_0_G1_MINI_ALU_nx461), .A0 (
          nx2606), .A1 (L1_1_L2_0_G1_MINI_ALU_BoothP_8), .S0 (
          L1_1_L2_0_G1_MINI_ALU_nx455)) ;
    inv01 ix2605 (.Y (nx2606), .A (L1_1_L2_0_G1_MINI_ALU_nx453)) ;
    mux21 L1_1_L2_0_G1_MINI_ALU_ix468 (.Y (L1_1_L2_0_G1_MINI_ALU_nx467), .A0 (
          nx2608), .A1 (L1_1_L2_0_G1_MINI_ALU_BoothP_9), .S0 (
          L1_1_L2_0_G1_MINI_ALU_nx463)) ;
    inv01 ix2607 (.Y (nx2608), .A (L1_1_L2_0_G1_MINI_ALU_nx461)) ;
    mux21 L1_1_L2_0_G1_MINI_ALU_ix476 (.Y (L1_1_L2_0_G1_MINI_ALU_nx475), .A0 (
          nx2610), .A1 (L1_1_L2_0_G1_MINI_ALU_BoothP_10), .S0 (
          L1_1_L2_0_G1_MINI_ALU_nx471)) ;
    inv01 ix2609 (.Y (nx2610), .A (L1_1_L2_0_G1_MINI_ALU_nx467)) ;
    mux21 L1_1_L2_0_G1_MINI_ALU_ix484 (.Y (L1_1_L2_0_G1_MINI_ALU_nx483), .A0 (
          nx2612), .A1 (L1_1_L2_0_G1_MINI_ALU_BoothP_11), .S0 (
          L1_1_L2_0_G1_MINI_ALU_nx479)) ;
    inv01 ix2611 (.Y (nx2612), .A (L1_1_L2_0_G1_MINI_ALU_nx475)) ;
    mux21 L1_1_L2_0_G1_MINI_ALU_ix492 (.Y (L1_1_L2_0_G1_MINI_ALU_nx491), .A0 (
          nx2614), .A1 (L1_1_L2_0_G1_MINI_ALU_BoothP_12), .S0 (
          L1_1_L2_0_G1_MINI_ALU_nx487)) ;
    inv01 ix2613 (.Y (nx2614), .A (L1_1_L2_0_G1_MINI_ALU_nx483)) ;
    mux21 L1_1_L2_0_G1_MINI_ALU_ix500 (.Y (L1_1_L2_0_G1_MINI_ALU_nx499), .A0 (
          nx2616), .A1 (L1_1_L2_0_G1_MINI_ALU_BoothP_13), .S0 (
          L1_1_L2_0_G1_MINI_ALU_nx495)) ;
    inv01 ix2615 (.Y (nx2616), .A (L1_1_L2_0_G1_MINI_ALU_nx491)) ;
    mux21 L1_1_L2_0_G1_MINI_ALU_ix508 (.Y (L1_1_L2_0_G1_MINI_ALU_nx507), .A0 (
          nx2618), .A1 (L1_1_L2_0_G1_MINI_ALU_BoothP_14), .S0 (
          L1_1_L2_0_G1_MINI_ALU_nx503)) ;
    inv01 ix2617 (.Y (nx2618), .A (L1_1_L2_0_G1_MINI_ALU_nx499)) ;
    mux21 L1_1_L2_0_G1_MINI_ALU_ix516 (.Y (L1_1_L2_0_G1_MINI_ALU_nx515), .A0 (
          nx2620), .A1 (L1_1_L2_0_G1_MINI_ALU_BoothP_15), .S0 (
          L1_1_L2_0_G1_MINI_ALU_nx511)) ;
    inv01 ix2619 (.Y (nx2620), .A (L1_1_L2_0_G1_MINI_ALU_nx507)) ;
    mux21 L1_1_L2_0_G1_MINI_ALU_ix161 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_1), .A0 (nx2622), .A1 (
          L1_1_L2_0_G1_MINI_ALU_nx379), .S0 (nx7798)) ;
    inv01 ix2621 (.Y (nx2622), .A (L1_1_L2_0_G1_MINI_ALU_BoothP_1)) ;
    mux21 L1_1_L2_0_G1_MINI_ALU_ix181 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_2), .A0 (
          L1_1_L2_0_G1_MINI_ALU_nx387), .A1 (L1_1_L2_0_G1_MINI_ALU_nx389), .S0 (
          nx7798)) ;
    mux21 L1_1_L2_0_G1_MINI_ALU_ix201 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_3), .A0 (
          L1_1_L2_0_G1_MINI_ALU_nx399), .A1 (L1_1_L2_0_G1_MINI_ALU_nx401), .S0 (
          nx7798)) ;
    mux21 L1_1_L2_0_G1_MINI_ALU_ix221 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_4), .A0 (
          L1_1_L2_0_G1_MINI_ALU_nx409), .A1 (L1_1_L2_0_G1_MINI_ALU_nx411), .S0 (
          nx7798)) ;
    mux21 L1_1_L2_0_G1_MINI_ALU_ix241 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_5), .A0 (
          L1_1_L2_0_G1_MINI_ALU_nx419), .A1 (L1_1_L2_0_G1_MINI_ALU_nx421), .S0 (
          nx7798)) ;
    mux21 L1_1_L2_0_G1_MINI_ALU_ix261 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_6), .A0 (
          L1_1_L2_0_G1_MINI_ALU_nx429), .A1 (L1_1_L2_0_G1_MINI_ALU_nx431), .S0 (
          nx7798)) ;
    mux21 L1_1_L2_0_G1_MINI_ALU_ix281 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_7), .A0 (
          L1_1_L2_0_G1_MINI_ALU_nx439), .A1 (L1_1_L2_0_G1_MINI_ALU_nx441), .S0 (
          nx7798)) ;
    mux21 L1_1_L2_0_G1_MINI_ALU_ix301 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_8), .A0 (
          L1_1_L2_0_G1_MINI_ALU_nx449), .A1 (L1_1_L2_0_G1_MINI_ALU_nx451), .S0 (
          nx7800)) ;
    mux21 L1_1_L2_0_G1_MINI_ALU_ix321 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_9), .A0 (
          L1_1_L2_0_G1_MINI_ALU_nx469), .A1 (nx2624), .S0 (nx7800)) ;
    inv01 ix2623 (.Y (nx2624), .A (L1_1_L2_0_G1_MINI_ALU_nx316)) ;
    mux21 L1_1_L2_0_G1_MINI_ALU_ix341 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_10), .A0 (
          L1_1_L2_0_G1_MINI_ALU_nx477), .A1 (nx2626), .S0 (nx7800)) ;
    inv01 ix2625 (.Y (nx2626), .A (L1_1_L2_0_G1_MINI_ALU_nx336)) ;
    mux21 L1_1_L2_0_G1_MINI_ALU_ix361 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_11), .A0 (
          L1_1_L2_0_G1_MINI_ALU_nx485), .A1 (nx2628), .S0 (nx7800)) ;
    inv01 ix2627 (.Y (nx2628), .A (L1_1_L2_0_G1_MINI_ALU_nx356)) ;
    mux21 L1_1_L2_0_G1_MINI_ALU_ix381 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_12), .A0 (
          L1_1_L2_0_G1_MINI_ALU_nx493), .A1 (nx2630), .S0 (nx7800)) ;
    inv01 ix2629 (.Y (nx2630), .A (L1_1_L2_0_G1_MINI_ALU_nx376)) ;
    mux21 L1_1_L2_0_G1_MINI_ALU_ix401 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_13), .A0 (
          L1_1_L2_0_G1_MINI_ALU_nx501), .A1 (nx2632), .S0 (nx7800)) ;
    inv01 ix2631 (.Y (nx2632), .A (L1_1_L2_0_G1_MINI_ALU_nx396)) ;
    mux21 L1_1_L2_0_G1_MINI_ALU_ix421 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_14), .A0 (
          L1_1_L2_0_G1_MINI_ALU_nx509), .A1 (nx2634), .S0 (nx7800)) ;
    inv01 ix2633 (.Y (nx2634), .A (L1_1_L2_0_G1_MINI_ALU_nx416)) ;
    mux21 L1_1_L2_0_G1_MINI_ALU_ix441 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_15), .A0 (
          L1_1_L2_0_G1_MINI_ALU_nx517), .A1 (nx2636), .S0 (nx7802)) ;
    inv01 ix2635 (.Y (nx2636), .A (L1_1_L2_0_G1_MINI_ALU_nx436)) ;
    mux21 L1_1_L2_0_G1_MINI_ALU_ix461 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_16), .A0 (nx2638), .A1 (nx2640
          ), .S0 (nx7802)) ;
    inv01 ix2637 (.Y (nx2638), .A (L1_1_L2_0_G1_MINI_ALU_BoothP_16)) ;
    inv01 ix2639 (.Y (nx2640), .A (L1_1_L2_0_G1_MINI_ALU_nx456)) ;
    nor02_2x L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix319 (.Y (
             L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642), .A0 (Start), .A1 (
             CalculatingBooth_dup_1084)) ;
    nor02_2x L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix85 (.Y (
             L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_0), .A0 (nx7812), .A1 (
             nx2642)) ;
    inv01 ix2641 (.Y (nx2642), .A (L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_1)) ;
    mux21 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix125 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_1), .A0 (nx2644), .A1 (
          nx2646), .S0 (nx7812)) ;
    inv01 ix2643 (.Y (nx2644), .A (L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_2)) ;
    inv01 ix2645 (.Y (nx2646), .A (WindowDin_1__0__0)) ;
    mux21 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix133 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_2), .A0 (nx2648), .A1 (
          nx2650), .S0 (nx7812)) ;
    inv01 ix2647 (.Y (nx2648), .A (L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_3)) ;
    inv01 ix2649 (.Y (nx2650), .A (WindowDin_1__0__1)) ;
    mux21 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix141 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_3), .A0 (nx2652), .A1 (
          nx2654), .S0 (nx7812)) ;
    inv01 ix2651 (.Y (nx2652), .A (L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_4)) ;
    inv01 ix2653 (.Y (nx2654), .A (WindowDin_1__0__2)) ;
    mux21 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix149 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_4), .A0 (nx2656), .A1 (
          nx2658), .S0 (nx7812)) ;
    inv01 ix2655 (.Y (nx2656), .A (L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_5)) ;
    inv01 ix2657 (.Y (nx2658), .A (WindowDin_1__0__3)) ;
    mux21 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix157 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_5), .A0 (nx2660), .A1 (
          nx2662), .S0 (nx7812)) ;
    inv01 ix2659 (.Y (nx2660), .A (L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_6)) ;
    inv01 ix2661 (.Y (nx2662), .A (WindowDin_1__0__4)) ;
    mux21 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix165 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_6), .A0 (nx2664), .A1 (
          nx2666), .S0 (nx7812)) ;
    inv01 ix2663 (.Y (nx2664), .A (L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_7)) ;
    inv01 ix2665 (.Y (nx2666), .A (WindowDin_1__0__5)) ;
    mux21 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix173 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_7), .A0 (nx2668), .A1 (
          nx2670), .S0 (nx7814)) ;
    inv01 ix2667 (.Y (nx2668), .A (L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_8)) ;
    inv01 ix2669 (.Y (nx2670), .A (WindowDin_1__0__6)) ;
    mux21 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix181 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_8), .A0 (nx2672), .A1 (
          nx2674), .S0 (nx7814)) ;
    inv01 ix2671 (.Y (nx2672), .A (L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_9)) ;
    inv01 ix2673 (.Y (nx2674), .A (WindowDin_1__0__7)) ;
    nor02_2x L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix89 (.Y (
             L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_9), .A0 (nx7814), .A1 (
             nx2676)) ;
    inv01 ix2675 (.Y (nx2676), .A (L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_10)
          ) ;
    nor02_2x L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix93 (.Y (
             L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_10), .A0 (nx7814), .A1 (
             nx2678)) ;
    inv01 ix2677 (.Y (nx2678), .A (L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_11)
          ) ;
    nor02_2x L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix97 (.Y (
             L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_11), .A0 (nx7814), .A1 (
             nx2680)) ;
    inv01 ix2679 (.Y (nx2680), .A (L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_12)
          ) ;
    nor02_2x L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix101 (.Y (
             L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_12), .A0 (nx7814), .A1 (
             nx2682)) ;
    inv01 ix2681 (.Y (nx2682), .A (L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_13)
          ) ;
    nor02_2x L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix105 (.Y (
             L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_13), .A0 (nx7814), .A1 (
             nx2684)) ;
    inv01 ix2683 (.Y (nx2684), .A (L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_14)
          ) ;
    nor02_2x L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix109 (.Y (
             L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_14), .A0 (nx7816), .A1 (
             nx2686)) ;
    inv01 ix2685 (.Y (nx2686), .A (L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_15)
          ) ;
    nor02_2x L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix113 (.Y (
             L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_15), .A0 (nx7816), .A1 (
             nx2688)) ;
    inv01 ix2687 (.Y (nx2688), .A (L1_1_L2_0_G1_MINI_ALU_BoothPBeforeShift_16)
          ) ;
    nor02_2x L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix117 (.Y (
             L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_16), .A0 (nx7816), .A1 (
             nx2688)) ;
    mux21 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix189 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BoothOperand_0), .A0 (nx2690), .A1 (nx2692), .S0 (
          nx7804)) ;
    inv01 ix2689 (.Y (nx2690), .A (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_0)) ;
    inv01 ix2691 (.Y (nx2692), .A (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_0)) ;
    mux21 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix197 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BoothOperand_1), .A0 (nx2694), .A1 (nx2696), .S0 (
          nx7804)) ;
    inv01 ix2693 (.Y (nx2694), .A (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_1)) ;
    inv01 ix2695 (.Y (nx2696), .A (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_1)) ;
    mux21 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix205 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BoothOperand_2), .A0 (nx2698), .A1 (nx2700), .S0 (
          nx7804)) ;
    inv01 ix2697 (.Y (nx2698), .A (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_2)) ;
    inv01 ix2699 (.Y (nx2700), .A (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_2)) ;
    mux21 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix213 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BoothOperand_3), .A0 (nx2702), .A1 (nx2704), .S0 (
          nx7804)) ;
    inv01 ix2701 (.Y (nx2702), .A (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_3)) ;
    inv01 ix2703 (.Y (nx2704), .A (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_3)) ;
    mux21 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix221 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BoothOperand_4), .A0 (nx2706), .A1 (nx2708), .S0 (
          nx7804)) ;
    inv01 ix2705 (.Y (nx2706), .A (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_4)) ;
    inv01 ix2707 (.Y (nx2708), .A (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_4)) ;
    mux21 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix229 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BoothOperand_5), .A0 (nx2710), .A1 (nx2712), .S0 (
          nx7806)) ;
    inv01 ix2709 (.Y (nx2710), .A (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_5)) ;
    inv01 ix2711 (.Y (nx2712), .A (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_5)) ;
    mux21 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix237 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BoothOperand_6), .A0 (nx2714), .A1 (nx2716), .S0 (
          nx7806)) ;
    inv01 ix2713 (.Y (nx2714), .A (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_6)) ;
    inv01 ix2715 (.Y (nx2716), .A (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_6)) ;
    mux21 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix245 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BoothOperand_7), .A0 (nx2718), .A1 (nx2720), .S0 (
          nx7806)) ;
    inv01 ix2717 (.Y (nx2718), .A (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_7)) ;
    inv01 ix2719 (.Y (nx2720), .A (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_7)) ;
    mux21 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix253 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BoothOperand_8), .A0 (nx2722), .A1 (nx2724), .S0 (
          nx7806)) ;
    inv01 ix2721 (.Y (nx2722), .A (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_8)) ;
    inv01 ix2723 (.Y (nx2724), .A (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_8)) ;
    mux21 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix261 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BoothOperand_9), .A0 (nx2726), .A1 (nx2728), .S0 (
          nx7806)) ;
    inv01 ix2725 (.Y (nx2726), .A (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_9)) ;
    inv01 ix2727 (.Y (nx2728), .A (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_9)) ;
    mux21 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix269 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BoothOperand_10), .A0 (nx2730), .A1 (nx2732), .S0 (
          nx7806)) ;
    inv01 ix2729 (.Y (nx2730), .A (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_10)) ;
    inv01 ix2731 (.Y (nx2732), .A (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_10)) ;
    mux21 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix277 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BoothOperand_11), .A0 (nx2734), .A1 (nx2736), .S0 (
          nx7806)) ;
    inv01 ix2733 (.Y (nx2734), .A (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_11)) ;
    inv01 ix2735 (.Y (nx2736), .A (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_11)) ;
    mux21 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix285 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BoothOperand_12), .A0 (nx2738), .A1 (nx2740), .S0 (
          nx7808)) ;
    inv01 ix2737 (.Y (nx2738), .A (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_12)) ;
    inv01 ix2739 (.Y (nx2740), .A (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_12)) ;
    mux21 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix293 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BoothOperand_13), .A0 (nx2742), .A1 (nx2744), .S0 (
          nx7808)) ;
    inv01 ix2741 (.Y (nx2742), .A (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_13)) ;
    inv01 ix2743 (.Y (nx2744), .A (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_13)) ;
    mux21 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix301 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BoothOperand_14), .A0 (nx2746), .A1 (nx2748), .S0 (
          nx7808)) ;
    inv01 ix2745 (.Y (nx2746), .A (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_14)) ;
    inv01 ix2747 (.Y (nx2748), .A (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_14)) ;
    mux21 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix309 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BoothOperand_15), .A0 (nx2750), .A1 (nx2752), .S0 (
          nx7808)) ;
    inv01 ix2749 (.Y (nx2750), .A (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_15)) ;
    inv01 ix2751 (.Y (nx2752), .A (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_15)) ;
    mux21 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix317 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BoothOperand_16), .A0 (nx2754), .A1 (nx2756), .S0 (
          nx7808)) ;
    inv01 ix2753 (.Y (nx2754), .A (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_16)) ;
    inv01 ix2755 (.Y (nx2756), .A (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_16)) ;
    xnor2 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix321 (.Y (
          L1_1_L2_0_G1_MINI_ALU_AddPToBoothOperand), .A0 (nx7808), .A1 (nx2622)
          ) ;
    oai32 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix393 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .A0 (nx8626), .A1 (
          RST), .A2 (nx7818), .B0 (nx2692), .B1 (nx2760)) ;
    oai32 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix403 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .A0 (nx8626), .A1 (
          RST), .A2 (nx7818), .B0 (nx2696), .B1 (nx2760)) ;
    oai32 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix413 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .A0 (nx8626), .A1 (
          RST), .A2 (nx7818), .B0 (nx2700), .B1 (nx2760)) ;
    oai32 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix423 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .A0 (nx8626), .A1 (
          RST), .A2 (nx7818), .B0 (nx2704), .B1 (nx2760)) ;
    oai32 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix433 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .A0 (nx8626), .A1 (
          RST), .A2 (nx7818), .B0 (nx2708), .B1 (nx2760)) ;
    oai32 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix443 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .A0 (nx8626), .A1 (
          RST), .A2 (nx7818), .B0 (nx2712), .B1 (nx2760)) ;
    oai32 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix453 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .A0 (nx8626), .A1 (
          RST), .A2 (nx7820), .B0 (nx2716), .B1 (nx2760)) ;
    oai32 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix463 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .A0 (nx8628), .A1 (
          RST), .A2 (nx7820), .B0 (nx2720), .B1 (nx2762)) ;
    oai32 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix473 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .A0 (nx8628), .A1 (
          RST), .A2 (nx7820), .B0 (nx2724), .B1 (nx2762)) ;
    oai32 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix483 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .A0 (nx2764), .A1 (
          RST), .A2 (nx7820), .B0 (nx2728), .B1 (nx2762)) ;
    inv01 ix2763 (.Y (nx2764), .A (FilterDin_1__0__0)) ;
    oai32 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix493 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .A0 (nx2766), .A1 (
          RST), .A2 (nx7820), .B0 (nx2732), .B1 (nx2762)) ;
    inv01 ix2765 (.Y (nx2766), .A (FilterDin_1__0__1)) ;
    oai32 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix503 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .A0 (nx2768), .A1 (
          RST), .A2 (nx7820), .B0 (nx2736), .B1 (nx2762)) ;
    inv01 ix2767 (.Y (nx2768), .A (FilterDin_1__0__2)) ;
    oai32 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix513 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .A0 (nx2770), .A1 (
          RST), .A2 (nx7820), .B0 (nx2740), .B1 (nx2762)) ;
    inv01 ix2769 (.Y (nx2770), .A (FilterDin_1__0__3)) ;
    oai32 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix523 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .A0 (nx2772), .A1 (
          RST), .A2 (nx7822), .B0 (nx2744), .B1 (nx2762)) ;
    inv01 ix2771 (.Y (nx2772), .A (FilterDin_1__0__4)) ;
    oai32 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix533 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .A0 (nx2774), .A1 (
          RST), .A2 (nx7822), .B0 (nx2748), .B1 (nx2776)) ;
    inv01 ix2773 (.Y (nx2774), .A (FilterDin_1__0__5)) ;
    inv01 ix2775 (.Y (nx2776), .A (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566)) ;
    oai32 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix543 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .A0 (nx2778), .A1 (
          RST), .A2 (nx7822), .B0 (nx2752), .B1 (nx2776)) ;
    inv01 ix2777 (.Y (nx2778), .A (FilterDin_1__0__6)) ;
    oai32 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix553 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .A0 (nx2780), .A1 (
          RST), .A2 (nx7822), .B0 (nx2756), .B1 (nx2776)) ;
    inv01 ix2779 (.Y (nx2780), .A (FilterDin_1__0__7)) ;
    nand02_2x L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix633 (.Y (nx2760), .A0 (
              nx7584), .A1 (nx7822)) ;
    nand02_2x L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix635 (.Y (nx2762), .A0 (
              nx7584), .A1 (nx7822)) ;
    oai32 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix393 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .A0 (nx8628), .A1 (
          RST), .A2 (nx7824), .B0 (nx2690), .B1 (nx2782)) ;
    oai32 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix403 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .A0 (nx8628), .A1 (
          RST), .A2 (nx7824), .B0 (nx2694), .B1 (nx2782)) ;
    oai32 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix413 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .A0 (nx8628), .A1 (
          RST), .A2 (nx7824), .B0 (nx2698), .B1 (nx2782)) ;
    oai32 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix423 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .A0 (nx8628), .A1 (
          RST), .A2 (nx7824), .B0 (nx2702), .B1 (nx2782)) ;
    oai32 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix433 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .A0 (nx8628), .A1 (
          RST), .A2 (nx7824), .B0 (nx2706), .B1 (nx2782)) ;
    oai32 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix443 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .A0 (nx8630), .A1 (
          RST), .A2 (nx7824), .B0 (nx2710), .B1 (nx2782)) ;
    oai32 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix453 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .A0 (nx8630), .A1 (
          RST), .A2 (nx7826), .B0 (nx2714), .B1 (nx2782)) ;
    oai32 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix463 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .A0 (nx8630), .A1 (
          RST), .A2 (nx7826), .B0 (nx2718), .B1 (nx2784)) ;
    oai32 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix473 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .A0 (nx8630), .A1 (
          RST), .A2 (nx7826), .B0 (nx2722), .B1 (nx2784)) ;
    oai32 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix483 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .A0 (nx2764), .A1 (
          RST), .A2 (nx7826), .B0 (nx2726), .B1 (nx2784)) ;
    oai32 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix493 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .A0 (nx2786), .A1 (
          RST), .A2 (nx7826), .B0 (nx2730), .B1 (nx2784)) ;
    inv01 ix2785 (.Y (nx2786), .A (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_10)) ;
    oai32 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix503 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .A0 (nx2788), .A1 (
          RST), .A2 (nx7826), .B0 (nx2734), .B1 (nx2784)) ;
    inv01 ix2787 (.Y (nx2788), .A (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_11)) ;
    oai32 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix513 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .A0 (nx2790), .A1 (
          RST), .A2 (nx7826), .B0 (nx2738), .B1 (nx2784)) ;
    inv01 ix2789 (.Y (nx2790), .A (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_12)) ;
    oai32 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix523 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .A0 (nx2792), .A1 (
          RST), .A2 (nx7828), .B0 (nx2742), .B1 (nx2784)) ;
    inv01 ix2791 (.Y (nx2792), .A (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_13)) ;
    oai32 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix533 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .A0 (nx2794), .A1 (
          RST), .A2 (nx7828), .B0 (nx2746), .B1 (nx2796)) ;
    inv01 ix2793 (.Y (nx2794), .A (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_14)) ;
    inv01 ix2795 (.Y (nx2796), .A (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566)) ;
    oai32 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix543 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .A0 (nx2798), .A1 (
          RST), .A2 (nx7828), .B0 (nx2750), .B1 (nx2796)) ;
    inv01 ix2797 (.Y (nx2798), .A (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_15)) ;
    oai32 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix553 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .A0 (nx2800), .A1 (
          RST), .A2 (nx7828), .B0 (nx2754), .B1 (nx2796)) ;
    inv01 ix2799 (.Y (nx2800), .A (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_16)) ;
    nand02_2x L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix633 (.Y (nx2782), .A0 (
              nx7584), .A1 (nx7828)) ;
    nand02_2x L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix635 (.Y (nx2784), .A0 (
              nx7584), .A1 (nx7828)) ;
    oai32 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix393 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .A0 (nx2802), .A1 (
          RST), .A2 (nx7830), .B0 (L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx384), .B1 (
          nx2804)) ;
    inv01 ix2801 (.Y (nx2802), .A (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_0)) ;
    oai32 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix403 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .A0 (nx2806), .A1 (
          RST), .A2 (nx7830), .B0 (nx2622), .B1 (nx2804)) ;
    inv01 ix2805 (.Y (nx2806), .A (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_1)) ;
    oai32 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix413 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .A0 (nx2808), .A1 (
          RST), .A2 (nx7830), .B0 (L1_1_L2_0_G1_MINI_ALU_nx387), .B1 (nx2804)) ;
    inv01 ix2807 (.Y (nx2808), .A (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_2)) ;
    oai32 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix423 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .A0 (nx2810), .A1 (
          RST), .A2 (nx7830), .B0 (L1_1_L2_0_G1_MINI_ALU_nx399), .B1 (nx2804)) ;
    inv01 ix2809 (.Y (nx2810), .A (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_3)) ;
    oai32 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix433 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .A0 (nx2812), .A1 (
          RST), .A2 (nx7830), .B0 (L1_1_L2_0_G1_MINI_ALU_nx409), .B1 (nx2804)) ;
    inv01 ix2811 (.Y (nx2812), .A (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_4)) ;
    oai32 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix443 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .A0 (nx2814), .A1 (
          RST), .A2 (nx7830), .B0 (L1_1_L2_0_G1_MINI_ALU_nx419), .B1 (nx2804)) ;
    inv01 ix2813 (.Y (nx2814), .A (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_5)) ;
    oai32 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix453 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .A0 (nx2816), .A1 (
          RST), .A2 (nx7830), .B0 (L1_1_L2_0_G1_MINI_ALU_nx429), .B1 (nx2804)) ;
    inv01 ix2815 (.Y (nx2816), .A (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_6)) ;
    oai32 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix463 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .A0 (nx2818), .A1 (
          RST), .A2 (nx7832), .B0 (L1_1_L2_0_G1_MINI_ALU_nx439), .B1 (nx2820)) ;
    inv01 ix2817 (.Y (nx2818), .A (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_7)) ;
    oai32 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix473 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .A0 (nx2822), .A1 (
          RST), .A2 (nx7832), .B0 (L1_1_L2_0_G1_MINI_ALU_nx449), .B1 (nx2820)) ;
    inv01 ix2821 (.Y (nx2822), .A (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_8)) ;
    oai32 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix483 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .A0 (nx2824), .A1 (
          RST), .A2 (nx7832), .B0 (L1_1_L2_0_G1_MINI_ALU_nx469), .B1 (nx2820)) ;
    inv01 ix2823 (.Y (nx2824), .A (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_9)) ;
    oai32 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix493 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .A0 (nx2826), .A1 (
          RST), .A2 (nx7832), .B0 (L1_1_L2_0_G1_MINI_ALU_nx477), .B1 (nx2820)) ;
    inv01 ix2825 (.Y (nx2826), .A (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_10)) ;
    oai32 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix503 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .A0 (nx2828), .A1 (
          RST), .A2 (nx7832), .B0 (L1_1_L2_0_G1_MINI_ALU_nx485), .B1 (nx2820)) ;
    inv01 ix2827 (.Y (nx2828), .A (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_11)) ;
    oai32 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix513 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .A0 (nx2830), .A1 (
          RST), .A2 (nx7832), .B0 (L1_1_L2_0_G1_MINI_ALU_nx493), .B1 (nx2820)) ;
    inv01 ix2829 (.Y (nx2830), .A (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_12)) ;
    oai32 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix523 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .A0 (nx2832), .A1 (
          RST), .A2 (nx7832), .B0 (L1_1_L2_0_G1_MINI_ALU_nx501), .B1 (nx2820)) ;
    inv01 ix2831 (.Y (nx2832), .A (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_13)) ;
    oai32 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix533 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .A0 (nx2834), .A1 (
          RST), .A2 (nx7834), .B0 (L1_1_L2_0_G1_MINI_ALU_nx509), .B1 (nx2836)) ;
    inv01 ix2833 (.Y (nx2834), .A (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_14)) ;
    inv01 ix2835 (.Y (nx2836), .A (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566)) ;
    oai32 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix543 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .A0 (nx2838), .A1 (
          RST), .A2 (nx7834), .B0 (L1_1_L2_0_G1_MINI_ALU_nx517), .B1 (nx2836)) ;
    inv01 ix2837 (.Y (nx2838), .A (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_15)) ;
    oai32 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix553 (.Y (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .A0 (nx2840), .A1 (
          RST), .A2 (nx7834), .B0 (nx2638), .B1 (nx2836)) ;
    inv01 ix2839 (.Y (nx2840), .A (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_16)) ;
    nand02_2x L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix633 (.Y (nx2804), .A0 (
              nx7584), .A1 (nx7834)) ;
    nand02_2x L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix635 (.Y (nx2820), .A0 (
              nx7586), .A1 (nx7834)) ;
    mux21 L1_1_L2_1_G1_MINI_ALU_ix404 (.Y (L1_1_L2_1_G1_MINI_ALU_nx403), .A0 (
          nx2842), .A1 (L1_1_L2_1_G1_MINI_ALU_BoothP_2), .S0 (
          L1_1_L2_1_G1_MINI_ALU_nx395)) ;
    inv01 ix2841 (.Y (nx2842), .A (L1_1_L2_1_G1_MINI_ALU_nx391)) ;
    mux21 L1_1_L2_1_G1_MINI_ALU_ix414 (.Y (L1_1_L2_1_G1_MINI_ALU_nx413), .A0 (
          nx2844), .A1 (L1_1_L2_1_G1_MINI_ALU_BoothP_3), .S0 (
          L1_1_L2_1_G1_MINI_ALU_nx405)) ;
    inv01 ix2843 (.Y (nx2844), .A (L1_1_L2_1_G1_MINI_ALU_nx403)) ;
    mux21 L1_1_L2_1_G1_MINI_ALU_ix424 (.Y (L1_1_L2_1_G1_MINI_ALU_nx423), .A0 (
          nx2846), .A1 (L1_1_L2_1_G1_MINI_ALU_BoothP_4), .S0 (
          L1_1_L2_1_G1_MINI_ALU_nx415)) ;
    inv01 ix2845 (.Y (nx2846), .A (L1_1_L2_1_G1_MINI_ALU_nx413)) ;
    mux21 L1_1_L2_1_G1_MINI_ALU_ix434 (.Y (L1_1_L2_1_G1_MINI_ALU_nx433), .A0 (
          nx2848), .A1 (L1_1_L2_1_G1_MINI_ALU_BoothP_5), .S0 (
          L1_1_L2_1_G1_MINI_ALU_nx425)) ;
    inv01 ix2847 (.Y (nx2848), .A (L1_1_L2_1_G1_MINI_ALU_nx423)) ;
    mux21 L1_1_L2_1_G1_MINI_ALU_ix444 (.Y (L1_1_L2_1_G1_MINI_ALU_nx443), .A0 (
          nx2850), .A1 (L1_1_L2_1_G1_MINI_ALU_BoothP_6), .S0 (
          L1_1_L2_1_G1_MINI_ALU_nx435)) ;
    inv01 ix2849 (.Y (nx2850), .A (L1_1_L2_1_G1_MINI_ALU_nx433)) ;
    mux21 L1_1_L2_1_G1_MINI_ALU_ix454 (.Y (L1_1_L2_1_G1_MINI_ALU_nx453), .A0 (
          nx2852), .A1 (L1_1_L2_1_G1_MINI_ALU_BoothP_7), .S0 (
          L1_1_L2_1_G1_MINI_ALU_nx445)) ;
    inv01 ix2851 (.Y (nx2852), .A (L1_1_L2_1_G1_MINI_ALU_nx443)) ;
    mux21 L1_1_L2_1_G1_MINI_ALU_ix462 (.Y (L1_1_L2_1_G1_MINI_ALU_nx461), .A0 (
          nx2854), .A1 (L1_1_L2_1_G1_MINI_ALU_BoothP_8), .S0 (
          L1_1_L2_1_G1_MINI_ALU_nx455)) ;
    inv01 ix2853 (.Y (nx2854), .A (L1_1_L2_1_G1_MINI_ALU_nx453)) ;
    mux21 L1_1_L2_1_G1_MINI_ALU_ix468 (.Y (L1_1_L2_1_G1_MINI_ALU_nx467), .A0 (
          nx2856), .A1 (L1_1_L2_1_G1_MINI_ALU_BoothP_9), .S0 (
          L1_1_L2_1_G1_MINI_ALU_nx463)) ;
    inv01 ix2855 (.Y (nx2856), .A (L1_1_L2_1_G1_MINI_ALU_nx461)) ;
    mux21 L1_1_L2_1_G1_MINI_ALU_ix476 (.Y (L1_1_L2_1_G1_MINI_ALU_nx475), .A0 (
          nx2858), .A1 (L1_1_L2_1_G1_MINI_ALU_BoothP_10), .S0 (
          L1_1_L2_1_G1_MINI_ALU_nx471)) ;
    inv01 ix2857 (.Y (nx2858), .A (L1_1_L2_1_G1_MINI_ALU_nx467)) ;
    mux21 L1_1_L2_1_G1_MINI_ALU_ix484 (.Y (L1_1_L2_1_G1_MINI_ALU_nx483), .A0 (
          nx2860), .A1 (L1_1_L2_1_G1_MINI_ALU_BoothP_11), .S0 (
          L1_1_L2_1_G1_MINI_ALU_nx479)) ;
    inv01 ix2859 (.Y (nx2860), .A (L1_1_L2_1_G1_MINI_ALU_nx475)) ;
    mux21 L1_1_L2_1_G1_MINI_ALU_ix492 (.Y (L1_1_L2_1_G1_MINI_ALU_nx491), .A0 (
          nx2862), .A1 (L1_1_L2_1_G1_MINI_ALU_BoothP_12), .S0 (
          L1_1_L2_1_G1_MINI_ALU_nx487)) ;
    inv01 ix2861 (.Y (nx2862), .A (L1_1_L2_1_G1_MINI_ALU_nx483)) ;
    mux21 L1_1_L2_1_G1_MINI_ALU_ix500 (.Y (L1_1_L2_1_G1_MINI_ALU_nx499), .A0 (
          nx2864), .A1 (L1_1_L2_1_G1_MINI_ALU_BoothP_13), .S0 (
          L1_1_L2_1_G1_MINI_ALU_nx495)) ;
    inv01 ix2863 (.Y (nx2864), .A (L1_1_L2_1_G1_MINI_ALU_nx491)) ;
    mux21 L1_1_L2_1_G1_MINI_ALU_ix508 (.Y (L1_1_L2_1_G1_MINI_ALU_nx507), .A0 (
          nx2866), .A1 (L1_1_L2_1_G1_MINI_ALU_BoothP_14), .S0 (
          L1_1_L2_1_G1_MINI_ALU_nx503)) ;
    inv01 ix2865 (.Y (nx2866), .A (L1_1_L2_1_G1_MINI_ALU_nx499)) ;
    mux21 L1_1_L2_1_G1_MINI_ALU_ix516 (.Y (L1_1_L2_1_G1_MINI_ALU_nx515), .A0 (
          nx2868), .A1 (L1_1_L2_1_G1_MINI_ALU_BoothP_15), .S0 (
          L1_1_L2_1_G1_MINI_ALU_nx511)) ;
    inv01 ix2867 (.Y (nx2868), .A (L1_1_L2_1_G1_MINI_ALU_nx507)) ;
    mux21 L1_1_L2_1_G1_MINI_ALU_ix161 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_1), .A0 (nx2870), .A1 (
          L1_1_L2_1_G1_MINI_ALU_nx379), .S0 (nx7838)) ;
    inv01 ix2869 (.Y (nx2870), .A (L1_1_L2_1_G1_MINI_ALU_BoothP_1)) ;
    mux21 L1_1_L2_1_G1_MINI_ALU_ix181 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_2), .A0 (
          L1_1_L2_1_G1_MINI_ALU_nx387), .A1 (L1_1_L2_1_G1_MINI_ALU_nx389), .S0 (
          nx7838)) ;
    mux21 L1_1_L2_1_G1_MINI_ALU_ix201 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_3), .A0 (
          L1_1_L2_1_G1_MINI_ALU_nx399), .A1 (L1_1_L2_1_G1_MINI_ALU_nx401), .S0 (
          nx7838)) ;
    mux21 L1_1_L2_1_G1_MINI_ALU_ix221 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_4), .A0 (
          L1_1_L2_1_G1_MINI_ALU_nx409), .A1 (L1_1_L2_1_G1_MINI_ALU_nx411), .S0 (
          nx7838)) ;
    mux21 L1_1_L2_1_G1_MINI_ALU_ix241 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_5), .A0 (
          L1_1_L2_1_G1_MINI_ALU_nx419), .A1 (L1_1_L2_1_G1_MINI_ALU_nx421), .S0 (
          nx7838)) ;
    mux21 L1_1_L2_1_G1_MINI_ALU_ix261 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_6), .A0 (
          L1_1_L2_1_G1_MINI_ALU_nx429), .A1 (L1_1_L2_1_G1_MINI_ALU_nx431), .S0 (
          nx7838)) ;
    mux21 L1_1_L2_1_G1_MINI_ALU_ix281 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_7), .A0 (
          L1_1_L2_1_G1_MINI_ALU_nx439), .A1 (L1_1_L2_1_G1_MINI_ALU_nx441), .S0 (
          nx7838)) ;
    mux21 L1_1_L2_1_G1_MINI_ALU_ix301 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_8), .A0 (
          L1_1_L2_1_G1_MINI_ALU_nx449), .A1 (L1_1_L2_1_G1_MINI_ALU_nx451), .S0 (
          nx7840)) ;
    mux21 L1_1_L2_1_G1_MINI_ALU_ix321 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_9), .A0 (
          L1_1_L2_1_G1_MINI_ALU_nx469), .A1 (nx2872), .S0 (nx7840)) ;
    inv01 ix2871 (.Y (nx2872), .A (L1_1_L2_1_G1_MINI_ALU_nx316)) ;
    mux21 L1_1_L2_1_G1_MINI_ALU_ix341 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_10), .A0 (
          L1_1_L2_1_G1_MINI_ALU_nx477), .A1 (nx2874), .S0 (nx7840)) ;
    inv01 ix2873 (.Y (nx2874), .A (L1_1_L2_1_G1_MINI_ALU_nx336)) ;
    mux21 L1_1_L2_1_G1_MINI_ALU_ix361 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_11), .A0 (
          L1_1_L2_1_G1_MINI_ALU_nx485), .A1 (nx2876), .S0 (nx7840)) ;
    inv01 ix2875 (.Y (nx2876), .A (L1_1_L2_1_G1_MINI_ALU_nx356)) ;
    mux21 L1_1_L2_1_G1_MINI_ALU_ix381 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_12), .A0 (
          L1_1_L2_1_G1_MINI_ALU_nx493), .A1 (nx2878), .S0 (nx7840)) ;
    inv01 ix2877 (.Y (nx2878), .A (L1_1_L2_1_G1_MINI_ALU_nx376)) ;
    mux21 L1_1_L2_1_G1_MINI_ALU_ix401 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_13), .A0 (
          L1_1_L2_1_G1_MINI_ALU_nx501), .A1 (nx2880), .S0 (nx7840)) ;
    inv01 ix2879 (.Y (nx2880), .A (L1_1_L2_1_G1_MINI_ALU_nx396)) ;
    mux21 L1_1_L2_1_G1_MINI_ALU_ix421 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_14), .A0 (
          L1_1_L2_1_G1_MINI_ALU_nx509), .A1 (nx2882), .S0 (nx7840)) ;
    inv01 ix2881 (.Y (nx2882), .A (L1_1_L2_1_G1_MINI_ALU_nx416)) ;
    mux21 L1_1_L2_1_G1_MINI_ALU_ix441 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_15), .A0 (
          L1_1_L2_1_G1_MINI_ALU_nx517), .A1 (nx2884), .S0 (nx7842)) ;
    inv01 ix2883 (.Y (nx2884), .A (L1_1_L2_1_G1_MINI_ALU_nx436)) ;
    mux21 L1_1_L2_1_G1_MINI_ALU_ix461 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_16), .A0 (nx2886), .A1 (nx2888
          ), .S0 (nx7842)) ;
    inv01 ix2885 (.Y (nx2886), .A (L1_1_L2_1_G1_MINI_ALU_BoothP_16)) ;
    inv01 ix2887 (.Y (nx2888), .A (L1_1_L2_1_G1_MINI_ALU_nx456)) ;
    nor02_2x L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix319 (.Y (
             L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642), .A0 (Start), .A1 (
             CalculatingBooth_dup_1084)) ;
    nor02_2x L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix85 (.Y (
             L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_0), .A0 (nx7852), .A1 (
             nx2890)) ;
    inv01 ix2889 (.Y (nx2890), .A (L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_1)) ;
    mux21 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix125 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_1), .A0 (nx2892), .A1 (
          nx2894), .S0 (nx7852)) ;
    inv01 ix2891 (.Y (nx2892), .A (L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_2)) ;
    inv01 ix2893 (.Y (nx2894), .A (WindowDin_1__1__0)) ;
    mux21 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix133 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_2), .A0 (nx2896), .A1 (
          nx2898), .S0 (nx7852)) ;
    inv01 ix2895 (.Y (nx2896), .A (L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_3)) ;
    inv01 ix2897 (.Y (nx2898), .A (WindowDin_1__1__1)) ;
    mux21 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix141 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_3), .A0 (nx2900), .A1 (
          nx2902), .S0 (nx7852)) ;
    inv01 ix2899 (.Y (nx2900), .A (L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_4)) ;
    inv01 ix2901 (.Y (nx2902), .A (WindowDin_1__1__2)) ;
    mux21 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix149 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_4), .A0 (nx2904), .A1 (
          nx2906), .S0 (nx7852)) ;
    inv01 ix2903 (.Y (nx2904), .A (L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_5)) ;
    inv01 ix2905 (.Y (nx2906), .A (WindowDin_1__1__3)) ;
    mux21 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix157 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_5), .A0 (nx2908), .A1 (
          nx2910), .S0 (nx7852)) ;
    inv01 ix2907 (.Y (nx2908), .A (L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_6)) ;
    inv01 ix2909 (.Y (nx2910), .A (WindowDin_1__1__4)) ;
    mux21 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix165 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_6), .A0 (nx2912), .A1 (
          nx2914), .S0 (nx7852)) ;
    inv01 ix2911 (.Y (nx2912), .A (L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_7)) ;
    inv01 ix2913 (.Y (nx2914), .A (WindowDin_1__1__5)) ;
    mux21 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix173 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_7), .A0 (nx2916), .A1 (
          nx2918), .S0 (nx7854)) ;
    inv01 ix2915 (.Y (nx2916), .A (L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_8)) ;
    inv01 ix2917 (.Y (nx2918), .A (WindowDin_1__1__6)) ;
    mux21 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix181 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_8), .A0 (nx2920), .A1 (
          nx2922), .S0 (nx7854)) ;
    inv01 ix2919 (.Y (nx2920), .A (L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_9)) ;
    inv01 ix2921 (.Y (nx2922), .A (WindowDin_1__1__7)) ;
    nor02_2x L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix89 (.Y (
             L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_9), .A0 (nx7854), .A1 (
             nx2924)) ;
    inv01 ix2923 (.Y (nx2924), .A (L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_10)
          ) ;
    nor02_2x L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix93 (.Y (
             L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_10), .A0 (nx7854), .A1 (
             nx2926)) ;
    inv01 ix2925 (.Y (nx2926), .A (L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_11)
          ) ;
    nor02_2x L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix97 (.Y (
             L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_11), .A0 (nx7854), .A1 (
             nx2928)) ;
    inv01 ix2927 (.Y (nx2928), .A (L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_12)
          ) ;
    nor02_2x L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix101 (.Y (
             L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_12), .A0 (nx7854), .A1 (
             nx2930)) ;
    inv01 ix2929 (.Y (nx2930), .A (L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_13)
          ) ;
    nor02_2x L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix105 (.Y (
             L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_13), .A0 (nx7854), .A1 (
             nx2932)) ;
    inv01 ix2931 (.Y (nx2932), .A (L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_14)
          ) ;
    nor02_2x L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix109 (.Y (
             L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_14), .A0 (nx7856), .A1 (
             nx2934)) ;
    inv01 ix2933 (.Y (nx2934), .A (L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_15)
          ) ;
    nor02_2x L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix113 (.Y (
             L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_15), .A0 (nx7856), .A1 (
             nx2936)) ;
    inv01 ix2935 (.Y (nx2936), .A (L1_1_L2_1_G1_MINI_ALU_BoothPBeforeShift_16)
          ) ;
    nor02_2x L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix117 (.Y (
             L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_16), .A0 (nx7856), .A1 (
             nx2936)) ;
    mux21 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix189 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BoothOperand_0), .A0 (nx2938), .A1 (nx2940), .S0 (
          nx7844)) ;
    inv01 ix2937 (.Y (nx2938), .A (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_0)) ;
    inv01 ix2939 (.Y (nx2940), .A (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_0)) ;
    mux21 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix197 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BoothOperand_1), .A0 (nx2942), .A1 (nx2944), .S0 (
          nx7844)) ;
    inv01 ix2941 (.Y (nx2942), .A (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_1)) ;
    inv01 ix2943 (.Y (nx2944), .A (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_1)) ;
    mux21 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix205 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BoothOperand_2), .A0 (nx2946), .A1 (nx2948), .S0 (
          nx7844)) ;
    inv01 ix2945 (.Y (nx2946), .A (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_2)) ;
    inv01 ix2947 (.Y (nx2948), .A (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_2)) ;
    mux21 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix213 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BoothOperand_3), .A0 (nx2950), .A1 (nx2952), .S0 (
          nx7844)) ;
    inv01 ix2949 (.Y (nx2950), .A (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_3)) ;
    inv01 ix2951 (.Y (nx2952), .A (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_3)) ;
    mux21 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix221 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BoothOperand_4), .A0 (nx2954), .A1 (nx2956), .S0 (
          nx7844)) ;
    inv01 ix2953 (.Y (nx2954), .A (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_4)) ;
    inv01 ix2955 (.Y (nx2956), .A (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_4)) ;
    mux21 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix229 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BoothOperand_5), .A0 (nx2958), .A1 (nx2960), .S0 (
          nx7846)) ;
    inv01 ix2957 (.Y (nx2958), .A (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_5)) ;
    inv01 ix2959 (.Y (nx2960), .A (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_5)) ;
    mux21 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix237 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BoothOperand_6), .A0 (nx2962), .A1 (nx2964), .S0 (
          nx7846)) ;
    inv01 ix2961 (.Y (nx2962), .A (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_6)) ;
    inv01 ix2963 (.Y (nx2964), .A (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_6)) ;
    mux21 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix245 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BoothOperand_7), .A0 (nx2966), .A1 (nx2968), .S0 (
          nx7846)) ;
    inv01 ix2965 (.Y (nx2966), .A (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_7)) ;
    inv01 ix2967 (.Y (nx2968), .A (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_7)) ;
    mux21 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix253 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BoothOperand_8), .A0 (nx2970), .A1 (nx2972), .S0 (
          nx7846)) ;
    inv01 ix2969 (.Y (nx2970), .A (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_8)) ;
    inv01 ix2971 (.Y (nx2972), .A (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_8)) ;
    mux21 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix261 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BoothOperand_9), .A0 (nx2974), .A1 (nx2976), .S0 (
          nx7846)) ;
    inv01 ix2973 (.Y (nx2974), .A (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_9)) ;
    inv01 ix2975 (.Y (nx2976), .A (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_9)) ;
    mux21 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix269 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BoothOperand_10), .A0 (nx2978), .A1 (nx2980), .S0 (
          nx7846)) ;
    inv01 ix2977 (.Y (nx2978), .A (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_10)) ;
    inv01 ix2979 (.Y (nx2980), .A (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_10)) ;
    mux21 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix277 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BoothOperand_11), .A0 (nx2982), .A1 (nx2984), .S0 (
          nx7846)) ;
    inv01 ix2981 (.Y (nx2982), .A (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_11)) ;
    inv01 ix2983 (.Y (nx2984), .A (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_11)) ;
    mux21 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix285 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BoothOperand_12), .A0 (nx2986), .A1 (nx2988), .S0 (
          nx7848)) ;
    inv01 ix2985 (.Y (nx2986), .A (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_12)) ;
    inv01 ix2987 (.Y (nx2988), .A (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_12)) ;
    mux21 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix293 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BoothOperand_13), .A0 (nx2990), .A1 (nx2992), .S0 (
          nx7848)) ;
    inv01 ix2989 (.Y (nx2990), .A (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_13)) ;
    inv01 ix2991 (.Y (nx2992), .A (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_13)) ;
    mux21 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix301 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BoothOperand_14), .A0 (nx2994), .A1 (nx2996), .S0 (
          nx7848)) ;
    inv01 ix2993 (.Y (nx2994), .A (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_14)) ;
    inv01 ix2995 (.Y (nx2996), .A (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_14)) ;
    mux21 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix309 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BoothOperand_15), .A0 (nx2998), .A1 (nx3000), .S0 (
          nx7848)) ;
    inv01 ix2997 (.Y (nx2998), .A (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_15)) ;
    inv01 ix2999 (.Y (nx3000), .A (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_15)) ;
    mux21 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix317 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BoothOperand_16), .A0 (nx3002), .A1 (nx3004), .S0 (
          nx7848)) ;
    inv01 ix3001 (.Y (nx3002), .A (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_16)) ;
    inv01 ix3003 (.Y (nx3004), .A (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_16)) ;
    xnor2 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix321 (.Y (
          L1_1_L2_1_G1_MINI_ALU_AddPToBoothOperand), .A0 (nx7848), .A1 (nx2870)
          ) ;
    oai32 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix393 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .A0 (nx8632), .A1 (
          RST), .A2 (nx7858), .B0 (nx2940), .B1 (nx3008)) ;
    oai32 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix403 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .A0 (nx8632), .A1 (
          RST), .A2 (nx7858), .B0 (nx2944), .B1 (nx3008)) ;
    oai32 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix413 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .A0 (nx8632), .A1 (
          RST), .A2 (nx7858), .B0 (nx2948), .B1 (nx3008)) ;
    oai32 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix423 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .A0 (nx8632), .A1 (
          RST), .A2 (nx7858), .B0 (nx2952), .B1 (nx3008)) ;
    oai32 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix433 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .A0 (nx8632), .A1 (
          RST), .A2 (nx7858), .B0 (nx2956), .B1 (nx3008)) ;
    oai32 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix443 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .A0 (nx8632), .A1 (
          RST), .A2 (nx7858), .B0 (nx2960), .B1 (nx3008)) ;
    oai32 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix453 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .A0 (nx8632), .A1 (
          RST), .A2 (nx7860), .B0 (nx2964), .B1 (nx3008)) ;
    oai32 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix463 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .A0 (nx8634), .A1 (
          RST), .A2 (nx7860), .B0 (nx2968), .B1 (nx3010)) ;
    oai32 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix473 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .A0 (nx8634), .A1 (
          RST), .A2 (nx7860), .B0 (nx2972), .B1 (nx3010)) ;
    oai32 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix483 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .A0 (nx3012), .A1 (
          RST), .A2 (nx7860), .B0 (nx2976), .B1 (nx3010)) ;
    inv01 ix3011 (.Y (nx3012), .A (FilterDin_1__1__0)) ;
    oai32 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix493 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .A0 (nx3014), .A1 (
          RST), .A2 (nx7860), .B0 (nx2980), .B1 (nx3010)) ;
    inv01 ix3013 (.Y (nx3014), .A (FilterDin_1__1__1)) ;
    oai32 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix503 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .A0 (nx3016), .A1 (
          RST), .A2 (nx7860), .B0 (nx2984), .B1 (nx3010)) ;
    inv01 ix3015 (.Y (nx3016), .A (FilterDin_1__1__2)) ;
    oai32 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix513 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .A0 (nx3018), .A1 (
          RST), .A2 (nx7860), .B0 (nx2988), .B1 (nx3010)) ;
    inv01 ix3017 (.Y (nx3018), .A (FilterDin_1__1__3)) ;
    oai32 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix523 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .A0 (nx3020), .A1 (
          RST), .A2 (nx7862), .B0 (nx2992), .B1 (nx3010)) ;
    inv01 ix3019 (.Y (nx3020), .A (FilterDin_1__1__4)) ;
    oai32 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix533 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .A0 (nx3022), .A1 (
          RST), .A2 (nx7862), .B0 (nx2996), .B1 (nx3024)) ;
    inv01 ix3021 (.Y (nx3022), .A (FilterDin_1__1__5)) ;
    inv01 ix3023 (.Y (nx3024), .A (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566)) ;
    oai32 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix543 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .A0 (nx3026), .A1 (
          RST), .A2 (nx7862), .B0 (nx3000), .B1 (nx3024)) ;
    inv01 ix3025 (.Y (nx3026), .A (FilterDin_1__1__6)) ;
    oai32 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix553 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .A0 (nx3028), .A1 (
          RST), .A2 (nx7862), .B0 (nx3004), .B1 (nx3024)) ;
    inv01 ix3027 (.Y (nx3028), .A (FilterDin_1__1__7)) ;
    nand02_2x L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix633 (.Y (nx3008), .A0 (
              nx7586), .A1 (nx7862)) ;
    nand02_2x L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix635 (.Y (nx3010), .A0 (
              nx7586), .A1 (nx7862)) ;
    oai32 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix393 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .A0 (nx8634), .A1 (
          RST), .A2 (nx7864), .B0 (nx2938), .B1 (nx3030)) ;
    oai32 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix403 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .A0 (nx8634), .A1 (
          RST), .A2 (nx7864), .B0 (nx2942), .B1 (nx3030)) ;
    oai32 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix413 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .A0 (nx8634), .A1 (
          RST), .A2 (nx7864), .B0 (nx2946), .B1 (nx3030)) ;
    oai32 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix423 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .A0 (nx8634), .A1 (
          RST), .A2 (nx7864), .B0 (nx2950), .B1 (nx3030)) ;
    oai32 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix433 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .A0 (nx8634), .A1 (
          RST), .A2 (nx7864), .B0 (nx2954), .B1 (nx3030)) ;
    oai32 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix443 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .A0 (nx8636), .A1 (
          RST), .A2 (nx7864), .B0 (nx2958), .B1 (nx3030)) ;
    oai32 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix453 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .A0 (nx8636), .A1 (
          RST), .A2 (nx7866), .B0 (nx2962), .B1 (nx3030)) ;
    oai32 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix463 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .A0 (nx8636), .A1 (
          RST), .A2 (nx7866), .B0 (nx2966), .B1 (nx3032)) ;
    oai32 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix473 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .A0 (nx8636), .A1 (
          RST), .A2 (nx7866), .B0 (nx2970), .B1 (nx3032)) ;
    oai32 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix483 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .A0 (nx3012), .A1 (
          RST), .A2 (nx7866), .B0 (nx2974), .B1 (nx3032)) ;
    oai32 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix493 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .A0 (nx3034), .A1 (
          RST), .A2 (nx7866), .B0 (nx2978), .B1 (nx3032)) ;
    inv01 ix3033 (.Y (nx3034), .A (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_10)) ;
    oai32 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix503 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .A0 (nx3036), .A1 (
          RST), .A2 (nx7866), .B0 (nx2982), .B1 (nx3032)) ;
    inv01 ix3035 (.Y (nx3036), .A (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_11)) ;
    oai32 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix513 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .A0 (nx3038), .A1 (
          RST), .A2 (nx7866), .B0 (nx2986), .B1 (nx3032)) ;
    inv01 ix3037 (.Y (nx3038), .A (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_12)) ;
    oai32 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix523 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .A0 (nx3040), .A1 (
          RST), .A2 (nx7868), .B0 (nx2990), .B1 (nx3032)) ;
    inv01 ix3039 (.Y (nx3040), .A (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_13)) ;
    oai32 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix533 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .A0 (nx3042), .A1 (
          RST), .A2 (nx7868), .B0 (nx2994), .B1 (nx3044)) ;
    inv01 ix3041 (.Y (nx3042), .A (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_14)) ;
    inv01 ix3043 (.Y (nx3044), .A (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566)) ;
    oai32 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix543 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .A0 (nx3046), .A1 (
          RST), .A2 (nx7868), .B0 (nx2998), .B1 (nx3044)) ;
    inv01 ix3045 (.Y (nx3046), .A (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_15)) ;
    oai32 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix553 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .A0 (nx3048), .A1 (
          RST), .A2 (nx7868), .B0 (nx3002), .B1 (nx3044)) ;
    inv01 ix3047 (.Y (nx3048), .A (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_16)) ;
    nand02_2x L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix633 (.Y (nx3030), .A0 (
              nx7586), .A1 (nx7868)) ;
    nand02_2x L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix635 (.Y (nx3032), .A0 (
              nx7586), .A1 (nx7868)) ;
    oai32 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix393 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .A0 (nx3050), .A1 (
          RST), .A2 (nx7870), .B0 (L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx384), .B1 (
          nx3052)) ;
    inv01 ix3049 (.Y (nx3050), .A (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_0)) ;
    oai32 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix403 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .A0 (nx3054), .A1 (
          RST), .A2 (nx7870), .B0 (nx2870), .B1 (nx3052)) ;
    inv01 ix3053 (.Y (nx3054), .A (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_1)) ;
    oai32 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix413 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .A0 (nx3056), .A1 (
          RST), .A2 (nx7870), .B0 (L1_1_L2_1_G1_MINI_ALU_nx387), .B1 (nx3052)) ;
    inv01 ix3055 (.Y (nx3056), .A (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_2)) ;
    oai32 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix423 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .A0 (nx3058), .A1 (
          RST), .A2 (nx7870), .B0 (L1_1_L2_1_G1_MINI_ALU_nx399), .B1 (nx3052)) ;
    inv01 ix3057 (.Y (nx3058), .A (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_3)) ;
    oai32 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix433 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .A0 (nx3060), .A1 (
          RST), .A2 (nx7870), .B0 (L1_1_L2_1_G1_MINI_ALU_nx409), .B1 (nx3052)) ;
    inv01 ix3059 (.Y (nx3060), .A (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_4)) ;
    oai32 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix443 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .A0 (nx3062), .A1 (
          RST), .A2 (nx7870), .B0 (L1_1_L2_1_G1_MINI_ALU_nx419), .B1 (nx3052)) ;
    inv01 ix3061 (.Y (nx3062), .A (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_5)) ;
    oai32 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix453 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .A0 (nx3064), .A1 (
          RST), .A2 (nx7870), .B0 (L1_1_L2_1_G1_MINI_ALU_nx429), .B1 (nx3052)) ;
    inv01 ix3063 (.Y (nx3064), .A (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_6)) ;
    oai32 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix463 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .A0 (nx3066), .A1 (
          RST), .A2 (nx7872), .B0 (L1_1_L2_1_G1_MINI_ALU_nx439), .B1 (nx3068)) ;
    inv01 ix3065 (.Y (nx3066), .A (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_7)) ;
    oai32 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix473 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .A0 (nx3070), .A1 (
          RST), .A2 (nx7872), .B0 (L1_1_L2_1_G1_MINI_ALU_nx449), .B1 (nx3068)) ;
    inv01 ix3069 (.Y (nx3070), .A (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_8)) ;
    oai32 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix483 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .A0 (nx3072), .A1 (
          RST), .A2 (nx7872), .B0 (L1_1_L2_1_G1_MINI_ALU_nx469), .B1 (nx3068)) ;
    inv01 ix3071 (.Y (nx3072), .A (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_9)) ;
    oai32 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix493 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .A0 (nx3074), .A1 (
          RST), .A2 (nx7872), .B0 (L1_1_L2_1_G1_MINI_ALU_nx477), .B1 (nx3068)) ;
    inv01 ix3073 (.Y (nx3074), .A (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_10)) ;
    oai32 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix503 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .A0 (nx3076), .A1 (
          RST), .A2 (nx7872), .B0 (L1_1_L2_1_G1_MINI_ALU_nx485), .B1 (nx3068)) ;
    inv01 ix3075 (.Y (nx3076), .A (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_11)) ;
    oai32 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix513 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .A0 (nx3078), .A1 (
          RST), .A2 (nx7872), .B0 (L1_1_L2_1_G1_MINI_ALU_nx493), .B1 (nx3068)) ;
    inv01 ix3077 (.Y (nx3078), .A (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_12)) ;
    oai32 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix523 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .A0 (nx3080), .A1 (
          RST), .A2 (nx7872), .B0 (L1_1_L2_1_G1_MINI_ALU_nx501), .B1 (nx3068)) ;
    inv01 ix3079 (.Y (nx3080), .A (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_13)) ;
    oai32 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix533 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .A0 (nx3082), .A1 (
          RST), .A2 (nx7874), .B0 (L1_1_L2_1_G1_MINI_ALU_nx509), .B1 (nx3084)) ;
    inv01 ix3081 (.Y (nx3082), .A (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_14)) ;
    inv01 ix3083 (.Y (nx3084), .A (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566)) ;
    oai32 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix543 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .A0 (nx3086), .A1 (
          RST), .A2 (nx7874), .B0 (L1_1_L2_1_G1_MINI_ALU_nx517), .B1 (nx3084)) ;
    inv01 ix3085 (.Y (nx3086), .A (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_15)) ;
    oai32 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix553 (.Y (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .A0 (nx3088), .A1 (
          RST), .A2 (nx7874), .B0 (nx2886), .B1 (nx3084)) ;
    inv01 ix3087 (.Y (nx3088), .A (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_16)) ;
    nand02_2x L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix633 (.Y (nx3052), .A0 (
              nx7586), .A1 (nx7874)) ;
    nand02_2x L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix635 (.Y (nx3068), .A0 (
              nx7586), .A1 (nx7874)) ;
    mux21 L1_1_L2_2_G1_MINI_ALU_ix404 (.Y (L1_1_L2_2_G1_MINI_ALU_nx403), .A0 (
          nx3090), .A1 (L1_1_L2_2_G1_MINI_ALU_BoothP_2), .S0 (
          L1_1_L2_2_G1_MINI_ALU_nx395)) ;
    inv01 ix3089 (.Y (nx3090), .A (L1_1_L2_2_G1_MINI_ALU_nx391)) ;
    mux21 L1_1_L2_2_G1_MINI_ALU_ix414 (.Y (L1_1_L2_2_G1_MINI_ALU_nx413), .A0 (
          nx3092), .A1 (L1_1_L2_2_G1_MINI_ALU_BoothP_3), .S0 (
          L1_1_L2_2_G1_MINI_ALU_nx405)) ;
    inv01 ix3091 (.Y (nx3092), .A (L1_1_L2_2_G1_MINI_ALU_nx403)) ;
    mux21 L1_1_L2_2_G1_MINI_ALU_ix424 (.Y (L1_1_L2_2_G1_MINI_ALU_nx423), .A0 (
          nx3094), .A1 (L1_1_L2_2_G1_MINI_ALU_BoothP_4), .S0 (
          L1_1_L2_2_G1_MINI_ALU_nx415)) ;
    inv01 ix3093 (.Y (nx3094), .A (L1_1_L2_2_G1_MINI_ALU_nx413)) ;
    mux21 L1_1_L2_2_G1_MINI_ALU_ix434 (.Y (L1_1_L2_2_G1_MINI_ALU_nx433), .A0 (
          nx3096), .A1 (L1_1_L2_2_G1_MINI_ALU_BoothP_5), .S0 (
          L1_1_L2_2_G1_MINI_ALU_nx425)) ;
    inv01 ix3095 (.Y (nx3096), .A (L1_1_L2_2_G1_MINI_ALU_nx423)) ;
    mux21 L1_1_L2_2_G1_MINI_ALU_ix444 (.Y (L1_1_L2_2_G1_MINI_ALU_nx443), .A0 (
          nx3098), .A1 (L1_1_L2_2_G1_MINI_ALU_BoothP_6), .S0 (
          L1_1_L2_2_G1_MINI_ALU_nx435)) ;
    inv01 ix3097 (.Y (nx3098), .A (L1_1_L2_2_G1_MINI_ALU_nx433)) ;
    mux21 L1_1_L2_2_G1_MINI_ALU_ix454 (.Y (L1_1_L2_2_G1_MINI_ALU_nx453), .A0 (
          nx3100), .A1 (L1_1_L2_2_G1_MINI_ALU_BoothP_7), .S0 (
          L1_1_L2_2_G1_MINI_ALU_nx445)) ;
    inv01 ix3099 (.Y (nx3100), .A (L1_1_L2_2_G1_MINI_ALU_nx443)) ;
    mux21 L1_1_L2_2_G1_MINI_ALU_ix462 (.Y (L1_1_L2_2_G1_MINI_ALU_nx461), .A0 (
          nx3102), .A1 (L1_1_L2_2_G1_MINI_ALU_BoothP_8), .S0 (
          L1_1_L2_2_G1_MINI_ALU_nx455)) ;
    inv01 ix3101 (.Y (nx3102), .A (L1_1_L2_2_G1_MINI_ALU_nx453)) ;
    mux21 L1_1_L2_2_G1_MINI_ALU_ix468 (.Y (L1_1_L2_2_G1_MINI_ALU_nx467), .A0 (
          nx3104), .A1 (L1_1_L2_2_G1_MINI_ALU_BoothP_9), .S0 (
          L1_1_L2_2_G1_MINI_ALU_nx463)) ;
    inv01 ix3103 (.Y (nx3104), .A (L1_1_L2_2_G1_MINI_ALU_nx461)) ;
    mux21 L1_1_L2_2_G1_MINI_ALU_ix476 (.Y (L1_1_L2_2_G1_MINI_ALU_nx475), .A0 (
          nx3106), .A1 (L1_1_L2_2_G1_MINI_ALU_BoothP_10), .S0 (
          L1_1_L2_2_G1_MINI_ALU_nx471)) ;
    inv01 ix3105 (.Y (nx3106), .A (L1_1_L2_2_G1_MINI_ALU_nx467)) ;
    mux21 L1_1_L2_2_G1_MINI_ALU_ix484 (.Y (L1_1_L2_2_G1_MINI_ALU_nx483), .A0 (
          nx3108), .A1 (L1_1_L2_2_G1_MINI_ALU_BoothP_11), .S0 (
          L1_1_L2_2_G1_MINI_ALU_nx479)) ;
    inv01 ix3107 (.Y (nx3108), .A (L1_1_L2_2_G1_MINI_ALU_nx475)) ;
    mux21 L1_1_L2_2_G1_MINI_ALU_ix492 (.Y (L1_1_L2_2_G1_MINI_ALU_nx491), .A0 (
          nx3110), .A1 (L1_1_L2_2_G1_MINI_ALU_BoothP_12), .S0 (
          L1_1_L2_2_G1_MINI_ALU_nx487)) ;
    inv01 ix3109 (.Y (nx3110), .A (L1_1_L2_2_G1_MINI_ALU_nx483)) ;
    mux21 L1_1_L2_2_G1_MINI_ALU_ix500 (.Y (L1_1_L2_2_G1_MINI_ALU_nx499), .A0 (
          nx3112), .A1 (L1_1_L2_2_G1_MINI_ALU_BoothP_13), .S0 (
          L1_1_L2_2_G1_MINI_ALU_nx495)) ;
    inv01 ix3111 (.Y (nx3112), .A (L1_1_L2_2_G1_MINI_ALU_nx491)) ;
    mux21 L1_1_L2_2_G1_MINI_ALU_ix508 (.Y (L1_1_L2_2_G1_MINI_ALU_nx507), .A0 (
          nx3114), .A1 (L1_1_L2_2_G1_MINI_ALU_BoothP_14), .S0 (
          L1_1_L2_2_G1_MINI_ALU_nx503)) ;
    inv01 ix3113 (.Y (nx3114), .A (L1_1_L2_2_G1_MINI_ALU_nx499)) ;
    mux21 L1_1_L2_2_G1_MINI_ALU_ix516 (.Y (L1_1_L2_2_G1_MINI_ALU_nx515), .A0 (
          nx3116), .A1 (L1_1_L2_2_G1_MINI_ALU_BoothP_15), .S0 (
          L1_1_L2_2_G1_MINI_ALU_nx511)) ;
    inv01 ix3115 (.Y (nx3116), .A (L1_1_L2_2_G1_MINI_ALU_nx507)) ;
    mux21 L1_1_L2_2_G1_MINI_ALU_ix161 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_1), .A0 (nx3118), .A1 (
          L1_1_L2_2_G1_MINI_ALU_nx379), .S0 (nx7878)) ;
    inv01 ix3117 (.Y (nx3118), .A (L1_1_L2_2_G1_MINI_ALU_BoothP_1)) ;
    mux21 L1_1_L2_2_G1_MINI_ALU_ix181 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_2), .A0 (
          L1_1_L2_2_G1_MINI_ALU_nx387), .A1 (L1_1_L2_2_G1_MINI_ALU_nx389), .S0 (
          nx7878)) ;
    mux21 L1_1_L2_2_G1_MINI_ALU_ix201 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_3), .A0 (
          L1_1_L2_2_G1_MINI_ALU_nx399), .A1 (L1_1_L2_2_G1_MINI_ALU_nx401), .S0 (
          nx7878)) ;
    mux21 L1_1_L2_2_G1_MINI_ALU_ix221 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_4), .A0 (
          L1_1_L2_2_G1_MINI_ALU_nx409), .A1 (L1_1_L2_2_G1_MINI_ALU_nx411), .S0 (
          nx7878)) ;
    mux21 L1_1_L2_2_G1_MINI_ALU_ix241 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_5), .A0 (
          L1_1_L2_2_G1_MINI_ALU_nx419), .A1 (L1_1_L2_2_G1_MINI_ALU_nx421), .S0 (
          nx7878)) ;
    mux21 L1_1_L2_2_G1_MINI_ALU_ix261 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_6), .A0 (
          L1_1_L2_2_G1_MINI_ALU_nx429), .A1 (L1_1_L2_2_G1_MINI_ALU_nx431), .S0 (
          nx7878)) ;
    mux21 L1_1_L2_2_G1_MINI_ALU_ix281 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_7), .A0 (
          L1_1_L2_2_G1_MINI_ALU_nx439), .A1 (L1_1_L2_2_G1_MINI_ALU_nx441), .S0 (
          nx7878)) ;
    mux21 L1_1_L2_2_G1_MINI_ALU_ix301 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_8), .A0 (
          L1_1_L2_2_G1_MINI_ALU_nx449), .A1 (L1_1_L2_2_G1_MINI_ALU_nx451), .S0 (
          nx7880)) ;
    mux21 L1_1_L2_2_G1_MINI_ALU_ix321 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_9), .A0 (
          L1_1_L2_2_G1_MINI_ALU_nx469), .A1 (nx3120), .S0 (nx7880)) ;
    inv01 ix3119 (.Y (nx3120), .A (L1_1_L2_2_G1_MINI_ALU_nx316)) ;
    mux21 L1_1_L2_2_G1_MINI_ALU_ix341 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_10), .A0 (
          L1_1_L2_2_G1_MINI_ALU_nx477), .A1 (nx3122), .S0 (nx7880)) ;
    inv01 ix3121 (.Y (nx3122), .A (L1_1_L2_2_G1_MINI_ALU_nx336)) ;
    mux21 L1_1_L2_2_G1_MINI_ALU_ix361 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_11), .A0 (
          L1_1_L2_2_G1_MINI_ALU_nx485), .A1 (nx3124), .S0 (nx7880)) ;
    inv01 ix3123 (.Y (nx3124), .A (L1_1_L2_2_G1_MINI_ALU_nx356)) ;
    mux21 L1_1_L2_2_G1_MINI_ALU_ix381 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_12), .A0 (
          L1_1_L2_2_G1_MINI_ALU_nx493), .A1 (nx3126), .S0 (nx7880)) ;
    inv01 ix3125 (.Y (nx3126), .A (L1_1_L2_2_G1_MINI_ALU_nx376)) ;
    mux21 L1_1_L2_2_G1_MINI_ALU_ix401 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_13), .A0 (
          L1_1_L2_2_G1_MINI_ALU_nx501), .A1 (nx3128), .S0 (nx7880)) ;
    inv01 ix3127 (.Y (nx3128), .A (L1_1_L2_2_G1_MINI_ALU_nx396)) ;
    mux21 L1_1_L2_2_G1_MINI_ALU_ix421 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_14), .A0 (
          L1_1_L2_2_G1_MINI_ALU_nx509), .A1 (nx3130), .S0 (nx7880)) ;
    inv01 ix3129 (.Y (nx3130), .A (L1_1_L2_2_G1_MINI_ALU_nx416)) ;
    mux21 L1_1_L2_2_G1_MINI_ALU_ix441 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_15), .A0 (
          L1_1_L2_2_G1_MINI_ALU_nx517), .A1 (nx3132), .S0 (nx7882)) ;
    inv01 ix3131 (.Y (nx3132), .A (L1_1_L2_2_G1_MINI_ALU_nx436)) ;
    mux21 L1_1_L2_2_G1_MINI_ALU_ix461 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_16), .A0 (nx3134), .A1 (nx3136
          ), .S0 (nx7882)) ;
    inv01 ix3133 (.Y (nx3134), .A (L1_1_L2_2_G1_MINI_ALU_BoothP_16)) ;
    inv01 ix3135 (.Y (nx3136), .A (L1_1_L2_2_G1_MINI_ALU_nx456)) ;
    nor02_2x L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix319 (.Y (
             L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642), .A0 (Start), .A1 (
             CalculatingBooth_dup_1119)) ;
    nor02_2x L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix85 (.Y (
             L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_0), .A0 (nx7892), .A1 (
             nx3138)) ;
    inv01 ix3137 (.Y (nx3138), .A (L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_1)) ;
    mux21 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix125 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_1), .A0 (nx3140), .A1 (
          nx3142), .S0 (nx7892)) ;
    inv01 ix3139 (.Y (nx3140), .A (L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_2)) ;
    inv01 ix3141 (.Y (nx3142), .A (WindowDin_1__2__0)) ;
    mux21 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix133 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_2), .A0 (nx3144), .A1 (
          nx3146), .S0 (nx7892)) ;
    inv01 ix3143 (.Y (nx3144), .A (L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_3)) ;
    inv01 ix3145 (.Y (nx3146), .A (WindowDin_1__2__1)) ;
    mux21 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix141 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_3), .A0 (nx3148), .A1 (
          nx3150), .S0 (nx7892)) ;
    inv01 ix3147 (.Y (nx3148), .A (L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_4)) ;
    inv01 ix3149 (.Y (nx3150), .A (WindowDin_1__2__2)) ;
    mux21 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix149 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_4), .A0 (nx3152), .A1 (
          nx3154), .S0 (nx7892)) ;
    inv01 ix3151 (.Y (nx3152), .A (L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_5)) ;
    inv01 ix3153 (.Y (nx3154), .A (WindowDin_1__2__3)) ;
    mux21 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix157 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_5), .A0 (nx3156), .A1 (
          nx3158), .S0 (nx7892)) ;
    inv01 ix3155 (.Y (nx3156), .A (L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_6)) ;
    inv01 ix3157 (.Y (nx3158), .A (WindowDin_1__2__4)) ;
    mux21 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix165 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_6), .A0 (nx3160), .A1 (
          nx3162), .S0 (nx7892)) ;
    inv01 ix3159 (.Y (nx3160), .A (L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_7)) ;
    inv01 ix3161 (.Y (nx3162), .A (WindowDin_1__2__5)) ;
    mux21 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix173 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_7), .A0 (nx3164), .A1 (
          nx3166), .S0 (nx7894)) ;
    inv01 ix3163 (.Y (nx3164), .A (L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_8)) ;
    inv01 ix3165 (.Y (nx3166), .A (WindowDin_1__2__6)) ;
    mux21 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix181 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_8), .A0 (nx3168), .A1 (
          nx3170), .S0 (nx7894)) ;
    inv01 ix3167 (.Y (nx3168), .A (L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_9)) ;
    inv01 ix3169 (.Y (nx3170), .A (WindowDin_1__2__7)) ;
    nor02_2x L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix89 (.Y (
             L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_9), .A0 (nx7894), .A1 (
             nx3172)) ;
    inv01 ix3171 (.Y (nx3172), .A (L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_10)
          ) ;
    nor02_2x L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix93 (.Y (
             L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_10), .A0 (nx7894), .A1 (
             nx3174)) ;
    inv01 ix3173 (.Y (nx3174), .A (L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_11)
          ) ;
    nor02_2x L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix97 (.Y (
             L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_11), .A0 (nx7894), .A1 (
             nx3176)) ;
    inv01 ix3175 (.Y (nx3176), .A (L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_12)
          ) ;
    nor02_2x L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix101 (.Y (
             L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_12), .A0 (nx7894), .A1 (
             nx3178)) ;
    inv01 ix3177 (.Y (nx3178), .A (L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_13)
          ) ;
    nor02_2x L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix105 (.Y (
             L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_13), .A0 (nx7894), .A1 (
             nx3180)) ;
    inv01 ix3179 (.Y (nx3180), .A (L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_14)
          ) ;
    nor02_2x L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix109 (.Y (
             L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_14), .A0 (nx7896), .A1 (
             nx3182)) ;
    inv01 ix3181 (.Y (nx3182), .A (L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_15)
          ) ;
    nor02_2x L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix113 (.Y (
             L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_15), .A0 (nx7896), .A1 (
             nx3184)) ;
    inv01 ix3183 (.Y (nx3184), .A (L1_1_L2_2_G1_MINI_ALU_BoothPBeforeShift_16)
          ) ;
    nor02_2x L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix117 (.Y (
             L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_16), .A0 (nx7896), .A1 (
             nx3184)) ;
    mux21 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix189 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BoothOperand_0), .A0 (nx3186), .A1 (nx3188), .S0 (
          nx7884)) ;
    inv01 ix3185 (.Y (nx3186), .A (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_0)) ;
    inv01 ix3187 (.Y (nx3188), .A (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_0)) ;
    mux21 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix197 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BoothOperand_1), .A0 (nx3190), .A1 (nx3192), .S0 (
          nx7884)) ;
    inv01 ix3189 (.Y (nx3190), .A (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_1)) ;
    inv01 ix3191 (.Y (nx3192), .A (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_1)) ;
    mux21 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix205 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BoothOperand_2), .A0 (nx3194), .A1 (nx3196), .S0 (
          nx7884)) ;
    inv01 ix3193 (.Y (nx3194), .A (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_2)) ;
    inv01 ix3195 (.Y (nx3196), .A (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_2)) ;
    mux21 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix213 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BoothOperand_3), .A0 (nx3198), .A1 (nx3200), .S0 (
          nx7884)) ;
    inv01 ix3197 (.Y (nx3198), .A (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_3)) ;
    inv01 ix3199 (.Y (nx3200), .A (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_3)) ;
    mux21 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix221 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BoothOperand_4), .A0 (nx3202), .A1 (nx3204), .S0 (
          nx7884)) ;
    inv01 ix3201 (.Y (nx3202), .A (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_4)) ;
    inv01 ix3203 (.Y (nx3204), .A (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_4)) ;
    mux21 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix229 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BoothOperand_5), .A0 (nx3206), .A1 (nx3208), .S0 (
          nx7886)) ;
    inv01 ix3205 (.Y (nx3206), .A (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_5)) ;
    inv01 ix3207 (.Y (nx3208), .A (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_5)) ;
    mux21 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix237 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BoothOperand_6), .A0 (nx3210), .A1 (nx3212), .S0 (
          nx7886)) ;
    inv01 ix3209 (.Y (nx3210), .A (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_6)) ;
    inv01 ix3211 (.Y (nx3212), .A (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_6)) ;
    mux21 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix245 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BoothOperand_7), .A0 (nx3214), .A1 (nx3216), .S0 (
          nx7886)) ;
    inv01 ix3213 (.Y (nx3214), .A (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_7)) ;
    inv01 ix3215 (.Y (nx3216), .A (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_7)) ;
    mux21 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix253 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BoothOperand_8), .A0 (nx3218), .A1 (nx3220), .S0 (
          nx7886)) ;
    inv01 ix3217 (.Y (nx3218), .A (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_8)) ;
    inv01 ix3219 (.Y (nx3220), .A (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_8)) ;
    mux21 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix261 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BoothOperand_9), .A0 (nx3222), .A1 (nx3224), .S0 (
          nx7886)) ;
    inv01 ix3221 (.Y (nx3222), .A (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_9)) ;
    inv01 ix3223 (.Y (nx3224), .A (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_9)) ;
    mux21 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix269 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BoothOperand_10), .A0 (nx3226), .A1 (nx3228), .S0 (
          nx7886)) ;
    inv01 ix3225 (.Y (nx3226), .A (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_10)) ;
    inv01 ix3227 (.Y (nx3228), .A (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_10)) ;
    mux21 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix277 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BoothOperand_11), .A0 (nx3230), .A1 (nx3232), .S0 (
          nx7886)) ;
    inv01 ix3229 (.Y (nx3230), .A (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_11)) ;
    inv01 ix3231 (.Y (nx3232), .A (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_11)) ;
    mux21 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix285 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BoothOperand_12), .A0 (nx3234), .A1 (nx3236), .S0 (
          nx7888)) ;
    inv01 ix3233 (.Y (nx3234), .A (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_12)) ;
    inv01 ix3235 (.Y (nx3236), .A (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_12)) ;
    mux21 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix293 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BoothOperand_13), .A0 (nx3238), .A1 (nx3240), .S0 (
          nx7888)) ;
    inv01 ix3237 (.Y (nx3238), .A (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_13)) ;
    inv01 ix3239 (.Y (nx3240), .A (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_13)) ;
    mux21 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix301 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BoothOperand_14), .A0 (nx3242), .A1 (nx3244), .S0 (
          nx7888)) ;
    inv01 ix3241 (.Y (nx3242), .A (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_14)) ;
    inv01 ix3243 (.Y (nx3244), .A (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_14)) ;
    mux21 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix309 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BoothOperand_15), .A0 (nx3246), .A1 (nx3248), .S0 (
          nx7888)) ;
    inv01 ix3245 (.Y (nx3246), .A (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_15)) ;
    inv01 ix3247 (.Y (nx3248), .A (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_15)) ;
    mux21 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix317 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BoothOperand_16), .A0 (nx3250), .A1 (nx3252), .S0 (
          nx7888)) ;
    inv01 ix3249 (.Y (nx3250), .A (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_16)) ;
    inv01 ix3251 (.Y (nx3252), .A (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_16)) ;
    xnor2 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix321 (.Y (
          L1_1_L2_2_G1_MINI_ALU_AddPToBoothOperand), .A0 (nx7888), .A1 (nx3118)
          ) ;
    oai32 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix393 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .A0 (nx8638), .A1 (
          RST), .A2 (nx7898), .B0 (nx3188), .B1 (nx3256)) ;
    oai32 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix403 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .A0 (nx8638), .A1 (
          RST), .A2 (nx7898), .B0 (nx3192), .B1 (nx3256)) ;
    oai32 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix413 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .A0 (nx8638), .A1 (
          RST), .A2 (nx7898), .B0 (nx3196), .B1 (nx3256)) ;
    oai32 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix423 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .A0 (nx8638), .A1 (
          RST), .A2 (nx7898), .B0 (nx3200), .B1 (nx3256)) ;
    oai32 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix433 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .A0 (nx8638), .A1 (
          RST), .A2 (nx7898), .B0 (nx3204), .B1 (nx3256)) ;
    oai32 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix443 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .A0 (nx8638), .A1 (
          RST), .A2 (nx7898), .B0 (nx3208), .B1 (nx3256)) ;
    oai32 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix453 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .A0 (nx8638), .A1 (
          RST), .A2 (nx7900), .B0 (nx3212), .B1 (nx3256)) ;
    oai32 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix463 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .A0 (nx8640), .A1 (
          RST), .A2 (nx7900), .B0 (nx3216), .B1 (nx3258)) ;
    oai32 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix473 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .A0 (nx8640), .A1 (
          RST), .A2 (nx7900), .B0 (nx3220), .B1 (nx3258)) ;
    oai32 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix483 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .A0 (nx3260), .A1 (
          RST), .A2 (nx7900), .B0 (nx3224), .B1 (nx3258)) ;
    inv01 ix3259 (.Y (nx3260), .A (FilterDin_1__2__0)) ;
    oai32 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix493 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .A0 (nx3262), .A1 (
          RST), .A2 (nx7900), .B0 (nx3228), .B1 (nx3258)) ;
    inv01 ix3261 (.Y (nx3262), .A (FilterDin_1__2__1)) ;
    oai32 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix503 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .A0 (nx3264), .A1 (
          RST), .A2 (nx7900), .B0 (nx3232), .B1 (nx3258)) ;
    inv01 ix3263 (.Y (nx3264), .A (FilterDin_1__2__2)) ;
    oai32 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix513 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .A0 (nx3266), .A1 (
          RST), .A2 (nx7900), .B0 (nx3236), .B1 (nx3258)) ;
    inv01 ix3265 (.Y (nx3266), .A (FilterDin_1__2__3)) ;
    oai32 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix523 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .A0 (nx3268), .A1 (
          RST), .A2 (nx7902), .B0 (nx3240), .B1 (nx3258)) ;
    inv01 ix3267 (.Y (nx3268), .A (FilterDin_1__2__4)) ;
    oai32 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix533 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .A0 (nx3270), .A1 (
          RST), .A2 (nx7902), .B0 (nx3244), .B1 (nx3272)) ;
    inv01 ix3269 (.Y (nx3270), .A (FilterDin_1__2__5)) ;
    inv01 ix3271 (.Y (nx3272), .A (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566)) ;
    oai32 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix543 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .A0 (nx3274), .A1 (
          RST), .A2 (nx7902), .B0 (nx3248), .B1 (nx3272)) ;
    inv01 ix3273 (.Y (nx3274), .A (FilterDin_1__2__6)) ;
    oai32 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix553 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .A0 (nx3276), .A1 (
          RST), .A2 (nx7902), .B0 (nx3252), .B1 (nx3272)) ;
    inv01 ix3275 (.Y (nx3276), .A (FilterDin_1__2__7)) ;
    nand02_2x L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix633 (.Y (nx3256), .A0 (
              nx7588), .A1 (nx7902)) ;
    nand02_2x L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix635 (.Y (nx3258), .A0 (
              nx7588), .A1 (nx7902)) ;
    oai32 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix393 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .A0 (nx8640), .A1 (
          RST), .A2 (nx7904), .B0 (nx3186), .B1 (nx3278)) ;
    oai32 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix403 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .A0 (nx8640), .A1 (
          RST), .A2 (nx7904), .B0 (nx3190), .B1 (nx3278)) ;
    oai32 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix413 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .A0 (nx8640), .A1 (
          RST), .A2 (nx7904), .B0 (nx3194), .B1 (nx3278)) ;
    oai32 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix423 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .A0 (nx8640), .A1 (
          RST), .A2 (nx7904), .B0 (nx3198), .B1 (nx3278)) ;
    oai32 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix433 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .A0 (nx8640), .A1 (
          RST), .A2 (nx7904), .B0 (nx3202), .B1 (nx3278)) ;
    oai32 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix443 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .A0 (nx8642), .A1 (
          RST), .A2 (nx7904), .B0 (nx3206), .B1 (nx3278)) ;
    oai32 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix453 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .A0 (nx8642), .A1 (
          RST), .A2 (nx7906), .B0 (nx3210), .B1 (nx3278)) ;
    oai32 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix463 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .A0 (nx8642), .A1 (
          RST), .A2 (nx7906), .B0 (nx3214), .B1 (nx3280)) ;
    oai32 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix473 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .A0 (nx8642), .A1 (
          RST), .A2 (nx7906), .B0 (nx3218), .B1 (nx3280)) ;
    oai32 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix483 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .A0 (nx3260), .A1 (
          RST), .A2 (nx7906), .B0 (nx3222), .B1 (nx3280)) ;
    oai32 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix493 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .A0 (nx3282), .A1 (
          RST), .A2 (nx7906), .B0 (nx3226), .B1 (nx3280)) ;
    inv01 ix3281 (.Y (nx3282), .A (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_10)) ;
    oai32 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix503 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .A0 (nx3284), .A1 (
          RST), .A2 (nx7906), .B0 (nx3230), .B1 (nx3280)) ;
    inv01 ix3283 (.Y (nx3284), .A (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_11)) ;
    oai32 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix513 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .A0 (nx3286), .A1 (
          RST), .A2 (nx7906), .B0 (nx3234), .B1 (nx3280)) ;
    inv01 ix3285 (.Y (nx3286), .A (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_12)) ;
    oai32 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix523 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .A0 (nx3288), .A1 (
          RST), .A2 (nx7908), .B0 (nx3238), .B1 (nx3280)) ;
    inv01 ix3287 (.Y (nx3288), .A (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_13)) ;
    oai32 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix533 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .A0 (nx3290), .A1 (
          RST), .A2 (nx7908), .B0 (nx3242), .B1 (nx3292)) ;
    inv01 ix3289 (.Y (nx3290), .A (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_14)) ;
    inv01 ix3291 (.Y (nx3292), .A (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566)) ;
    oai32 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix543 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .A0 (nx3294), .A1 (
          RST), .A2 (nx7908), .B0 (nx3246), .B1 (nx3292)) ;
    inv01 ix3293 (.Y (nx3294), .A (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_15)) ;
    oai32 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix553 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .A0 (nx3296), .A1 (
          RST), .A2 (nx7908), .B0 (nx3250), .B1 (nx3292)) ;
    inv01 ix3295 (.Y (nx3296), .A (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_16)) ;
    nand02_2x L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix633 (.Y (nx3278), .A0 (
              nx7588), .A1 (nx7908)) ;
    nand02_2x L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix635 (.Y (nx3280), .A0 (
              nx7588), .A1 (nx7908)) ;
    oai32 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix393 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .A0 (nx3298), .A1 (
          RST), .A2 (nx7910), .B0 (L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx384), .B1 (
          nx3300)) ;
    inv01 ix3297 (.Y (nx3298), .A (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_0)) ;
    oai32 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix403 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .A0 (nx3302), .A1 (
          RST), .A2 (nx7910), .B0 (nx3118), .B1 (nx3300)) ;
    inv01 ix3301 (.Y (nx3302), .A (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_1)) ;
    oai32 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix413 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .A0 (nx3304), .A1 (
          RST), .A2 (nx7910), .B0 (L1_1_L2_2_G1_MINI_ALU_nx387), .B1 (nx3300)) ;
    inv01 ix3303 (.Y (nx3304), .A (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_2)) ;
    oai32 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix423 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .A0 (nx3306), .A1 (
          RST), .A2 (nx7910), .B0 (L1_1_L2_2_G1_MINI_ALU_nx399), .B1 (nx3300)) ;
    inv01 ix3305 (.Y (nx3306), .A (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_3)) ;
    oai32 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix433 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .A0 (nx3308), .A1 (
          RST), .A2 (nx7910), .B0 (L1_1_L2_2_G1_MINI_ALU_nx409), .B1 (nx3300)) ;
    inv01 ix3307 (.Y (nx3308), .A (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_4)) ;
    oai32 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix443 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .A0 (nx3310), .A1 (
          RST), .A2 (nx7910), .B0 (L1_1_L2_2_G1_MINI_ALU_nx419), .B1 (nx3300)) ;
    inv01 ix3309 (.Y (nx3310), .A (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_5)) ;
    oai32 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix453 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .A0 (nx3312), .A1 (
          RST), .A2 (nx7910), .B0 (L1_1_L2_2_G1_MINI_ALU_nx429), .B1 (nx3300)) ;
    inv01 ix3311 (.Y (nx3312), .A (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_6)) ;
    oai32 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix463 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .A0 (nx3314), .A1 (
          RST), .A2 (nx7912), .B0 (L1_1_L2_2_G1_MINI_ALU_nx439), .B1 (nx3316)) ;
    inv01 ix3313 (.Y (nx3314), .A (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_7)) ;
    oai32 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix473 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .A0 (nx3318), .A1 (
          RST), .A2 (nx7912), .B0 (L1_1_L2_2_G1_MINI_ALU_nx449), .B1 (nx3316)) ;
    inv01 ix3317 (.Y (nx3318), .A (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_8)) ;
    oai32 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix483 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .A0 (nx3320), .A1 (
          RST), .A2 (nx7912), .B0 (L1_1_L2_2_G1_MINI_ALU_nx469), .B1 (nx3316)) ;
    inv01 ix3319 (.Y (nx3320), .A (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_9)) ;
    oai32 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix493 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .A0 (nx3322), .A1 (
          RST), .A2 (nx7912), .B0 (L1_1_L2_2_G1_MINI_ALU_nx477), .B1 (nx3316)) ;
    inv01 ix3321 (.Y (nx3322), .A (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_10)) ;
    oai32 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix503 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .A0 (nx3324), .A1 (
          RST), .A2 (nx7912), .B0 (L1_1_L2_2_G1_MINI_ALU_nx485), .B1 (nx3316)) ;
    inv01 ix3323 (.Y (nx3324), .A (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_11)) ;
    oai32 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix513 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .A0 (nx3326), .A1 (
          RST), .A2 (nx7912), .B0 (L1_1_L2_2_G1_MINI_ALU_nx493), .B1 (nx3316)) ;
    inv01 ix3325 (.Y (nx3326), .A (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_12)) ;
    oai32 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix523 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .A0 (nx3328), .A1 (
          RST), .A2 (nx7912), .B0 (L1_1_L2_2_G1_MINI_ALU_nx501), .B1 (nx3316)) ;
    inv01 ix3327 (.Y (nx3328), .A (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_13)) ;
    oai32 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix533 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .A0 (nx3330), .A1 (
          RST), .A2 (nx7914), .B0 (L1_1_L2_2_G1_MINI_ALU_nx509), .B1 (nx3332)) ;
    inv01 ix3329 (.Y (nx3330), .A (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_14)) ;
    inv01 ix3331 (.Y (nx3332), .A (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566)) ;
    oai32 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix543 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .A0 (nx3334), .A1 (
          RST), .A2 (nx7914), .B0 (L1_1_L2_2_G1_MINI_ALU_nx517), .B1 (nx3332)) ;
    inv01 ix3333 (.Y (nx3334), .A (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_15)) ;
    oai32 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix553 (.Y (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .A0 (nx3336), .A1 (
          RST), .A2 (nx7914), .B0 (nx3134), .B1 (nx3332)) ;
    inv01 ix3335 (.Y (nx3336), .A (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_16)) ;
    nand02_2x L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix633 (.Y (nx3300), .A0 (
              nx7588), .A1 (nx7914)) ;
    nand02_2x L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix635 (.Y (nx3316), .A0 (
              nx7588), .A1 (nx7914)) ;
    mux21 L1_1_L2_3_G1_MINI_ALU_ix404 (.Y (L1_1_L2_3_G1_MINI_ALU_nx403), .A0 (
          nx3338), .A1 (L1_1_L2_3_G1_MINI_ALU_BoothP_2), .S0 (
          L1_1_L2_3_G1_MINI_ALU_nx395)) ;
    inv01 ix3337 (.Y (nx3338), .A (L1_1_L2_3_G1_MINI_ALU_nx391)) ;
    mux21 L1_1_L2_3_G1_MINI_ALU_ix414 (.Y (L1_1_L2_3_G1_MINI_ALU_nx413), .A0 (
          nx3340), .A1 (L1_1_L2_3_G1_MINI_ALU_BoothP_3), .S0 (
          L1_1_L2_3_G1_MINI_ALU_nx405)) ;
    inv01 ix3339 (.Y (nx3340), .A (L1_1_L2_3_G1_MINI_ALU_nx403)) ;
    mux21 L1_1_L2_3_G1_MINI_ALU_ix424 (.Y (L1_1_L2_3_G1_MINI_ALU_nx423), .A0 (
          nx3342), .A1 (L1_1_L2_3_G1_MINI_ALU_BoothP_4), .S0 (
          L1_1_L2_3_G1_MINI_ALU_nx415)) ;
    inv01 ix3341 (.Y (nx3342), .A (L1_1_L2_3_G1_MINI_ALU_nx413)) ;
    mux21 L1_1_L2_3_G1_MINI_ALU_ix434 (.Y (L1_1_L2_3_G1_MINI_ALU_nx433), .A0 (
          nx3344), .A1 (L1_1_L2_3_G1_MINI_ALU_BoothP_5), .S0 (
          L1_1_L2_3_G1_MINI_ALU_nx425)) ;
    inv01 ix3343 (.Y (nx3344), .A (L1_1_L2_3_G1_MINI_ALU_nx423)) ;
    mux21 L1_1_L2_3_G1_MINI_ALU_ix444 (.Y (L1_1_L2_3_G1_MINI_ALU_nx443), .A0 (
          nx3346), .A1 (L1_1_L2_3_G1_MINI_ALU_BoothP_6), .S0 (
          L1_1_L2_3_G1_MINI_ALU_nx435)) ;
    inv01 ix3345 (.Y (nx3346), .A (L1_1_L2_3_G1_MINI_ALU_nx433)) ;
    mux21 L1_1_L2_3_G1_MINI_ALU_ix454 (.Y (L1_1_L2_3_G1_MINI_ALU_nx453), .A0 (
          nx3348), .A1 (L1_1_L2_3_G1_MINI_ALU_BoothP_7), .S0 (
          L1_1_L2_3_G1_MINI_ALU_nx445)) ;
    inv01 ix3347 (.Y (nx3348), .A (L1_1_L2_3_G1_MINI_ALU_nx443)) ;
    mux21 L1_1_L2_3_G1_MINI_ALU_ix462 (.Y (L1_1_L2_3_G1_MINI_ALU_nx461), .A0 (
          nx3350), .A1 (L1_1_L2_3_G1_MINI_ALU_BoothP_8), .S0 (
          L1_1_L2_3_G1_MINI_ALU_nx455)) ;
    inv01 ix3349 (.Y (nx3350), .A (L1_1_L2_3_G1_MINI_ALU_nx453)) ;
    mux21 L1_1_L2_3_G1_MINI_ALU_ix468 (.Y (L1_1_L2_3_G1_MINI_ALU_nx467), .A0 (
          nx3352), .A1 (L1_1_L2_3_G1_MINI_ALU_BoothP_9), .S0 (
          L1_1_L2_3_G1_MINI_ALU_nx463)) ;
    inv01 ix3351 (.Y (nx3352), .A (L1_1_L2_3_G1_MINI_ALU_nx461)) ;
    mux21 L1_1_L2_3_G1_MINI_ALU_ix476 (.Y (L1_1_L2_3_G1_MINI_ALU_nx475), .A0 (
          nx3354), .A1 (L1_1_L2_3_G1_MINI_ALU_BoothP_10), .S0 (
          L1_1_L2_3_G1_MINI_ALU_nx471)) ;
    inv01 ix3353 (.Y (nx3354), .A (L1_1_L2_3_G1_MINI_ALU_nx467)) ;
    mux21 L1_1_L2_3_G1_MINI_ALU_ix484 (.Y (L1_1_L2_3_G1_MINI_ALU_nx483), .A0 (
          nx3356), .A1 (L1_1_L2_3_G1_MINI_ALU_BoothP_11), .S0 (
          L1_1_L2_3_G1_MINI_ALU_nx479)) ;
    inv01 ix3355 (.Y (nx3356), .A (L1_1_L2_3_G1_MINI_ALU_nx475)) ;
    mux21 L1_1_L2_3_G1_MINI_ALU_ix492 (.Y (L1_1_L2_3_G1_MINI_ALU_nx491), .A0 (
          nx3358), .A1 (L1_1_L2_3_G1_MINI_ALU_BoothP_12), .S0 (
          L1_1_L2_3_G1_MINI_ALU_nx487)) ;
    inv01 ix3357 (.Y (nx3358), .A (L1_1_L2_3_G1_MINI_ALU_nx483)) ;
    mux21 L1_1_L2_3_G1_MINI_ALU_ix500 (.Y (L1_1_L2_3_G1_MINI_ALU_nx499), .A0 (
          nx3360), .A1 (L1_1_L2_3_G1_MINI_ALU_BoothP_13), .S0 (
          L1_1_L2_3_G1_MINI_ALU_nx495)) ;
    inv01 ix3359 (.Y (nx3360), .A (L1_1_L2_3_G1_MINI_ALU_nx491)) ;
    mux21 L1_1_L2_3_G1_MINI_ALU_ix508 (.Y (L1_1_L2_3_G1_MINI_ALU_nx507), .A0 (
          nx3362), .A1 (L1_1_L2_3_G1_MINI_ALU_BoothP_14), .S0 (
          L1_1_L2_3_G1_MINI_ALU_nx503)) ;
    inv01 ix3361 (.Y (nx3362), .A (L1_1_L2_3_G1_MINI_ALU_nx499)) ;
    mux21 L1_1_L2_3_G1_MINI_ALU_ix516 (.Y (L1_1_L2_3_G1_MINI_ALU_nx515), .A0 (
          nx3364), .A1 (L1_1_L2_3_G1_MINI_ALU_BoothP_15), .S0 (
          L1_1_L2_3_G1_MINI_ALU_nx511)) ;
    inv01 ix3363 (.Y (nx3364), .A (L1_1_L2_3_G1_MINI_ALU_nx507)) ;
    mux21 L1_1_L2_3_G1_MINI_ALU_ix161 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_1), .A0 (nx3366), .A1 (
          L1_1_L2_3_G1_MINI_ALU_nx379), .S0 (nx7918)) ;
    inv01 ix3365 (.Y (nx3366), .A (L1_1_L2_3_G1_MINI_ALU_BoothP_1)) ;
    mux21 L1_1_L2_3_G1_MINI_ALU_ix181 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_2), .A0 (
          L1_1_L2_3_G1_MINI_ALU_nx387), .A1 (L1_1_L2_3_G1_MINI_ALU_nx389), .S0 (
          nx7918)) ;
    mux21 L1_1_L2_3_G1_MINI_ALU_ix201 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_3), .A0 (
          L1_1_L2_3_G1_MINI_ALU_nx399), .A1 (L1_1_L2_3_G1_MINI_ALU_nx401), .S0 (
          nx7918)) ;
    mux21 L1_1_L2_3_G1_MINI_ALU_ix221 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_4), .A0 (
          L1_1_L2_3_G1_MINI_ALU_nx409), .A1 (L1_1_L2_3_G1_MINI_ALU_nx411), .S0 (
          nx7918)) ;
    mux21 L1_1_L2_3_G1_MINI_ALU_ix241 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_5), .A0 (
          L1_1_L2_3_G1_MINI_ALU_nx419), .A1 (L1_1_L2_3_G1_MINI_ALU_nx421), .S0 (
          nx7918)) ;
    mux21 L1_1_L2_3_G1_MINI_ALU_ix261 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_6), .A0 (
          L1_1_L2_3_G1_MINI_ALU_nx429), .A1 (L1_1_L2_3_G1_MINI_ALU_nx431), .S0 (
          nx7918)) ;
    mux21 L1_1_L2_3_G1_MINI_ALU_ix281 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_7), .A0 (
          L1_1_L2_3_G1_MINI_ALU_nx439), .A1 (L1_1_L2_3_G1_MINI_ALU_nx441), .S0 (
          nx7918)) ;
    mux21 L1_1_L2_3_G1_MINI_ALU_ix301 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_8), .A0 (
          L1_1_L2_3_G1_MINI_ALU_nx449), .A1 (L1_1_L2_3_G1_MINI_ALU_nx451), .S0 (
          nx7920)) ;
    mux21 L1_1_L2_3_G1_MINI_ALU_ix321 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_9), .A0 (
          L1_1_L2_3_G1_MINI_ALU_nx469), .A1 (nx3368), .S0 (nx7920)) ;
    inv01 ix3367 (.Y (nx3368), .A (L1_1_L2_3_G1_MINI_ALU_nx316)) ;
    mux21 L1_1_L2_3_G1_MINI_ALU_ix341 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_10), .A0 (
          L1_1_L2_3_G1_MINI_ALU_nx477), .A1 (nx3370), .S0 (nx7920)) ;
    inv01 ix3369 (.Y (nx3370), .A (L1_1_L2_3_G1_MINI_ALU_nx336)) ;
    mux21 L1_1_L2_3_G1_MINI_ALU_ix361 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_11), .A0 (
          L1_1_L2_3_G1_MINI_ALU_nx485), .A1 (nx3372), .S0 (nx7920)) ;
    inv01 ix3371 (.Y (nx3372), .A (L1_1_L2_3_G1_MINI_ALU_nx356)) ;
    mux21 L1_1_L2_3_G1_MINI_ALU_ix381 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_12), .A0 (
          L1_1_L2_3_G1_MINI_ALU_nx493), .A1 (nx3374), .S0 (nx7920)) ;
    inv01 ix3373 (.Y (nx3374), .A (L1_1_L2_3_G1_MINI_ALU_nx376)) ;
    mux21 L1_1_L2_3_G1_MINI_ALU_ix401 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_13), .A0 (
          L1_1_L2_3_G1_MINI_ALU_nx501), .A1 (nx3376), .S0 (nx7920)) ;
    inv01 ix3375 (.Y (nx3376), .A (L1_1_L2_3_G1_MINI_ALU_nx396)) ;
    mux21 L1_1_L2_3_G1_MINI_ALU_ix421 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_14), .A0 (
          L1_1_L2_3_G1_MINI_ALU_nx509), .A1 (nx3378), .S0 (nx7920)) ;
    inv01 ix3377 (.Y (nx3378), .A (L1_1_L2_3_G1_MINI_ALU_nx416)) ;
    mux21 L1_1_L2_3_G1_MINI_ALU_ix441 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_15), .A0 (
          L1_1_L2_3_G1_MINI_ALU_nx517), .A1 (nx3380), .S0 (nx7922)) ;
    inv01 ix3379 (.Y (nx3380), .A (L1_1_L2_3_G1_MINI_ALU_nx436)) ;
    mux21 L1_1_L2_3_G1_MINI_ALU_ix461 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_16), .A0 (nx3382), .A1 (nx3384
          ), .S0 (nx7922)) ;
    inv01 ix3381 (.Y (nx3382), .A (L1_1_L2_3_G1_MINI_ALU_BoothP_16)) ;
    inv01 ix3383 (.Y (nx3384), .A (L1_1_L2_3_G1_MINI_ALU_nx456)) ;
    nor02_2x L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix319 (.Y (
             L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642), .A0 (Start), .A1 (
             CalculatingBooth_dup_1119)) ;
    nor02_2x L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix85 (.Y (
             L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_0), .A0 (nx7932), .A1 (
             nx3386)) ;
    inv01 ix3385 (.Y (nx3386), .A (L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_1)) ;
    mux21 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix125 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_1), .A0 (nx3388), .A1 (
          nx3390), .S0 (nx7932)) ;
    inv01 ix3387 (.Y (nx3388), .A (L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_2)) ;
    inv01 ix3389 (.Y (nx3390), .A (WindowDin_1__3__0)) ;
    mux21 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix133 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_2), .A0 (nx3392), .A1 (
          nx3394), .S0 (nx7932)) ;
    inv01 ix3391 (.Y (nx3392), .A (L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_3)) ;
    inv01 ix3393 (.Y (nx3394), .A (WindowDin_1__3__1)) ;
    mux21 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix141 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_3), .A0 (nx3396), .A1 (
          nx3398), .S0 (nx7932)) ;
    inv01 ix3395 (.Y (nx3396), .A (L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_4)) ;
    inv01 ix3397 (.Y (nx3398), .A (WindowDin_1__3__2)) ;
    mux21 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix149 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_4), .A0 (nx3400), .A1 (
          nx3402), .S0 (nx7932)) ;
    inv01 ix3399 (.Y (nx3400), .A (L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_5)) ;
    inv01 ix3401 (.Y (nx3402), .A (WindowDin_1__3__3)) ;
    mux21 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix157 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_5), .A0 (nx3404), .A1 (
          nx3406), .S0 (nx7932)) ;
    inv01 ix3403 (.Y (nx3404), .A (L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_6)) ;
    inv01 ix3405 (.Y (nx3406), .A (WindowDin_1__3__4)) ;
    mux21 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix165 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_6), .A0 (nx3408), .A1 (
          nx3410), .S0 (nx7932)) ;
    inv01 ix3407 (.Y (nx3408), .A (L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_7)) ;
    inv01 ix3409 (.Y (nx3410), .A (WindowDin_1__3__5)) ;
    mux21 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix173 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_7), .A0 (nx3412), .A1 (
          nx3414), .S0 (nx7934)) ;
    inv01 ix3411 (.Y (nx3412), .A (L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_8)) ;
    inv01 ix3413 (.Y (nx3414), .A (WindowDin_1__3__6)) ;
    mux21 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix181 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_8), .A0 (nx3416), .A1 (
          nx3418), .S0 (nx7934)) ;
    inv01 ix3415 (.Y (nx3416), .A (L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_9)) ;
    inv01 ix3417 (.Y (nx3418), .A (WindowDin_1__3__7)) ;
    nor02_2x L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix89 (.Y (
             L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_9), .A0 (nx7934), .A1 (
             nx3420)) ;
    inv01 ix3419 (.Y (nx3420), .A (L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_10)
          ) ;
    nor02_2x L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix93 (.Y (
             L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_10), .A0 (nx7934), .A1 (
             nx3422)) ;
    inv01 ix3421 (.Y (nx3422), .A (L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_11)
          ) ;
    nor02_2x L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix97 (.Y (
             L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_11), .A0 (nx7934), .A1 (
             nx3424)) ;
    inv01 ix3423 (.Y (nx3424), .A (L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_12)
          ) ;
    nor02_2x L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix101 (.Y (
             L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_12), .A0 (nx7934), .A1 (
             nx3426)) ;
    inv01 ix3425 (.Y (nx3426), .A (L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_13)
          ) ;
    nor02_2x L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix105 (.Y (
             L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_13), .A0 (nx7934), .A1 (
             nx3428)) ;
    inv01 ix3427 (.Y (nx3428), .A (L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_14)
          ) ;
    nor02_2x L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix109 (.Y (
             L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_14), .A0 (nx7936), .A1 (
             nx3430)) ;
    inv01 ix3429 (.Y (nx3430), .A (L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_15)
          ) ;
    nor02_2x L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix113 (.Y (
             L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_15), .A0 (nx7936), .A1 (
             nx3432)) ;
    inv01 ix3431 (.Y (nx3432), .A (L1_1_L2_3_G1_MINI_ALU_BoothPBeforeShift_16)
          ) ;
    nor02_2x L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix117 (.Y (
             L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_16), .A0 (nx7936), .A1 (
             nx3432)) ;
    mux21 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix189 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BoothOperand_0), .A0 (nx3434), .A1 (nx3436), .S0 (
          nx7924)) ;
    inv01 ix3433 (.Y (nx3434), .A (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_0)) ;
    inv01 ix3435 (.Y (nx3436), .A (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_0)) ;
    mux21 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix197 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BoothOperand_1), .A0 (nx3438), .A1 (nx3440), .S0 (
          nx7924)) ;
    inv01 ix3437 (.Y (nx3438), .A (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_1)) ;
    inv01 ix3439 (.Y (nx3440), .A (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_1)) ;
    mux21 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix205 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BoothOperand_2), .A0 (nx3442), .A1 (nx3444), .S0 (
          nx7924)) ;
    inv01 ix3441 (.Y (nx3442), .A (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_2)) ;
    inv01 ix3443 (.Y (nx3444), .A (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_2)) ;
    mux21 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix213 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BoothOperand_3), .A0 (nx3446), .A1 (nx3448), .S0 (
          nx7924)) ;
    inv01 ix3445 (.Y (nx3446), .A (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_3)) ;
    inv01 ix3447 (.Y (nx3448), .A (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_3)) ;
    mux21 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix221 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BoothOperand_4), .A0 (nx3450), .A1 (nx3452), .S0 (
          nx7924)) ;
    inv01 ix3449 (.Y (nx3450), .A (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_4)) ;
    inv01 ix3451 (.Y (nx3452), .A (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_4)) ;
    mux21 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix229 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BoothOperand_5), .A0 (nx3454), .A1 (nx3456), .S0 (
          nx7926)) ;
    inv01 ix3453 (.Y (nx3454), .A (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_5)) ;
    inv01 ix3455 (.Y (nx3456), .A (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_5)) ;
    mux21 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix237 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BoothOperand_6), .A0 (nx3458), .A1 (nx3460), .S0 (
          nx7926)) ;
    inv01 ix3457 (.Y (nx3458), .A (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_6)) ;
    inv01 ix3459 (.Y (nx3460), .A (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_6)) ;
    mux21 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix245 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BoothOperand_7), .A0 (nx3462), .A1 (nx3464), .S0 (
          nx7926)) ;
    inv01 ix3461 (.Y (nx3462), .A (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_7)) ;
    inv01 ix3463 (.Y (nx3464), .A (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_7)) ;
    mux21 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix253 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BoothOperand_8), .A0 (nx3466), .A1 (nx3468), .S0 (
          nx7926)) ;
    inv01 ix3465 (.Y (nx3466), .A (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_8)) ;
    inv01 ix3467 (.Y (nx3468), .A (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_8)) ;
    mux21 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix261 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BoothOperand_9), .A0 (nx3470), .A1 (nx3472), .S0 (
          nx7926)) ;
    inv01 ix3469 (.Y (nx3470), .A (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_9)) ;
    inv01 ix3471 (.Y (nx3472), .A (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_9)) ;
    mux21 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix269 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BoothOperand_10), .A0 (nx3474), .A1 (nx3476), .S0 (
          nx7926)) ;
    inv01 ix3473 (.Y (nx3474), .A (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_10)) ;
    inv01 ix3475 (.Y (nx3476), .A (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_10)) ;
    mux21 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix277 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BoothOperand_11), .A0 (nx3478), .A1 (nx3480), .S0 (
          nx7926)) ;
    inv01 ix3477 (.Y (nx3478), .A (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_11)) ;
    inv01 ix3479 (.Y (nx3480), .A (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_11)) ;
    mux21 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix285 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BoothOperand_12), .A0 (nx3482), .A1 (nx3484), .S0 (
          nx7928)) ;
    inv01 ix3481 (.Y (nx3482), .A (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_12)) ;
    inv01 ix3483 (.Y (nx3484), .A (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_12)) ;
    mux21 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix293 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BoothOperand_13), .A0 (nx3486), .A1 (nx3488), .S0 (
          nx7928)) ;
    inv01 ix3485 (.Y (nx3486), .A (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_13)) ;
    inv01 ix3487 (.Y (nx3488), .A (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_13)) ;
    mux21 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix301 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BoothOperand_14), .A0 (nx3490), .A1 (nx3492), .S0 (
          nx7928)) ;
    inv01 ix3489 (.Y (nx3490), .A (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_14)) ;
    inv01 ix3491 (.Y (nx3492), .A (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_14)) ;
    mux21 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix309 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BoothOperand_15), .A0 (nx3494), .A1 (nx3496), .S0 (
          nx7928)) ;
    inv01 ix3493 (.Y (nx3494), .A (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_15)) ;
    inv01 ix3495 (.Y (nx3496), .A (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_15)) ;
    mux21 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix317 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BoothOperand_16), .A0 (nx3498), .A1 (nx3500), .S0 (
          nx7928)) ;
    inv01 ix3497 (.Y (nx3498), .A (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_16)) ;
    inv01 ix3499 (.Y (nx3500), .A (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_16)) ;
    xnor2 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_ix321 (.Y (
          L1_1_L2_3_G1_MINI_ALU_AddPToBoothOperand), .A0 (nx7928), .A1 (nx3366)
          ) ;
    oai32 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix393 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .A0 (nx8644), .A1 (
          RST), .A2 (nx7938), .B0 (nx3436), .B1 (nx3504)) ;
    oai32 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix403 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .A0 (nx8644), .A1 (
          RST), .A2 (nx7938), .B0 (nx3440), .B1 (nx3504)) ;
    oai32 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix413 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .A0 (nx8644), .A1 (
          RST), .A2 (nx7938), .B0 (nx3444), .B1 (nx3504)) ;
    oai32 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix423 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .A0 (nx8644), .A1 (
          RST), .A2 (nx7938), .B0 (nx3448), .B1 (nx3504)) ;
    oai32 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix433 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .A0 (nx8644), .A1 (
          RST), .A2 (nx7938), .B0 (nx3452), .B1 (nx3504)) ;
    oai32 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix443 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .A0 (nx8644), .A1 (
          RST), .A2 (nx7938), .B0 (nx3456), .B1 (nx3504)) ;
    oai32 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix453 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .A0 (nx8644), .A1 (
          RST), .A2 (nx7940), .B0 (nx3460), .B1 (nx3504)) ;
    oai32 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix463 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .A0 (nx8646), .A1 (
          RST), .A2 (nx7940), .B0 (nx3464), .B1 (nx3506)) ;
    oai32 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix473 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .A0 (nx8646), .A1 (
          RST), .A2 (nx7940), .B0 (nx3468), .B1 (nx3506)) ;
    oai32 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix483 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .A0 (nx3508), .A1 (
          RST), .A2 (nx7940), .B0 (nx3472), .B1 (nx3506)) ;
    inv01 ix3507 (.Y (nx3508), .A (FilterDin_1__3__0)) ;
    oai32 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix493 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .A0 (nx3510), .A1 (
          RST), .A2 (nx7940), .B0 (nx3476), .B1 (nx3506)) ;
    inv01 ix3509 (.Y (nx3510), .A (FilterDin_1__3__1)) ;
    oai32 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix503 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .A0 (nx3512), .A1 (
          RST), .A2 (nx7940), .B0 (nx3480), .B1 (nx3506)) ;
    inv01 ix3511 (.Y (nx3512), .A (FilterDin_1__3__2)) ;
    oai32 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix513 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .A0 (nx3514), .A1 (
          RST), .A2 (nx7940), .B0 (nx3484), .B1 (nx3506)) ;
    inv01 ix3513 (.Y (nx3514), .A (FilterDin_1__3__3)) ;
    oai32 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix523 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .A0 (nx3516), .A1 (
          RST), .A2 (nx7942), .B0 (nx3488), .B1 (nx3506)) ;
    inv01 ix3515 (.Y (nx3516), .A (FilterDin_1__3__4)) ;
    oai32 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix533 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .A0 (nx3518), .A1 (
          RST), .A2 (nx7942), .B0 (nx3492), .B1 (nx3520)) ;
    inv01 ix3517 (.Y (nx3518), .A (FilterDin_1__3__5)) ;
    inv01 ix3519 (.Y (nx3520), .A (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566)) ;
    oai32 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix543 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .A0 (nx3522), .A1 (
          RST), .A2 (nx7942), .B0 (nx3496), .B1 (nx3520)) ;
    inv01 ix3521 (.Y (nx3522), .A (FilterDin_1__3__6)) ;
    oai32 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix553 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .A0 (nx3524), .A1 (
          RST), .A2 (nx7942), .B0 (nx3500), .B1 (nx3520)) ;
    inv01 ix3523 (.Y (nx3524), .A (FilterDin_1__3__7)) ;
    nand02_2x L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix633 (.Y (nx3504), .A0 (
              nx7588), .A1 (nx7942)) ;
    nand02_2x L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix635 (.Y (nx3506), .A0 (
              nx7590), .A1 (nx7942)) ;
    oai32 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix393 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .A0 (nx8646), .A1 (
          RST), .A2 (nx7944), .B0 (nx3434), .B1 (nx3526)) ;
    oai32 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix403 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .A0 (nx8646), .A1 (
          RST), .A2 (nx7944), .B0 (nx3438), .B1 (nx3526)) ;
    oai32 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix413 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .A0 (nx8646), .A1 (
          RST), .A2 (nx7944), .B0 (nx3442), .B1 (nx3526)) ;
    oai32 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix423 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .A0 (nx8646), .A1 (
          RST), .A2 (nx7944), .B0 (nx3446), .B1 (nx3526)) ;
    oai32 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix433 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .A0 (nx8646), .A1 (
          RST), .A2 (nx7944), .B0 (nx3450), .B1 (nx3526)) ;
    oai32 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix443 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .A0 (nx8648), .A1 (
          RST), .A2 (nx7944), .B0 (nx3454), .B1 (nx3526)) ;
    oai32 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix453 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .A0 (nx8648), .A1 (
          RST), .A2 (nx7946), .B0 (nx3458), .B1 (nx3526)) ;
    oai32 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix463 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .A0 (nx8648), .A1 (
          RST), .A2 (nx7946), .B0 (nx3462), .B1 (nx3528)) ;
    oai32 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix473 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .A0 (nx8648), .A1 (
          RST), .A2 (nx7946), .B0 (nx3466), .B1 (nx3528)) ;
    oai32 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix483 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .A0 (nx3508), .A1 (
          RST), .A2 (nx7946), .B0 (nx3470), .B1 (nx3528)) ;
    oai32 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix493 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .A0 (nx3530), .A1 (
          RST), .A2 (nx7946), .B0 (nx3474), .B1 (nx3528)) ;
    inv01 ix3529 (.Y (nx3530), .A (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_10)) ;
    oai32 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix503 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .A0 (nx3532), .A1 (
          RST), .A2 (nx7946), .B0 (nx3478), .B1 (nx3528)) ;
    inv01 ix3531 (.Y (nx3532), .A (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_11)) ;
    oai32 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix513 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .A0 (nx3534), .A1 (
          RST), .A2 (nx7946), .B0 (nx3482), .B1 (nx3528)) ;
    inv01 ix3533 (.Y (nx3534), .A (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_12)) ;
    oai32 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix523 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .A0 (nx3536), .A1 (
          RST), .A2 (nx7948), .B0 (nx3486), .B1 (nx3528)) ;
    inv01 ix3535 (.Y (nx3536), .A (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_13)) ;
    oai32 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix533 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .A0 (nx3538), .A1 (
          RST), .A2 (nx7948), .B0 (nx3490), .B1 (nx3540)) ;
    inv01 ix3537 (.Y (nx3538), .A (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_14)) ;
    inv01 ix3539 (.Y (nx3540), .A (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566)) ;
    oai32 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix543 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .A0 (nx3542), .A1 (
          RST), .A2 (nx7948), .B0 (nx3494), .B1 (nx3540)) ;
    inv01 ix3541 (.Y (nx3542), .A (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_15)) ;
    oai32 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix553 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .A0 (nx3544), .A1 (
          RST), .A2 (nx7948), .B0 (nx3498), .B1 (nx3540)) ;
    inv01 ix3543 (.Y (nx3544), .A (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_16)) ;
    nand02_2x L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix633 (.Y (nx3526), .A0 (
              nx7590), .A1 (nx7948)) ;
    nand02_2x L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix635 (.Y (nx3528), .A0 (
              nx7590), .A1 (nx7948)) ;
    oai32 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix393 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .A0 (nx3546), .A1 (
          RST), .A2 (nx7950), .B0 (L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx384), .B1 (
          nx3548)) ;
    inv01 ix3545 (.Y (nx3546), .A (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_0)) ;
    oai32 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix403 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .A0 (nx3550), .A1 (
          RST), .A2 (nx7950), .B0 (nx3366), .B1 (nx3548)) ;
    inv01 ix3549 (.Y (nx3550), .A (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_1)) ;
    oai32 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix413 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .A0 (nx3552), .A1 (
          RST), .A2 (nx7950), .B0 (L1_1_L2_3_G1_MINI_ALU_nx387), .B1 (nx3548)) ;
    inv01 ix3551 (.Y (nx3552), .A (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_2)) ;
    oai32 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix423 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .A0 (nx3554), .A1 (
          RST), .A2 (nx7950), .B0 (L1_1_L2_3_G1_MINI_ALU_nx399), .B1 (nx3548)) ;
    inv01 ix3553 (.Y (nx3554), .A (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_3)) ;
    oai32 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix433 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .A0 (nx3556), .A1 (
          RST), .A2 (nx7950), .B0 (L1_1_L2_3_G1_MINI_ALU_nx409), .B1 (nx3548)) ;
    inv01 ix3555 (.Y (nx3556), .A (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_4)) ;
    oai32 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix443 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .A0 (nx3558), .A1 (
          RST), .A2 (nx7950), .B0 (L1_1_L2_3_G1_MINI_ALU_nx419), .B1 (nx3548)) ;
    inv01 ix3557 (.Y (nx3558), .A (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_5)) ;
    oai32 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix453 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .A0 (nx3560), .A1 (
          RST), .A2 (nx7950), .B0 (L1_1_L2_3_G1_MINI_ALU_nx429), .B1 (nx3548)) ;
    inv01 ix3559 (.Y (nx3560), .A (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_6)) ;
    oai32 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix463 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .A0 (nx3562), .A1 (
          RST), .A2 (nx7952), .B0 (L1_1_L2_3_G1_MINI_ALU_nx439), .B1 (nx3564)) ;
    inv01 ix3561 (.Y (nx3562), .A (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_7)) ;
    oai32 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix473 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .A0 (nx3566), .A1 (
          RST), .A2 (nx7952), .B0 (L1_1_L2_3_G1_MINI_ALU_nx449), .B1 (nx3564)) ;
    inv01 ix3565 (.Y (nx3566), .A (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_8)) ;
    oai32 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix483 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .A0 (nx3568), .A1 (
          RST), .A2 (nx7952), .B0 (L1_1_L2_3_G1_MINI_ALU_nx469), .B1 (nx3564)) ;
    inv01 ix3567 (.Y (nx3568), .A (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_9)) ;
    oai32 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix493 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .A0 (nx3570), .A1 (
          RST), .A2 (nx7952), .B0 (L1_1_L2_3_G1_MINI_ALU_nx477), .B1 (nx3564)) ;
    inv01 ix3569 (.Y (nx3570), .A (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_10)) ;
    oai32 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix503 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .A0 (nx3572), .A1 (
          RST), .A2 (nx7952), .B0 (L1_1_L2_3_G1_MINI_ALU_nx485), .B1 (nx3564)) ;
    inv01 ix3571 (.Y (nx3572), .A (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_11)) ;
    oai32 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix513 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .A0 (nx3574), .A1 (
          RST), .A2 (nx7952), .B0 (L1_1_L2_3_G1_MINI_ALU_nx493), .B1 (nx3564)) ;
    inv01 ix3573 (.Y (nx3574), .A (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_12)) ;
    oai32 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix523 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .A0 (nx3576), .A1 (
          RST), .A2 (nx7952), .B0 (L1_1_L2_3_G1_MINI_ALU_nx501), .B1 (nx3564)) ;
    inv01 ix3575 (.Y (nx3576), .A (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_13)) ;
    oai32 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix533 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .A0 (nx3578), .A1 (
          RST), .A2 (nx7954), .B0 (L1_1_L2_3_G1_MINI_ALU_nx509), .B1 (nx3580)) ;
    inv01 ix3577 (.Y (nx3578), .A (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_14)) ;
    inv01 ix3579 (.Y (nx3580), .A (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566)) ;
    oai32 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix543 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .A0 (nx3582), .A1 (
          RST), .A2 (nx7954), .B0 (L1_1_L2_3_G1_MINI_ALU_nx517), .B1 (nx3580)) ;
    inv01 ix3581 (.Y (nx3582), .A (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_15)) ;
    oai32 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix553 (.Y (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .A0 (nx3584), .A1 (
          RST), .A2 (nx7954), .B0 (nx3382), .B1 (nx3580)) ;
    inv01 ix3583 (.Y (nx3584), .A (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_16)) ;
    nand02_2x L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix633 (.Y (nx3548), .A0 (
              nx7590), .A1 (nx7954)) ;
    nand02_2x L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix635 (.Y (nx3564), .A0 (
              nx7590), .A1 (nx7954)) ;
    mux21 L1_1_L2_4_G1_MINI_ALU_ix404 (.Y (L1_1_L2_4_G1_MINI_ALU_nx403), .A0 (
          nx3586), .A1 (L1_1_L2_4_G1_MINI_ALU_BoothP_2), .S0 (
          L1_1_L2_4_G1_MINI_ALU_nx395)) ;
    inv01 ix3585 (.Y (nx3586), .A (L1_1_L2_4_G1_MINI_ALU_nx391)) ;
    mux21 L1_1_L2_4_G1_MINI_ALU_ix414 (.Y (L1_1_L2_4_G1_MINI_ALU_nx413), .A0 (
          nx3588), .A1 (L1_1_L2_4_G1_MINI_ALU_BoothP_3), .S0 (
          L1_1_L2_4_G1_MINI_ALU_nx405)) ;
    inv01 ix3587 (.Y (nx3588), .A (L1_1_L2_4_G1_MINI_ALU_nx403)) ;
    mux21 L1_1_L2_4_G1_MINI_ALU_ix424 (.Y (L1_1_L2_4_G1_MINI_ALU_nx423), .A0 (
          nx3590), .A1 (L1_1_L2_4_G1_MINI_ALU_BoothP_4), .S0 (
          L1_1_L2_4_G1_MINI_ALU_nx415)) ;
    inv01 ix3589 (.Y (nx3590), .A (L1_1_L2_4_G1_MINI_ALU_nx413)) ;
    mux21 L1_1_L2_4_G1_MINI_ALU_ix434 (.Y (L1_1_L2_4_G1_MINI_ALU_nx433), .A0 (
          nx3592), .A1 (L1_1_L2_4_G1_MINI_ALU_BoothP_5), .S0 (
          L1_1_L2_4_G1_MINI_ALU_nx425)) ;
    inv01 ix3591 (.Y (nx3592), .A (L1_1_L2_4_G1_MINI_ALU_nx423)) ;
    mux21 L1_1_L2_4_G1_MINI_ALU_ix444 (.Y (L1_1_L2_4_G1_MINI_ALU_nx443), .A0 (
          nx3594), .A1 (L1_1_L2_4_G1_MINI_ALU_BoothP_6), .S0 (
          L1_1_L2_4_G1_MINI_ALU_nx435)) ;
    inv01 ix3593 (.Y (nx3594), .A (L1_1_L2_4_G1_MINI_ALU_nx433)) ;
    mux21 L1_1_L2_4_G1_MINI_ALU_ix454 (.Y (L1_1_L2_4_G1_MINI_ALU_nx453), .A0 (
          nx3596), .A1 (L1_1_L2_4_G1_MINI_ALU_BoothP_7), .S0 (
          L1_1_L2_4_G1_MINI_ALU_nx445)) ;
    inv01 ix3595 (.Y (nx3596), .A (L1_1_L2_4_G1_MINI_ALU_nx443)) ;
    mux21 L1_1_L2_4_G1_MINI_ALU_ix462 (.Y (L1_1_L2_4_G1_MINI_ALU_nx461), .A0 (
          nx3598), .A1 (L1_1_L2_4_G1_MINI_ALU_BoothP_8), .S0 (
          L1_1_L2_4_G1_MINI_ALU_nx455)) ;
    inv01 ix3597 (.Y (nx3598), .A (L1_1_L2_4_G1_MINI_ALU_nx453)) ;
    mux21 L1_1_L2_4_G1_MINI_ALU_ix468 (.Y (L1_1_L2_4_G1_MINI_ALU_nx467), .A0 (
          nx3600), .A1 (L1_1_L2_4_G1_MINI_ALU_BoothP_9), .S0 (
          L1_1_L2_4_G1_MINI_ALU_nx463)) ;
    inv01 ix3599 (.Y (nx3600), .A (L1_1_L2_4_G1_MINI_ALU_nx461)) ;
    mux21 L1_1_L2_4_G1_MINI_ALU_ix476 (.Y (L1_1_L2_4_G1_MINI_ALU_nx475), .A0 (
          nx3602), .A1 (L1_1_L2_4_G1_MINI_ALU_BoothP_10), .S0 (
          L1_1_L2_4_G1_MINI_ALU_nx471)) ;
    inv01 ix3601 (.Y (nx3602), .A (L1_1_L2_4_G1_MINI_ALU_nx467)) ;
    mux21 L1_1_L2_4_G1_MINI_ALU_ix484 (.Y (L1_1_L2_4_G1_MINI_ALU_nx483), .A0 (
          nx3604), .A1 (L1_1_L2_4_G1_MINI_ALU_BoothP_11), .S0 (
          L1_1_L2_4_G1_MINI_ALU_nx479)) ;
    inv01 ix3603 (.Y (nx3604), .A (L1_1_L2_4_G1_MINI_ALU_nx475)) ;
    mux21 L1_1_L2_4_G1_MINI_ALU_ix492 (.Y (L1_1_L2_4_G1_MINI_ALU_nx491), .A0 (
          nx3606), .A1 (L1_1_L2_4_G1_MINI_ALU_BoothP_12), .S0 (
          L1_1_L2_4_G1_MINI_ALU_nx487)) ;
    inv01 ix3605 (.Y (nx3606), .A (L1_1_L2_4_G1_MINI_ALU_nx483)) ;
    mux21 L1_1_L2_4_G1_MINI_ALU_ix500 (.Y (L1_1_L2_4_G1_MINI_ALU_nx499), .A0 (
          nx3608), .A1 (L1_1_L2_4_G1_MINI_ALU_BoothP_13), .S0 (
          L1_1_L2_4_G1_MINI_ALU_nx495)) ;
    inv01 ix3607 (.Y (nx3608), .A (L1_1_L2_4_G1_MINI_ALU_nx491)) ;
    mux21 L1_1_L2_4_G1_MINI_ALU_ix508 (.Y (L1_1_L2_4_G1_MINI_ALU_nx507), .A0 (
          nx3610), .A1 (L1_1_L2_4_G1_MINI_ALU_BoothP_14), .S0 (
          L1_1_L2_4_G1_MINI_ALU_nx503)) ;
    inv01 ix3609 (.Y (nx3610), .A (L1_1_L2_4_G1_MINI_ALU_nx499)) ;
    mux21 L1_1_L2_4_G1_MINI_ALU_ix516 (.Y (L1_1_L2_4_G1_MINI_ALU_nx515), .A0 (
          nx3612), .A1 (L1_1_L2_4_G1_MINI_ALU_BoothP_15), .S0 (
          L1_1_L2_4_G1_MINI_ALU_nx511)) ;
    inv01 ix3611 (.Y (nx3612), .A (L1_1_L2_4_G1_MINI_ALU_nx507)) ;
    mux21 L1_1_L2_4_G1_MINI_ALU_ix161 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_1), .A0 (nx3614), .A1 (
          L1_1_L2_4_G1_MINI_ALU_nx379), .S0 (nx7958)) ;
    inv01 ix3613 (.Y (nx3614), .A (L1_1_L2_4_G1_MINI_ALU_BoothP_1)) ;
    mux21 L1_1_L2_4_G1_MINI_ALU_ix181 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_2), .A0 (
          L1_1_L2_4_G1_MINI_ALU_nx387), .A1 (L1_1_L2_4_G1_MINI_ALU_nx389), .S0 (
          nx7958)) ;
    mux21 L1_1_L2_4_G1_MINI_ALU_ix201 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_3), .A0 (
          L1_1_L2_4_G1_MINI_ALU_nx399), .A1 (L1_1_L2_4_G1_MINI_ALU_nx401), .S0 (
          nx7958)) ;
    mux21 L1_1_L2_4_G1_MINI_ALU_ix221 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_4), .A0 (
          L1_1_L2_4_G1_MINI_ALU_nx409), .A1 (L1_1_L2_4_G1_MINI_ALU_nx411), .S0 (
          nx7958)) ;
    mux21 L1_1_L2_4_G1_MINI_ALU_ix241 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_5), .A0 (
          L1_1_L2_4_G1_MINI_ALU_nx419), .A1 (L1_1_L2_4_G1_MINI_ALU_nx421), .S0 (
          nx7958)) ;
    mux21 L1_1_L2_4_G1_MINI_ALU_ix261 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_6), .A0 (
          L1_1_L2_4_G1_MINI_ALU_nx429), .A1 (L1_1_L2_4_G1_MINI_ALU_nx431), .S0 (
          nx7958)) ;
    mux21 L1_1_L2_4_G1_MINI_ALU_ix281 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_7), .A0 (
          L1_1_L2_4_G1_MINI_ALU_nx439), .A1 (L1_1_L2_4_G1_MINI_ALU_nx441), .S0 (
          nx7958)) ;
    mux21 L1_1_L2_4_G1_MINI_ALU_ix301 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_8), .A0 (
          L1_1_L2_4_G1_MINI_ALU_nx449), .A1 (L1_1_L2_4_G1_MINI_ALU_nx451), .S0 (
          nx7960)) ;
    mux21 L1_1_L2_4_G1_MINI_ALU_ix321 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_9), .A0 (
          L1_1_L2_4_G1_MINI_ALU_nx469), .A1 (nx3616), .S0 (nx7960)) ;
    inv01 ix3615 (.Y (nx3616), .A (L1_1_L2_4_G1_MINI_ALU_nx316)) ;
    mux21 L1_1_L2_4_G1_MINI_ALU_ix341 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_10), .A0 (
          L1_1_L2_4_G1_MINI_ALU_nx477), .A1 (nx3618), .S0 (nx7960)) ;
    inv01 ix3617 (.Y (nx3618), .A (L1_1_L2_4_G1_MINI_ALU_nx336)) ;
    mux21 L1_1_L2_4_G1_MINI_ALU_ix361 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_11), .A0 (
          L1_1_L2_4_G1_MINI_ALU_nx485), .A1 (nx3620), .S0 (nx7960)) ;
    inv01 ix3619 (.Y (nx3620), .A (L1_1_L2_4_G1_MINI_ALU_nx356)) ;
    mux21 L1_1_L2_4_G1_MINI_ALU_ix381 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_12), .A0 (
          L1_1_L2_4_G1_MINI_ALU_nx493), .A1 (nx3622), .S0 (nx7960)) ;
    inv01 ix3621 (.Y (nx3622), .A (L1_1_L2_4_G1_MINI_ALU_nx376)) ;
    mux21 L1_1_L2_4_G1_MINI_ALU_ix401 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_13), .A0 (
          L1_1_L2_4_G1_MINI_ALU_nx501), .A1 (nx3624), .S0 (nx7960)) ;
    inv01 ix3623 (.Y (nx3624), .A (L1_1_L2_4_G1_MINI_ALU_nx396)) ;
    mux21 L1_1_L2_4_G1_MINI_ALU_ix421 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_14), .A0 (
          L1_1_L2_4_G1_MINI_ALU_nx509), .A1 (nx3626), .S0 (nx7960)) ;
    inv01 ix3625 (.Y (nx3626), .A (L1_1_L2_4_G1_MINI_ALU_nx416)) ;
    mux21 L1_1_L2_4_G1_MINI_ALU_ix441 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_15), .A0 (
          L1_1_L2_4_G1_MINI_ALU_nx517), .A1 (nx3628), .S0 (nx7962)) ;
    inv01 ix3627 (.Y (nx3628), .A (L1_1_L2_4_G1_MINI_ALU_nx436)) ;
    mux21 L1_1_L2_4_G1_MINI_ALU_ix461 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_16), .A0 (nx3630), .A1 (nx3632
          ), .S0 (nx7962)) ;
    inv01 ix3629 (.Y (nx3630), .A (L1_1_L2_4_G1_MINI_ALU_BoothP_16)) ;
    inv01 ix3631 (.Y (nx3632), .A (L1_1_L2_4_G1_MINI_ALU_nx456)) ;
    nor02_2x L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix319 (.Y (
             L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642), .A0 (Start), .A1 (
             CalculatingBooth_dup_1119)) ;
    nor02_2x L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix85 (.Y (
             L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_0), .A0 (nx7972), .A1 (
             nx3634)) ;
    inv01 ix3633 (.Y (nx3634), .A (L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_1)) ;
    mux21 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix125 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_1), .A0 (nx3636), .A1 (
          nx3638), .S0 (nx7972)) ;
    inv01 ix3635 (.Y (nx3636), .A (L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_2)) ;
    inv01 ix3637 (.Y (nx3638), .A (WindowDin_1__4__0)) ;
    mux21 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix133 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_2), .A0 (nx3640), .A1 (
          nx3642), .S0 (nx7972)) ;
    inv01 ix3639 (.Y (nx3640), .A (L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_3)) ;
    inv01 ix3641 (.Y (nx3642), .A (WindowDin_1__4__1)) ;
    mux21 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix141 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_3), .A0 (nx3644), .A1 (
          nx3646), .S0 (nx7972)) ;
    inv01 ix3643 (.Y (nx3644), .A (L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_4)) ;
    inv01 ix3645 (.Y (nx3646), .A (WindowDin_1__4__2)) ;
    mux21 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix149 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_4), .A0 (nx3648), .A1 (
          nx3650), .S0 (nx7972)) ;
    inv01 ix3647 (.Y (nx3648), .A (L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_5)) ;
    inv01 ix3649 (.Y (nx3650), .A (WindowDin_1__4__3)) ;
    mux21 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix157 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_5), .A0 (nx3652), .A1 (
          nx3654), .S0 (nx7972)) ;
    inv01 ix3651 (.Y (nx3652), .A (L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_6)) ;
    inv01 ix3653 (.Y (nx3654), .A (WindowDin_1__4__4)) ;
    mux21 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix165 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_6), .A0 (nx3656), .A1 (
          nx3658), .S0 (nx7972)) ;
    inv01 ix3655 (.Y (nx3656), .A (L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_7)) ;
    inv01 ix3657 (.Y (nx3658), .A (WindowDin_1__4__5)) ;
    mux21 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix173 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_7), .A0 (nx3660), .A1 (
          nx3662), .S0 (nx7974)) ;
    inv01 ix3659 (.Y (nx3660), .A (L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_8)) ;
    inv01 ix3661 (.Y (nx3662), .A (WindowDin_1__4__6)) ;
    mux21 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix181 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_8), .A0 (nx3664), .A1 (
          nx3666), .S0 (nx7974)) ;
    inv01 ix3663 (.Y (nx3664), .A (L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_9)) ;
    inv01 ix3665 (.Y (nx3666), .A (WindowDin_1__4__7)) ;
    nor02_2x L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix89 (.Y (
             L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_9), .A0 (nx7974), .A1 (
             nx3668)) ;
    inv01 ix3667 (.Y (nx3668), .A (L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_10)
          ) ;
    nor02_2x L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix93 (.Y (
             L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_10), .A0 (nx7974), .A1 (
             nx3670)) ;
    inv01 ix3669 (.Y (nx3670), .A (L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_11)
          ) ;
    nor02_2x L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix97 (.Y (
             L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_11), .A0 (nx7974), .A1 (
             nx3672)) ;
    inv01 ix3671 (.Y (nx3672), .A (L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_12)
          ) ;
    nor02_2x L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix101 (.Y (
             L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_12), .A0 (nx7974), .A1 (
             nx3674)) ;
    inv01 ix3673 (.Y (nx3674), .A (L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_13)
          ) ;
    nor02_2x L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix105 (.Y (
             L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_13), .A0 (nx7974), .A1 (
             nx3676)) ;
    inv01 ix3675 (.Y (nx3676), .A (L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_14)
          ) ;
    nor02_2x L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix109 (.Y (
             L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_14), .A0 (nx7976), .A1 (
             nx3678)) ;
    inv01 ix3677 (.Y (nx3678), .A (L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_15)
          ) ;
    nor02_2x L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix113 (.Y (
             L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_15), .A0 (nx7976), .A1 (
             nx3680)) ;
    inv01 ix3679 (.Y (nx3680), .A (L1_1_L2_4_G1_MINI_ALU_BoothPBeforeShift_16)
          ) ;
    nor02_2x L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix117 (.Y (
             L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_16), .A0 (nx7976), .A1 (
             nx3680)) ;
    mux21 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix189 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BoothOperand_0), .A0 (nx3682), .A1 (nx3684), .S0 (
          nx7964)) ;
    inv01 ix3681 (.Y (nx3682), .A (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_0)) ;
    inv01 ix3683 (.Y (nx3684), .A (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_0)) ;
    mux21 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix197 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BoothOperand_1), .A0 (nx3686), .A1 (nx3688), .S0 (
          nx7964)) ;
    inv01 ix3685 (.Y (nx3686), .A (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_1)) ;
    inv01 ix3687 (.Y (nx3688), .A (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_1)) ;
    mux21 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix205 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BoothOperand_2), .A0 (nx3690), .A1 (nx3692), .S0 (
          nx7964)) ;
    inv01 ix3689 (.Y (nx3690), .A (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_2)) ;
    inv01 ix3691 (.Y (nx3692), .A (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_2)) ;
    mux21 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix213 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BoothOperand_3), .A0 (nx3694), .A1 (nx3696), .S0 (
          nx7964)) ;
    inv01 ix3693 (.Y (nx3694), .A (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_3)) ;
    inv01 ix3695 (.Y (nx3696), .A (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_3)) ;
    mux21 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix221 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BoothOperand_4), .A0 (nx3698), .A1 (nx3700), .S0 (
          nx7964)) ;
    inv01 ix3697 (.Y (nx3698), .A (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_4)) ;
    inv01 ix3699 (.Y (nx3700), .A (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_4)) ;
    mux21 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix229 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BoothOperand_5), .A0 (nx3702), .A1 (nx3704), .S0 (
          nx7966)) ;
    inv01 ix3701 (.Y (nx3702), .A (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_5)) ;
    inv01 ix3703 (.Y (nx3704), .A (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_5)) ;
    mux21 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix237 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BoothOperand_6), .A0 (nx3706), .A1 (nx3708), .S0 (
          nx7966)) ;
    inv01 ix3705 (.Y (nx3706), .A (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_6)) ;
    inv01 ix3707 (.Y (nx3708), .A (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_6)) ;
    mux21 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix245 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BoothOperand_7), .A0 (nx3710), .A1 (nx3712), .S0 (
          nx7966)) ;
    inv01 ix3709 (.Y (nx3710), .A (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_7)) ;
    inv01 ix3711 (.Y (nx3712), .A (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_7)) ;
    mux21 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix253 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BoothOperand_8), .A0 (nx3714), .A1 (nx3716), .S0 (
          nx7966)) ;
    inv01 ix3713 (.Y (nx3714), .A (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_8)) ;
    inv01 ix3715 (.Y (nx3716), .A (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_8)) ;
    mux21 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix261 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BoothOperand_9), .A0 (nx3718), .A1 (nx3720), .S0 (
          nx7966)) ;
    inv01 ix3717 (.Y (nx3718), .A (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_9)) ;
    inv01 ix3719 (.Y (nx3720), .A (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_9)) ;
    mux21 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix269 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BoothOperand_10), .A0 (nx3722), .A1 (nx3724), .S0 (
          nx7966)) ;
    inv01 ix3721 (.Y (nx3722), .A (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_10)) ;
    inv01 ix3723 (.Y (nx3724), .A (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_10)) ;
    mux21 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix277 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BoothOperand_11), .A0 (nx3726), .A1 (nx3728), .S0 (
          nx7966)) ;
    inv01 ix3725 (.Y (nx3726), .A (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_11)) ;
    inv01 ix3727 (.Y (nx3728), .A (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_11)) ;
    mux21 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix285 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BoothOperand_12), .A0 (nx3730), .A1 (nx3732), .S0 (
          nx7968)) ;
    inv01 ix3729 (.Y (nx3730), .A (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_12)) ;
    inv01 ix3731 (.Y (nx3732), .A (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_12)) ;
    mux21 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix293 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BoothOperand_13), .A0 (nx3734), .A1 (nx3736), .S0 (
          nx7968)) ;
    inv01 ix3733 (.Y (nx3734), .A (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_13)) ;
    inv01 ix3735 (.Y (nx3736), .A (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_13)) ;
    mux21 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix301 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BoothOperand_14), .A0 (nx3738), .A1 (nx3740), .S0 (
          nx7968)) ;
    inv01 ix3737 (.Y (nx3738), .A (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_14)) ;
    inv01 ix3739 (.Y (nx3740), .A (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_14)) ;
    mux21 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix309 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BoothOperand_15), .A0 (nx3742), .A1 (nx3744), .S0 (
          nx7968)) ;
    inv01 ix3741 (.Y (nx3742), .A (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_15)) ;
    inv01 ix3743 (.Y (nx3744), .A (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_15)) ;
    mux21 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix317 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BoothOperand_16), .A0 (nx3746), .A1 (nx3748), .S0 (
          nx7968)) ;
    inv01 ix3745 (.Y (nx3746), .A (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_16)) ;
    inv01 ix3747 (.Y (nx3748), .A (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_16)) ;
    xnor2 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_ix321 (.Y (
          L1_1_L2_4_G1_MINI_ALU_AddPToBoothOperand), .A0 (nx7968), .A1 (nx3614)
          ) ;
    oai32 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix393 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .A0 (nx8650), .A1 (
          RST), .A2 (nx7978), .B0 (nx3684), .B1 (nx3752)) ;
    oai32 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix403 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .A0 (nx8650), .A1 (
          RST), .A2 (nx7978), .B0 (nx3688), .B1 (nx3752)) ;
    oai32 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix413 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .A0 (nx8650), .A1 (
          RST), .A2 (nx7978), .B0 (nx3692), .B1 (nx3752)) ;
    oai32 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix423 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .A0 (nx8650), .A1 (
          RST), .A2 (nx7978), .B0 (nx3696), .B1 (nx3752)) ;
    oai32 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix433 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .A0 (nx8650), .A1 (
          RST), .A2 (nx7978), .B0 (nx3700), .B1 (nx3752)) ;
    oai32 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix443 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .A0 (nx8650), .A1 (
          RST), .A2 (nx7978), .B0 (nx3704), .B1 (nx3752)) ;
    oai32 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix453 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .A0 (nx8650), .A1 (
          RST), .A2 (nx7980), .B0 (nx3708), .B1 (nx3752)) ;
    oai32 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix463 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .A0 (nx8652), .A1 (
          RST), .A2 (nx7980), .B0 (nx3712), .B1 (nx3754)) ;
    oai32 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix473 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .A0 (nx8652), .A1 (
          RST), .A2 (nx7980), .B0 (nx3716), .B1 (nx3754)) ;
    oai32 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix483 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .A0 (nx3756), .A1 (
          RST), .A2 (nx7980), .B0 (nx3720), .B1 (nx3754)) ;
    inv01 ix3755 (.Y (nx3756), .A (FilterDin_1__4__0)) ;
    oai32 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix493 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .A0 (nx3758), .A1 (
          RST), .A2 (nx7980), .B0 (nx3724), .B1 (nx3754)) ;
    inv01 ix3757 (.Y (nx3758), .A (FilterDin_1__4__1)) ;
    oai32 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix503 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .A0 (nx3760), .A1 (
          RST), .A2 (nx7980), .B0 (nx3728), .B1 (nx3754)) ;
    inv01 ix3759 (.Y (nx3760), .A (FilterDin_1__4__2)) ;
    oai32 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix513 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .A0 (nx3762), .A1 (
          RST), .A2 (nx7980), .B0 (nx3732), .B1 (nx3754)) ;
    inv01 ix3761 (.Y (nx3762), .A (FilterDin_1__4__3)) ;
    oai32 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix523 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .A0 (nx3764), .A1 (
          RST), .A2 (nx7982), .B0 (nx3736), .B1 (nx3754)) ;
    inv01 ix3763 (.Y (nx3764), .A (FilterDin_1__4__4)) ;
    oai32 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix533 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .A0 (nx3766), .A1 (
          RST), .A2 (nx7982), .B0 (nx3740), .B1 (nx3768)) ;
    inv01 ix3765 (.Y (nx3766), .A (FilterDin_1__4__5)) ;
    inv01 ix3767 (.Y (nx3768), .A (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566)) ;
    oai32 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix543 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .A0 (nx3770), .A1 (
          RST), .A2 (nx7982), .B0 (nx3744), .B1 (nx3768)) ;
    inv01 ix3769 (.Y (nx3770), .A (FilterDin_1__4__6)) ;
    oai32 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix553 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .A0 (nx3772), .A1 (
          RST), .A2 (nx7982), .B0 (nx3748), .B1 (nx3768)) ;
    inv01 ix3771 (.Y (nx3772), .A (FilterDin_1__4__7)) ;
    nand02_2x L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix633 (.Y (nx3752), .A0 (
              nx7590), .A1 (nx7982)) ;
    nand02_2x L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix635 (.Y (nx3754), .A0 (
              nx7590), .A1 (nx7982)) ;
    oai32 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix393 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .A0 (nx8652), .A1 (
          RST), .A2 (nx7984), .B0 (nx3682), .B1 (nx3774)) ;
    oai32 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix403 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .A0 (nx8652), .A1 (
          RST), .A2 (nx7984), .B0 (nx3686), .B1 (nx3774)) ;
    oai32 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix413 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .A0 (nx8652), .A1 (
          RST), .A2 (nx7984), .B0 (nx3690), .B1 (nx3774)) ;
    oai32 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix423 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .A0 (nx8652), .A1 (
          RST), .A2 (nx7984), .B0 (nx3694), .B1 (nx3774)) ;
    oai32 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix433 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .A0 (nx8652), .A1 (
          RST), .A2 (nx7984), .B0 (nx3698), .B1 (nx3774)) ;
    oai32 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix443 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .A0 (nx8654), .A1 (
          RST), .A2 (nx7984), .B0 (nx3702), .B1 (nx3774)) ;
    oai32 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix453 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .A0 (nx8654), .A1 (
          RST), .A2 (nx7986), .B0 (nx3706), .B1 (nx3774)) ;
    oai32 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix463 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .A0 (nx8654), .A1 (
          RST), .A2 (nx7986), .B0 (nx3710), .B1 (nx3776)) ;
    oai32 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix473 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .A0 (nx8654), .A1 (
          RST), .A2 (nx7986), .B0 (nx3714), .B1 (nx3776)) ;
    oai32 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix483 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .A0 (nx3756), .A1 (
          RST), .A2 (nx7986), .B0 (nx3718), .B1 (nx3776)) ;
    oai32 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix493 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .A0 (nx3778), .A1 (
          RST), .A2 (nx7986), .B0 (nx3722), .B1 (nx3776)) ;
    inv01 ix3777 (.Y (nx3778), .A (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_10)) ;
    oai32 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix503 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .A0 (nx3780), .A1 (
          RST), .A2 (nx7986), .B0 (nx3726), .B1 (nx3776)) ;
    inv01 ix3779 (.Y (nx3780), .A (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_11)) ;
    oai32 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix513 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .A0 (nx3782), .A1 (
          RST), .A2 (nx7986), .B0 (nx3730), .B1 (nx3776)) ;
    inv01 ix3781 (.Y (nx3782), .A (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_12)) ;
    oai32 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix523 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .A0 (nx3784), .A1 (
          RST), .A2 (nx7988), .B0 (nx3734), .B1 (nx3776)) ;
    inv01 ix3783 (.Y (nx3784), .A (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_13)) ;
    oai32 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix533 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .A0 (nx3786), .A1 (
          RST), .A2 (nx7988), .B0 (nx3738), .B1 (nx3788)) ;
    inv01 ix3785 (.Y (nx3786), .A (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_14)) ;
    inv01 ix3787 (.Y (nx3788), .A (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566)) ;
    oai32 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix543 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .A0 (nx3790), .A1 (
          RST), .A2 (nx7988), .B0 (nx3742), .B1 (nx3788)) ;
    inv01 ix3789 (.Y (nx3790), .A (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_15)) ;
    oai32 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix553 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .A0 (nx3792), .A1 (
          RST), .A2 (nx7988), .B0 (nx3746), .B1 (nx3788)) ;
    inv01 ix3791 (.Y (nx3792), .A (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_16)) ;
    nand02_2x L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix633 (.Y (nx3774), .A0 (
              nx7592), .A1 (nx7988)) ;
    nand02_2x L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix635 (.Y (nx3776), .A0 (
              nx7592), .A1 (nx7988)) ;
    oai32 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix393 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .A0 (nx3794), .A1 (
          RST), .A2 (nx7990), .B0 (L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx384), .B1 (
          nx3796)) ;
    inv01 ix3793 (.Y (nx3794), .A (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_0)) ;
    oai32 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix403 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .A0 (nx3798), .A1 (
          RST), .A2 (nx7990), .B0 (nx3614), .B1 (nx3796)) ;
    inv01 ix3797 (.Y (nx3798), .A (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_1)) ;
    oai32 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix413 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .A0 (nx3800), .A1 (
          RST), .A2 (nx7990), .B0 (L1_1_L2_4_G1_MINI_ALU_nx387), .B1 (nx3796)) ;
    inv01 ix3799 (.Y (nx3800), .A (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_2)) ;
    oai32 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix423 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .A0 (nx3802), .A1 (
          RST), .A2 (nx7990), .B0 (L1_1_L2_4_G1_MINI_ALU_nx399), .B1 (nx3796)) ;
    inv01 ix3801 (.Y (nx3802), .A (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_3)) ;
    oai32 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix433 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .A0 (nx3804), .A1 (
          RST), .A2 (nx7990), .B0 (L1_1_L2_4_G1_MINI_ALU_nx409), .B1 (nx3796)) ;
    inv01 ix3803 (.Y (nx3804), .A (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_4)) ;
    oai32 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix443 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .A0 (nx3806), .A1 (
          RST), .A2 (nx7990), .B0 (L1_1_L2_4_G1_MINI_ALU_nx419), .B1 (nx3796)) ;
    inv01 ix3805 (.Y (nx3806), .A (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_5)) ;
    oai32 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix453 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .A0 (nx3808), .A1 (
          RST), .A2 (nx7990), .B0 (L1_1_L2_4_G1_MINI_ALU_nx429), .B1 (nx3796)) ;
    inv01 ix3807 (.Y (nx3808), .A (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_6)) ;
    oai32 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix463 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .A0 (nx3810), .A1 (
          RST), .A2 (nx7992), .B0 (L1_1_L2_4_G1_MINI_ALU_nx439), .B1 (nx3812)) ;
    inv01 ix3809 (.Y (nx3810), .A (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_7)) ;
    oai32 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix473 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .A0 (nx3814), .A1 (
          RST), .A2 (nx7992), .B0 (L1_1_L2_4_G1_MINI_ALU_nx449), .B1 (nx3812)) ;
    inv01 ix3813 (.Y (nx3814), .A (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_8)) ;
    oai32 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix483 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .A0 (nx3816), .A1 (
          RST), .A2 (nx7992), .B0 (L1_1_L2_4_G1_MINI_ALU_nx469), .B1 (nx3812)) ;
    inv01 ix3815 (.Y (nx3816), .A (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_9)) ;
    oai32 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix493 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .A0 (nx3818), .A1 (
          RST), .A2 (nx7992), .B0 (L1_1_L2_4_G1_MINI_ALU_nx477), .B1 (nx3812)) ;
    inv01 ix3817 (.Y (nx3818), .A (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_10)) ;
    oai32 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix503 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .A0 (nx3820), .A1 (
          RST), .A2 (nx7992), .B0 (L1_1_L2_4_G1_MINI_ALU_nx485), .B1 (nx3812)) ;
    inv01 ix3819 (.Y (nx3820), .A (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_11)) ;
    oai32 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix513 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .A0 (nx3822), .A1 (
          RST), .A2 (nx7992), .B0 (L1_1_L2_4_G1_MINI_ALU_nx493), .B1 (nx3812)) ;
    inv01 ix3821 (.Y (nx3822), .A (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_12)) ;
    oai32 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix523 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .A0 (nx3824), .A1 (
          RST), .A2 (nx7992), .B0 (L1_1_L2_4_G1_MINI_ALU_nx501), .B1 (nx3812)) ;
    inv01 ix3823 (.Y (nx3824), .A (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_13)) ;
    oai32 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix533 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .A0 (nx3826), .A1 (
          RST), .A2 (nx7994), .B0 (L1_1_L2_4_G1_MINI_ALU_nx509), .B1 (nx3828)) ;
    inv01 ix3825 (.Y (nx3826), .A (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_14)) ;
    inv01 ix3827 (.Y (nx3828), .A (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566)) ;
    oai32 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix543 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .A0 (nx3830), .A1 (
          RST), .A2 (nx7994), .B0 (L1_1_L2_4_G1_MINI_ALU_nx517), .B1 (nx3828)) ;
    inv01 ix3829 (.Y (nx3830), .A (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_15)) ;
    oai32 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix553 (.Y (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .A0 (nx3832), .A1 (
          RST), .A2 (nx7994), .B0 (nx3630), .B1 (nx3828)) ;
    inv01 ix3831 (.Y (nx3832), .A (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_16)) ;
    nand02_2x L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix633 (.Y (nx3796), .A0 (
              nx7592), .A1 (nx7994)) ;
    nand02_2x L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix635 (.Y (nx3812), .A0 (
              nx7592), .A1 (nx7994)) ;
    mux21 L1_2_L2_0_G1_MINI_ALU_ix404 (.Y (L1_2_L2_0_G1_MINI_ALU_nx403), .A0 (
          nx3834), .A1 (L1_2_L2_0_G1_MINI_ALU_BoothP_2), .S0 (
          L1_2_L2_0_G1_MINI_ALU_nx395)) ;
    inv01 ix3833 (.Y (nx3834), .A (L1_2_L2_0_G1_MINI_ALU_nx391)) ;
    mux21 L1_2_L2_0_G1_MINI_ALU_ix414 (.Y (L1_2_L2_0_G1_MINI_ALU_nx413), .A0 (
          nx3836), .A1 (L1_2_L2_0_G1_MINI_ALU_BoothP_3), .S0 (
          L1_2_L2_0_G1_MINI_ALU_nx405)) ;
    inv01 ix3835 (.Y (nx3836), .A (L1_2_L2_0_G1_MINI_ALU_nx403)) ;
    mux21 L1_2_L2_0_G1_MINI_ALU_ix424 (.Y (L1_2_L2_0_G1_MINI_ALU_nx423), .A0 (
          nx3838), .A1 (L1_2_L2_0_G1_MINI_ALU_BoothP_4), .S0 (
          L1_2_L2_0_G1_MINI_ALU_nx415)) ;
    inv01 ix3837 (.Y (nx3838), .A (L1_2_L2_0_G1_MINI_ALU_nx413)) ;
    mux21 L1_2_L2_0_G1_MINI_ALU_ix434 (.Y (L1_2_L2_0_G1_MINI_ALU_nx433), .A0 (
          nx3840), .A1 (L1_2_L2_0_G1_MINI_ALU_BoothP_5), .S0 (
          L1_2_L2_0_G1_MINI_ALU_nx425)) ;
    inv01 ix3839 (.Y (nx3840), .A (L1_2_L2_0_G1_MINI_ALU_nx423)) ;
    mux21 L1_2_L2_0_G1_MINI_ALU_ix444 (.Y (L1_2_L2_0_G1_MINI_ALU_nx443), .A0 (
          nx3842), .A1 (L1_2_L2_0_G1_MINI_ALU_BoothP_6), .S0 (
          L1_2_L2_0_G1_MINI_ALU_nx435)) ;
    inv01 ix3841 (.Y (nx3842), .A (L1_2_L2_0_G1_MINI_ALU_nx433)) ;
    mux21 L1_2_L2_0_G1_MINI_ALU_ix454 (.Y (L1_2_L2_0_G1_MINI_ALU_nx453), .A0 (
          nx3844), .A1 (L1_2_L2_0_G1_MINI_ALU_BoothP_7), .S0 (
          L1_2_L2_0_G1_MINI_ALU_nx445)) ;
    inv01 ix3843 (.Y (nx3844), .A (L1_2_L2_0_G1_MINI_ALU_nx443)) ;
    mux21 L1_2_L2_0_G1_MINI_ALU_ix462 (.Y (L1_2_L2_0_G1_MINI_ALU_nx461), .A0 (
          nx3846), .A1 (L1_2_L2_0_G1_MINI_ALU_BoothP_8), .S0 (
          L1_2_L2_0_G1_MINI_ALU_nx455)) ;
    inv01 ix3845 (.Y (nx3846), .A (L1_2_L2_0_G1_MINI_ALU_nx453)) ;
    mux21 L1_2_L2_0_G1_MINI_ALU_ix468 (.Y (L1_2_L2_0_G1_MINI_ALU_nx467), .A0 (
          nx3848), .A1 (L1_2_L2_0_G1_MINI_ALU_BoothP_9), .S0 (
          L1_2_L2_0_G1_MINI_ALU_nx463)) ;
    inv01 ix3847 (.Y (nx3848), .A (L1_2_L2_0_G1_MINI_ALU_nx461)) ;
    mux21 L1_2_L2_0_G1_MINI_ALU_ix476 (.Y (L1_2_L2_0_G1_MINI_ALU_nx475), .A0 (
          nx3850), .A1 (L1_2_L2_0_G1_MINI_ALU_BoothP_10), .S0 (
          L1_2_L2_0_G1_MINI_ALU_nx471)) ;
    inv01 ix3849 (.Y (nx3850), .A (L1_2_L2_0_G1_MINI_ALU_nx467)) ;
    mux21 L1_2_L2_0_G1_MINI_ALU_ix484 (.Y (L1_2_L2_0_G1_MINI_ALU_nx483), .A0 (
          nx3852), .A1 (L1_2_L2_0_G1_MINI_ALU_BoothP_11), .S0 (
          L1_2_L2_0_G1_MINI_ALU_nx479)) ;
    inv01 ix3851 (.Y (nx3852), .A (L1_2_L2_0_G1_MINI_ALU_nx475)) ;
    mux21 L1_2_L2_0_G1_MINI_ALU_ix492 (.Y (L1_2_L2_0_G1_MINI_ALU_nx491), .A0 (
          nx3854), .A1 (L1_2_L2_0_G1_MINI_ALU_BoothP_12), .S0 (
          L1_2_L2_0_G1_MINI_ALU_nx487)) ;
    inv01 ix3853 (.Y (nx3854), .A (L1_2_L2_0_G1_MINI_ALU_nx483)) ;
    mux21 L1_2_L2_0_G1_MINI_ALU_ix500 (.Y (L1_2_L2_0_G1_MINI_ALU_nx499), .A0 (
          nx3856), .A1 (L1_2_L2_0_G1_MINI_ALU_BoothP_13), .S0 (
          L1_2_L2_0_G1_MINI_ALU_nx495)) ;
    inv01 ix3855 (.Y (nx3856), .A (L1_2_L2_0_G1_MINI_ALU_nx491)) ;
    mux21 L1_2_L2_0_G1_MINI_ALU_ix508 (.Y (L1_2_L2_0_G1_MINI_ALU_nx507), .A0 (
          nx3858), .A1 (L1_2_L2_0_G1_MINI_ALU_BoothP_14), .S0 (
          L1_2_L2_0_G1_MINI_ALU_nx503)) ;
    inv01 ix3857 (.Y (nx3858), .A (L1_2_L2_0_G1_MINI_ALU_nx499)) ;
    mux21 L1_2_L2_0_G1_MINI_ALU_ix516 (.Y (L1_2_L2_0_G1_MINI_ALU_nx515), .A0 (
          nx3860), .A1 (L1_2_L2_0_G1_MINI_ALU_BoothP_15), .S0 (
          L1_2_L2_0_G1_MINI_ALU_nx511)) ;
    inv01 ix3859 (.Y (nx3860), .A (L1_2_L2_0_G1_MINI_ALU_nx507)) ;
    mux21 L1_2_L2_0_G1_MINI_ALU_ix161 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_1), .A0 (nx3862), .A1 (
          L1_2_L2_0_G1_MINI_ALU_nx379), .S0 (nx7998)) ;
    inv01 ix3861 (.Y (nx3862), .A (L1_2_L2_0_G1_MINI_ALU_BoothP_1)) ;
    mux21 L1_2_L2_0_G1_MINI_ALU_ix181 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_2), .A0 (
          L1_2_L2_0_G1_MINI_ALU_nx387), .A1 (L1_2_L2_0_G1_MINI_ALU_nx389), .S0 (
          nx7998)) ;
    mux21 L1_2_L2_0_G1_MINI_ALU_ix201 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_3), .A0 (
          L1_2_L2_0_G1_MINI_ALU_nx399), .A1 (L1_2_L2_0_G1_MINI_ALU_nx401), .S0 (
          nx7998)) ;
    mux21 L1_2_L2_0_G1_MINI_ALU_ix221 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_4), .A0 (
          L1_2_L2_0_G1_MINI_ALU_nx409), .A1 (L1_2_L2_0_G1_MINI_ALU_nx411), .S0 (
          nx7998)) ;
    mux21 L1_2_L2_0_G1_MINI_ALU_ix241 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_5), .A0 (
          L1_2_L2_0_G1_MINI_ALU_nx419), .A1 (L1_2_L2_0_G1_MINI_ALU_nx421), .S0 (
          nx7998)) ;
    mux21 L1_2_L2_0_G1_MINI_ALU_ix261 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_6), .A0 (
          L1_2_L2_0_G1_MINI_ALU_nx429), .A1 (L1_2_L2_0_G1_MINI_ALU_nx431), .S0 (
          nx7998)) ;
    mux21 L1_2_L2_0_G1_MINI_ALU_ix281 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_7), .A0 (
          L1_2_L2_0_G1_MINI_ALU_nx439), .A1 (L1_2_L2_0_G1_MINI_ALU_nx441), .S0 (
          nx7998)) ;
    mux21 L1_2_L2_0_G1_MINI_ALU_ix301 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_8), .A0 (
          L1_2_L2_0_G1_MINI_ALU_nx449), .A1 (L1_2_L2_0_G1_MINI_ALU_nx451), .S0 (
          nx8000)) ;
    mux21 L1_2_L2_0_G1_MINI_ALU_ix321 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_9), .A0 (
          L1_2_L2_0_G1_MINI_ALU_nx469), .A1 (nx3864), .S0 (nx8000)) ;
    inv01 ix3863 (.Y (nx3864), .A (L1_2_L2_0_G1_MINI_ALU_nx316)) ;
    mux21 L1_2_L2_0_G1_MINI_ALU_ix341 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_10), .A0 (
          L1_2_L2_0_G1_MINI_ALU_nx477), .A1 (nx3866), .S0 (nx8000)) ;
    inv01 ix3865 (.Y (nx3866), .A (L1_2_L2_0_G1_MINI_ALU_nx336)) ;
    mux21 L1_2_L2_0_G1_MINI_ALU_ix361 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_11), .A0 (
          L1_2_L2_0_G1_MINI_ALU_nx485), .A1 (nx3868), .S0 (nx8000)) ;
    inv01 ix3867 (.Y (nx3868), .A (L1_2_L2_0_G1_MINI_ALU_nx356)) ;
    mux21 L1_2_L2_0_G1_MINI_ALU_ix381 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_12), .A0 (
          L1_2_L2_0_G1_MINI_ALU_nx493), .A1 (nx3870), .S0 (nx8000)) ;
    inv01 ix3869 (.Y (nx3870), .A (L1_2_L2_0_G1_MINI_ALU_nx376)) ;
    mux21 L1_2_L2_0_G1_MINI_ALU_ix401 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_13), .A0 (
          L1_2_L2_0_G1_MINI_ALU_nx501), .A1 (nx3872), .S0 (nx8000)) ;
    inv01 ix3871 (.Y (nx3872), .A (L1_2_L2_0_G1_MINI_ALU_nx396)) ;
    mux21 L1_2_L2_0_G1_MINI_ALU_ix421 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_14), .A0 (
          L1_2_L2_0_G1_MINI_ALU_nx509), .A1 (nx3874), .S0 (nx8000)) ;
    inv01 ix3873 (.Y (nx3874), .A (L1_2_L2_0_G1_MINI_ALU_nx416)) ;
    mux21 L1_2_L2_0_G1_MINI_ALU_ix441 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_15), .A0 (
          L1_2_L2_0_G1_MINI_ALU_nx517), .A1 (nx3876), .S0 (nx8002)) ;
    inv01 ix3875 (.Y (nx3876), .A (L1_2_L2_0_G1_MINI_ALU_nx436)) ;
    mux21 L1_2_L2_0_G1_MINI_ALU_ix461 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_16), .A0 (nx3878), .A1 (nx3880
          ), .S0 (nx8002)) ;
    inv01 ix3877 (.Y (nx3878), .A (L1_2_L2_0_G1_MINI_ALU_BoothP_16)) ;
    inv01 ix3879 (.Y (nx3880), .A (L1_2_L2_0_G1_MINI_ALU_nx456)) ;
    nor02_2x L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix319 (.Y (
             L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642), .A0 (Start), .A1 (
             CalculatingBooth_dup_1119)) ;
    nor02_2x L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix85 (.Y (
             L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_0), .A0 (nx8012), .A1 (
             nx3882)) ;
    inv01 ix3881 (.Y (nx3882), .A (L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_1)) ;
    mux21 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix125 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_1), .A0 (nx3884), .A1 (
          nx3886), .S0 (nx8012)) ;
    inv01 ix3883 (.Y (nx3884), .A (L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_2)) ;
    inv01 ix3885 (.Y (nx3886), .A (WindowDin_2__0__0)) ;
    mux21 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix133 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_2), .A0 (nx3888), .A1 (
          nx3890), .S0 (nx8012)) ;
    inv01 ix3887 (.Y (nx3888), .A (L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_3)) ;
    inv01 ix3889 (.Y (nx3890), .A (WindowDin_2__0__1)) ;
    mux21 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix141 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_3), .A0 (nx3892), .A1 (
          nx3894), .S0 (nx8012)) ;
    inv01 ix3891 (.Y (nx3892), .A (L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_4)) ;
    inv01 ix3893 (.Y (nx3894), .A (WindowDin_2__0__2)) ;
    mux21 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix149 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_4), .A0 (nx3896), .A1 (
          nx3898), .S0 (nx8012)) ;
    inv01 ix3895 (.Y (nx3896), .A (L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_5)) ;
    inv01 ix3897 (.Y (nx3898), .A (WindowDin_2__0__3)) ;
    mux21 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix157 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_5), .A0 (nx3900), .A1 (
          nx3902), .S0 (nx8012)) ;
    inv01 ix3899 (.Y (nx3900), .A (L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_6)) ;
    inv01 ix3901 (.Y (nx3902), .A (WindowDin_2__0__4)) ;
    mux21 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix165 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_6), .A0 (nx3904), .A1 (
          nx3906), .S0 (nx8012)) ;
    inv01 ix3903 (.Y (nx3904), .A (L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_7)) ;
    inv01 ix3905 (.Y (nx3906), .A (WindowDin_2__0__5)) ;
    mux21 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix173 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_7), .A0 (nx3908), .A1 (
          nx3910), .S0 (nx8014)) ;
    inv01 ix3907 (.Y (nx3908), .A (L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_8)) ;
    inv01 ix3909 (.Y (nx3910), .A (WindowDin_2__0__6)) ;
    mux21 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix181 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_8), .A0 (nx3912), .A1 (
          nx3914), .S0 (nx8014)) ;
    inv01 ix3911 (.Y (nx3912), .A (L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_9)) ;
    inv01 ix3913 (.Y (nx3914), .A (WindowDin_2__0__7)) ;
    nor02_2x L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix89 (.Y (
             L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_9), .A0 (nx8014), .A1 (
             nx3916)) ;
    inv01 ix3915 (.Y (nx3916), .A (L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_10)
          ) ;
    nor02_2x L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix93 (.Y (
             L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_10), .A0 (nx8014), .A1 (
             nx3918)) ;
    inv01 ix3917 (.Y (nx3918), .A (L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_11)
          ) ;
    nor02_2x L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix97 (.Y (
             L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_11), .A0 (nx8014), .A1 (
             nx3920)) ;
    inv01 ix3919 (.Y (nx3920), .A (L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_12)
          ) ;
    nor02_2x L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix101 (.Y (
             L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_12), .A0 (nx8014), .A1 (
             nx3922)) ;
    inv01 ix3921 (.Y (nx3922), .A (L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_13)
          ) ;
    nor02_2x L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix105 (.Y (
             L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_13), .A0 (nx8014), .A1 (
             nx3924)) ;
    inv01 ix3923 (.Y (nx3924), .A (L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_14)
          ) ;
    nor02_2x L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix109 (.Y (
             L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_14), .A0 (nx8016), .A1 (
             nx3926)) ;
    inv01 ix3925 (.Y (nx3926), .A (L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_15)
          ) ;
    nor02_2x L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix113 (.Y (
             L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_15), .A0 (nx8016), .A1 (
             nx3928)) ;
    inv01 ix3927 (.Y (nx3928), .A (L1_2_L2_0_G1_MINI_ALU_BoothPBeforeShift_16)
          ) ;
    nor02_2x L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix117 (.Y (
             L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_16), .A0 (nx8016), .A1 (
             nx3928)) ;
    mux21 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix189 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BoothOperand_0), .A0 (nx3930), .A1 (nx3932), .S0 (
          nx8004)) ;
    inv01 ix3929 (.Y (nx3930), .A (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_0)) ;
    inv01 ix3931 (.Y (nx3932), .A (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_0)) ;
    mux21 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix197 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BoothOperand_1), .A0 (nx3934), .A1 (nx3936), .S0 (
          nx8004)) ;
    inv01 ix3933 (.Y (nx3934), .A (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_1)) ;
    inv01 ix3935 (.Y (nx3936), .A (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_1)) ;
    mux21 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix205 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BoothOperand_2), .A0 (nx3938), .A1 (nx3940), .S0 (
          nx8004)) ;
    inv01 ix3937 (.Y (nx3938), .A (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_2)) ;
    inv01 ix3939 (.Y (nx3940), .A (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_2)) ;
    mux21 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix213 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BoothOperand_3), .A0 (nx3942), .A1 (nx3944), .S0 (
          nx8004)) ;
    inv01 ix3941 (.Y (nx3942), .A (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_3)) ;
    inv01 ix3943 (.Y (nx3944), .A (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_3)) ;
    mux21 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix221 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BoothOperand_4), .A0 (nx3946), .A1 (nx3948), .S0 (
          nx8004)) ;
    inv01 ix3945 (.Y (nx3946), .A (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_4)) ;
    inv01 ix3947 (.Y (nx3948), .A (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_4)) ;
    mux21 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix229 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BoothOperand_5), .A0 (nx3950), .A1 (nx3952), .S0 (
          nx8006)) ;
    inv01 ix3949 (.Y (nx3950), .A (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_5)) ;
    inv01 ix3951 (.Y (nx3952), .A (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_5)) ;
    mux21 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix237 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BoothOperand_6), .A0 (nx3954), .A1 (nx3956), .S0 (
          nx8006)) ;
    inv01 ix3953 (.Y (nx3954), .A (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_6)) ;
    inv01 ix3955 (.Y (nx3956), .A (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_6)) ;
    mux21 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix245 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BoothOperand_7), .A0 (nx3958), .A1 (nx3960), .S0 (
          nx8006)) ;
    inv01 ix3957 (.Y (nx3958), .A (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_7)) ;
    inv01 ix3959 (.Y (nx3960), .A (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_7)) ;
    mux21 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix253 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BoothOperand_8), .A0 (nx3962), .A1 (nx3964), .S0 (
          nx8006)) ;
    inv01 ix3961 (.Y (nx3962), .A (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_8)) ;
    inv01 ix3963 (.Y (nx3964), .A (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_8)) ;
    mux21 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix261 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BoothOperand_9), .A0 (nx3966), .A1 (nx3968), .S0 (
          nx8006)) ;
    inv01 ix3965 (.Y (nx3966), .A (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_9)) ;
    inv01 ix3967 (.Y (nx3968), .A (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_9)) ;
    mux21 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix269 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BoothOperand_10), .A0 (nx3970), .A1 (nx3972), .S0 (
          nx8006)) ;
    inv01 ix3969 (.Y (nx3970), .A (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_10)) ;
    inv01 ix3971 (.Y (nx3972), .A (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_10)) ;
    mux21 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix277 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BoothOperand_11), .A0 (nx3974), .A1 (nx3976), .S0 (
          nx8006)) ;
    inv01 ix3973 (.Y (nx3974), .A (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_11)) ;
    inv01 ix3975 (.Y (nx3976), .A (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_11)) ;
    mux21 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix285 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BoothOperand_12), .A0 (nx3978), .A1 (nx3980), .S0 (
          nx8008)) ;
    inv01 ix3977 (.Y (nx3978), .A (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_12)) ;
    inv01 ix3979 (.Y (nx3980), .A (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_12)) ;
    mux21 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix293 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BoothOperand_13), .A0 (nx3982), .A1 (nx3984), .S0 (
          nx8008)) ;
    inv01 ix3981 (.Y (nx3982), .A (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_13)) ;
    inv01 ix3983 (.Y (nx3984), .A (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_13)) ;
    mux21 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix301 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BoothOperand_14), .A0 (nx3986), .A1 (nx3988), .S0 (
          nx8008)) ;
    inv01 ix3985 (.Y (nx3986), .A (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_14)) ;
    inv01 ix3987 (.Y (nx3988), .A (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_14)) ;
    mux21 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix309 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BoothOperand_15), .A0 (nx3990), .A1 (nx3992), .S0 (
          nx8008)) ;
    inv01 ix3989 (.Y (nx3990), .A (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_15)) ;
    inv01 ix3991 (.Y (nx3992), .A (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_15)) ;
    mux21 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix317 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BoothOperand_16), .A0 (nx3994), .A1 (nx3996), .S0 (
          nx8008)) ;
    inv01 ix3993 (.Y (nx3994), .A (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_16)) ;
    inv01 ix3995 (.Y (nx3996), .A (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_16)) ;
    xnor2 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_ix321 (.Y (
          L1_2_L2_0_G1_MINI_ALU_AddPToBoothOperand), .A0 (nx8008), .A1 (nx3862)
          ) ;
    oai32 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix393 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .A0 (nx8656), .A1 (
          RST), .A2 (nx8018), .B0 (nx3932), .B1 (nx4000)) ;
    oai32 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix403 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .A0 (nx8656), .A1 (
          RST), .A2 (nx8018), .B0 (nx3936), .B1 (nx4000)) ;
    oai32 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix413 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .A0 (nx8656), .A1 (
          RST), .A2 (nx8018), .B0 (nx3940), .B1 (nx4000)) ;
    oai32 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix423 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .A0 (nx8656), .A1 (
          RST), .A2 (nx8018), .B0 (nx3944), .B1 (nx4000)) ;
    oai32 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix433 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .A0 (nx8656), .A1 (
          RST), .A2 (nx8018), .B0 (nx3948), .B1 (nx4000)) ;
    oai32 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix443 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .A0 (nx8656), .A1 (
          RST), .A2 (nx8018), .B0 (nx3952), .B1 (nx4000)) ;
    oai32 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix453 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .A0 (nx8656), .A1 (
          RST), .A2 (nx8020), .B0 (nx3956), .B1 (nx4000)) ;
    oai32 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix463 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .A0 (nx8658), .A1 (
          RST), .A2 (nx8020), .B0 (nx3960), .B1 (nx4002)) ;
    oai32 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix473 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .A0 (nx8658), .A1 (
          RST), .A2 (nx8020), .B0 (nx3964), .B1 (nx4002)) ;
    oai32 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix483 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .A0 (nx4004), .A1 (
          RST), .A2 (nx8020), .B0 (nx3968), .B1 (nx4002)) ;
    inv01 ix4003 (.Y (nx4004), .A (FilterDin_2__0__0)) ;
    oai32 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix493 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .A0 (nx4006), .A1 (
          RST), .A2 (nx8020), .B0 (nx3972), .B1 (nx4002)) ;
    inv01 ix4005 (.Y (nx4006), .A (FilterDin_2__0__1)) ;
    oai32 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix503 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .A0 (nx4008), .A1 (
          RST), .A2 (nx8020), .B0 (nx3976), .B1 (nx4002)) ;
    inv01 ix4007 (.Y (nx4008), .A (FilterDin_2__0__2)) ;
    oai32 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix513 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .A0 (nx4010), .A1 (
          RST), .A2 (nx8020), .B0 (nx3980), .B1 (nx4002)) ;
    inv01 ix4009 (.Y (nx4010), .A (FilterDin_2__0__3)) ;
    oai32 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix523 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .A0 (nx4012), .A1 (
          RST), .A2 (nx8022), .B0 (nx3984), .B1 (nx4002)) ;
    inv01 ix4011 (.Y (nx4012), .A (FilterDin_2__0__4)) ;
    oai32 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix533 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .A0 (nx4014), .A1 (
          RST), .A2 (nx8022), .B0 (nx3988), .B1 (nx4016)) ;
    inv01 ix4013 (.Y (nx4014), .A (FilterDin_2__0__5)) ;
    inv01 ix4015 (.Y (nx4016), .A (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566)) ;
    oai32 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix543 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .A0 (nx4018), .A1 (
          RST), .A2 (nx8022), .B0 (nx3992), .B1 (nx4016)) ;
    inv01 ix4017 (.Y (nx4018), .A (FilterDin_2__0__6)) ;
    oai32 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix553 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .A0 (nx4020), .A1 (
          RST), .A2 (nx8022), .B0 (nx3996), .B1 (nx4016)) ;
    inv01 ix4019 (.Y (nx4020), .A (FilterDin_2__0__7)) ;
    nand02_2x L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix633 (.Y (nx4000), .A0 (
              nx7592), .A1 (nx8022)) ;
    nand02_2x L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix635 (.Y (nx4002), .A0 (
              nx7592), .A1 (nx8022)) ;
    oai32 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix393 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .A0 (nx8658), .A1 (
          RST), .A2 (nx8024), .B0 (nx3930), .B1 (nx4022)) ;
    oai32 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix403 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .A0 (nx8658), .A1 (
          RST), .A2 (nx8024), .B0 (nx3934), .B1 (nx4022)) ;
    oai32 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix413 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .A0 (nx8658), .A1 (
          RST), .A2 (nx8024), .B0 (nx3938), .B1 (nx4022)) ;
    oai32 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix423 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .A0 (nx8658), .A1 (
          RST), .A2 (nx8024), .B0 (nx3942), .B1 (nx4022)) ;
    oai32 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix433 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .A0 (nx8658), .A1 (
          RST), .A2 (nx8024), .B0 (nx3946), .B1 (nx4022)) ;
    oai32 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix443 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .A0 (nx8660), .A1 (
          RST), .A2 (nx8024), .B0 (nx3950), .B1 (nx4022)) ;
    oai32 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix453 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .A0 (nx8660), .A1 (
          RST), .A2 (nx8026), .B0 (nx3954), .B1 (nx4022)) ;
    oai32 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix463 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .A0 (nx8660), .A1 (
          RST), .A2 (nx8026), .B0 (nx3958), .B1 (nx4024)) ;
    oai32 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix473 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .A0 (nx8660), .A1 (
          RST), .A2 (nx8026), .B0 (nx3962), .B1 (nx4024)) ;
    oai32 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix483 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .A0 (nx4004), .A1 (
          RST), .A2 (nx8026), .B0 (nx3966), .B1 (nx4024)) ;
    oai32 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix493 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .A0 (nx4026), .A1 (
          RST), .A2 (nx8026), .B0 (nx3970), .B1 (nx4024)) ;
    inv01 ix4025 (.Y (nx4026), .A (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_10)) ;
    oai32 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix503 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .A0 (nx4028), .A1 (
          RST), .A2 (nx8026), .B0 (nx3974), .B1 (nx4024)) ;
    inv01 ix4027 (.Y (nx4028), .A (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_11)) ;
    oai32 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix513 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .A0 (nx4030), .A1 (
          RST), .A2 (nx8026), .B0 (nx3978), .B1 (nx4024)) ;
    inv01 ix4029 (.Y (nx4030), .A (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_12)) ;
    oai32 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix523 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .A0 (nx4032), .A1 (
          RST), .A2 (nx8028), .B0 (nx3982), .B1 (nx4024)) ;
    inv01 ix4031 (.Y (nx4032), .A (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_13)) ;
    oai32 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix533 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .A0 (nx4034), .A1 (
          RST), .A2 (nx8028), .B0 (nx3986), .B1 (nx4036)) ;
    inv01 ix4033 (.Y (nx4034), .A (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_14)) ;
    inv01 ix4035 (.Y (nx4036), .A (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566)) ;
    oai32 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix543 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .A0 (nx4038), .A1 (
          RST), .A2 (nx8028), .B0 (nx3990), .B1 (nx4036)) ;
    inv01 ix4037 (.Y (nx4038), .A (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_15)) ;
    oai32 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix553 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .A0 (nx4040), .A1 (
          RST), .A2 (nx8028), .B0 (nx3994), .B1 (nx4036)) ;
    inv01 ix4039 (.Y (nx4040), .A (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_16)) ;
    nand02_2x L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix633 (.Y (nx4022), .A0 (
              nx7592), .A1 (nx8028)) ;
    nand02_2x L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix635 (.Y (nx4024), .A0 (
              nx7594), .A1 (nx8028)) ;
    oai32 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix393 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .A0 (nx4042), .A1 (
          RST), .A2 (nx8030), .B0 (L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx384), .B1 (
          nx4044)) ;
    inv01 ix4041 (.Y (nx4042), .A (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_0)) ;
    oai32 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix403 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .A0 (nx4046), .A1 (
          RST), .A2 (nx8030), .B0 (nx3862), .B1 (nx4044)) ;
    inv01 ix4045 (.Y (nx4046), .A (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_1)) ;
    oai32 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix413 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .A0 (nx4048), .A1 (
          RST), .A2 (nx8030), .B0 (L1_2_L2_0_G1_MINI_ALU_nx387), .B1 (nx4044)) ;
    inv01 ix4047 (.Y (nx4048), .A (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_2)) ;
    oai32 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix423 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .A0 (nx4050), .A1 (
          RST), .A2 (nx8030), .B0 (L1_2_L2_0_G1_MINI_ALU_nx399), .B1 (nx4044)) ;
    inv01 ix4049 (.Y (nx4050), .A (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_3)) ;
    oai32 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix433 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .A0 (nx4052), .A1 (
          RST), .A2 (nx8030), .B0 (L1_2_L2_0_G1_MINI_ALU_nx409), .B1 (nx4044)) ;
    inv01 ix4051 (.Y (nx4052), .A (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_4)) ;
    oai32 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix443 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .A0 (nx4054), .A1 (
          RST), .A2 (nx8030), .B0 (L1_2_L2_0_G1_MINI_ALU_nx419), .B1 (nx4044)) ;
    inv01 ix4053 (.Y (nx4054), .A (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_5)) ;
    oai32 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix453 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .A0 (nx4056), .A1 (
          RST), .A2 (nx8030), .B0 (L1_2_L2_0_G1_MINI_ALU_nx429), .B1 (nx4044)) ;
    inv01 ix4055 (.Y (nx4056), .A (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_6)) ;
    oai32 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix463 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .A0 (nx4058), .A1 (
          RST), .A2 (nx8032), .B0 (L1_2_L2_0_G1_MINI_ALU_nx439), .B1 (nx4060)) ;
    inv01 ix4057 (.Y (nx4058), .A (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_7)) ;
    oai32 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix473 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .A0 (nx4062), .A1 (
          RST), .A2 (nx8032), .B0 (L1_2_L2_0_G1_MINI_ALU_nx449), .B1 (nx4060)) ;
    inv01 ix4061 (.Y (nx4062), .A (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_8)) ;
    oai32 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix483 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .A0 (nx4064), .A1 (
          RST), .A2 (nx8032), .B0 (L1_2_L2_0_G1_MINI_ALU_nx469), .B1 (nx4060)) ;
    inv01 ix4063 (.Y (nx4064), .A (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_9)) ;
    oai32 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix493 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .A0 (nx4066), .A1 (
          RST), .A2 (nx8032), .B0 (L1_2_L2_0_G1_MINI_ALU_nx477), .B1 (nx4060)) ;
    inv01 ix4065 (.Y (nx4066), .A (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_10)) ;
    oai32 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix503 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .A0 (nx4068), .A1 (
          RST), .A2 (nx8032), .B0 (L1_2_L2_0_G1_MINI_ALU_nx485), .B1 (nx4060)) ;
    inv01 ix4067 (.Y (nx4068), .A (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_11)) ;
    oai32 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix513 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .A0 (nx4070), .A1 (
          RST), .A2 (nx8032), .B0 (L1_2_L2_0_G1_MINI_ALU_nx493), .B1 (nx4060)) ;
    inv01 ix4069 (.Y (nx4070), .A (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_12)) ;
    oai32 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix523 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .A0 (nx4072), .A1 (
          RST), .A2 (nx8032), .B0 (L1_2_L2_0_G1_MINI_ALU_nx501), .B1 (nx4060)) ;
    inv01 ix4071 (.Y (nx4072), .A (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_13)) ;
    oai32 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix533 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .A0 (nx4074), .A1 (
          RST), .A2 (nx8034), .B0 (L1_2_L2_0_G1_MINI_ALU_nx509), .B1 (nx4076)) ;
    inv01 ix4073 (.Y (nx4074), .A (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_14)) ;
    inv01 ix4075 (.Y (nx4076), .A (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566)) ;
    oai32 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix543 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .A0 (nx4078), .A1 (
          RST), .A2 (nx8034), .B0 (L1_2_L2_0_G1_MINI_ALU_nx517), .B1 (nx4076)) ;
    inv01 ix4077 (.Y (nx4078), .A (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_15)) ;
    oai32 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix553 (.Y (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .A0 (nx4080), .A1 (
          RST), .A2 (nx8034), .B0 (nx3878), .B1 (nx4076)) ;
    inv01 ix4079 (.Y (nx4080), .A (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_16)) ;
    nand02_2x L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix633 (.Y (nx4044), .A0 (
              nx7594), .A1 (nx8034)) ;
    nand02_2x L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix635 (.Y (nx4060), .A0 (
              nx7594), .A1 (nx8034)) ;
    mux21 L1_2_L2_1_G1_MINI_ALU_ix404 (.Y (L1_2_L2_1_G1_MINI_ALU_nx403), .A0 (
          nx4082), .A1 (L1_2_L2_1_G1_MINI_ALU_BoothP_2), .S0 (
          L1_2_L2_1_G1_MINI_ALU_nx395)) ;
    inv01 ix4081 (.Y (nx4082), .A (L1_2_L2_1_G1_MINI_ALU_nx391)) ;
    mux21 L1_2_L2_1_G1_MINI_ALU_ix414 (.Y (L1_2_L2_1_G1_MINI_ALU_nx413), .A0 (
          nx4084), .A1 (L1_2_L2_1_G1_MINI_ALU_BoothP_3), .S0 (
          L1_2_L2_1_G1_MINI_ALU_nx405)) ;
    inv01 ix4083 (.Y (nx4084), .A (L1_2_L2_1_G1_MINI_ALU_nx403)) ;
    mux21 L1_2_L2_1_G1_MINI_ALU_ix424 (.Y (L1_2_L2_1_G1_MINI_ALU_nx423), .A0 (
          nx4086), .A1 (L1_2_L2_1_G1_MINI_ALU_BoothP_4), .S0 (
          L1_2_L2_1_G1_MINI_ALU_nx415)) ;
    inv01 ix4085 (.Y (nx4086), .A (L1_2_L2_1_G1_MINI_ALU_nx413)) ;
    mux21 L1_2_L2_1_G1_MINI_ALU_ix434 (.Y (L1_2_L2_1_G1_MINI_ALU_nx433), .A0 (
          nx4088), .A1 (L1_2_L2_1_G1_MINI_ALU_BoothP_5), .S0 (
          L1_2_L2_1_G1_MINI_ALU_nx425)) ;
    inv01 ix4087 (.Y (nx4088), .A (L1_2_L2_1_G1_MINI_ALU_nx423)) ;
    mux21 L1_2_L2_1_G1_MINI_ALU_ix444 (.Y (L1_2_L2_1_G1_MINI_ALU_nx443), .A0 (
          nx4090), .A1 (L1_2_L2_1_G1_MINI_ALU_BoothP_6), .S0 (
          L1_2_L2_1_G1_MINI_ALU_nx435)) ;
    inv01 ix4089 (.Y (nx4090), .A (L1_2_L2_1_G1_MINI_ALU_nx433)) ;
    mux21 L1_2_L2_1_G1_MINI_ALU_ix454 (.Y (L1_2_L2_1_G1_MINI_ALU_nx453), .A0 (
          nx4092), .A1 (L1_2_L2_1_G1_MINI_ALU_BoothP_7), .S0 (
          L1_2_L2_1_G1_MINI_ALU_nx445)) ;
    inv01 ix4091 (.Y (nx4092), .A (L1_2_L2_1_G1_MINI_ALU_nx443)) ;
    mux21 L1_2_L2_1_G1_MINI_ALU_ix462 (.Y (L1_2_L2_1_G1_MINI_ALU_nx461), .A0 (
          nx4094), .A1 (L1_2_L2_1_G1_MINI_ALU_BoothP_8), .S0 (
          L1_2_L2_1_G1_MINI_ALU_nx455)) ;
    inv01 ix4093 (.Y (nx4094), .A (L1_2_L2_1_G1_MINI_ALU_nx453)) ;
    mux21 L1_2_L2_1_G1_MINI_ALU_ix468 (.Y (L1_2_L2_1_G1_MINI_ALU_nx467), .A0 (
          nx4096), .A1 (L1_2_L2_1_G1_MINI_ALU_BoothP_9), .S0 (
          L1_2_L2_1_G1_MINI_ALU_nx463)) ;
    inv01 ix4095 (.Y (nx4096), .A (L1_2_L2_1_G1_MINI_ALU_nx461)) ;
    mux21 L1_2_L2_1_G1_MINI_ALU_ix476 (.Y (L1_2_L2_1_G1_MINI_ALU_nx475), .A0 (
          nx4098), .A1 (L1_2_L2_1_G1_MINI_ALU_BoothP_10), .S0 (
          L1_2_L2_1_G1_MINI_ALU_nx471)) ;
    inv01 ix4097 (.Y (nx4098), .A (L1_2_L2_1_G1_MINI_ALU_nx467)) ;
    mux21 L1_2_L2_1_G1_MINI_ALU_ix484 (.Y (L1_2_L2_1_G1_MINI_ALU_nx483), .A0 (
          nx4100), .A1 (L1_2_L2_1_G1_MINI_ALU_BoothP_11), .S0 (
          L1_2_L2_1_G1_MINI_ALU_nx479)) ;
    inv01 ix4099 (.Y (nx4100), .A (L1_2_L2_1_G1_MINI_ALU_nx475)) ;
    mux21 L1_2_L2_1_G1_MINI_ALU_ix492 (.Y (L1_2_L2_1_G1_MINI_ALU_nx491), .A0 (
          nx4102), .A1 (L1_2_L2_1_G1_MINI_ALU_BoothP_12), .S0 (
          L1_2_L2_1_G1_MINI_ALU_nx487)) ;
    inv01 ix4101 (.Y (nx4102), .A (L1_2_L2_1_G1_MINI_ALU_nx483)) ;
    mux21 L1_2_L2_1_G1_MINI_ALU_ix500 (.Y (L1_2_L2_1_G1_MINI_ALU_nx499), .A0 (
          nx4104), .A1 (L1_2_L2_1_G1_MINI_ALU_BoothP_13), .S0 (
          L1_2_L2_1_G1_MINI_ALU_nx495)) ;
    inv01 ix4103 (.Y (nx4104), .A (L1_2_L2_1_G1_MINI_ALU_nx491)) ;
    mux21 L1_2_L2_1_G1_MINI_ALU_ix508 (.Y (L1_2_L2_1_G1_MINI_ALU_nx507), .A0 (
          nx4106), .A1 (L1_2_L2_1_G1_MINI_ALU_BoothP_14), .S0 (
          L1_2_L2_1_G1_MINI_ALU_nx503)) ;
    inv01 ix4105 (.Y (nx4106), .A (L1_2_L2_1_G1_MINI_ALU_nx499)) ;
    mux21 L1_2_L2_1_G1_MINI_ALU_ix516 (.Y (L1_2_L2_1_G1_MINI_ALU_nx515), .A0 (
          nx4108), .A1 (L1_2_L2_1_G1_MINI_ALU_BoothP_15), .S0 (
          L1_2_L2_1_G1_MINI_ALU_nx511)) ;
    inv01 ix4107 (.Y (nx4108), .A (L1_2_L2_1_G1_MINI_ALU_nx507)) ;
    mux21 L1_2_L2_1_G1_MINI_ALU_ix161 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_1), .A0 (nx4110), .A1 (
          L1_2_L2_1_G1_MINI_ALU_nx379), .S0 (nx8038)) ;
    inv01 ix4109 (.Y (nx4110), .A (L1_2_L2_1_G1_MINI_ALU_BoothP_1)) ;
    mux21 L1_2_L2_1_G1_MINI_ALU_ix181 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_2), .A0 (
          L1_2_L2_1_G1_MINI_ALU_nx387), .A1 (L1_2_L2_1_G1_MINI_ALU_nx389), .S0 (
          nx8038)) ;
    mux21 L1_2_L2_1_G1_MINI_ALU_ix201 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_3), .A0 (
          L1_2_L2_1_G1_MINI_ALU_nx399), .A1 (L1_2_L2_1_G1_MINI_ALU_nx401), .S0 (
          nx8038)) ;
    mux21 L1_2_L2_1_G1_MINI_ALU_ix221 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_4), .A0 (
          L1_2_L2_1_G1_MINI_ALU_nx409), .A1 (L1_2_L2_1_G1_MINI_ALU_nx411), .S0 (
          nx8038)) ;
    mux21 L1_2_L2_1_G1_MINI_ALU_ix241 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_5), .A0 (
          L1_2_L2_1_G1_MINI_ALU_nx419), .A1 (L1_2_L2_1_G1_MINI_ALU_nx421), .S0 (
          nx8038)) ;
    mux21 L1_2_L2_1_G1_MINI_ALU_ix261 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_6), .A0 (
          L1_2_L2_1_G1_MINI_ALU_nx429), .A1 (L1_2_L2_1_G1_MINI_ALU_nx431), .S0 (
          nx8038)) ;
    mux21 L1_2_L2_1_G1_MINI_ALU_ix281 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_7), .A0 (
          L1_2_L2_1_G1_MINI_ALU_nx439), .A1 (L1_2_L2_1_G1_MINI_ALU_nx441), .S0 (
          nx8038)) ;
    mux21 L1_2_L2_1_G1_MINI_ALU_ix301 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_8), .A0 (
          L1_2_L2_1_G1_MINI_ALU_nx449), .A1 (L1_2_L2_1_G1_MINI_ALU_nx451), .S0 (
          nx8040)) ;
    mux21 L1_2_L2_1_G1_MINI_ALU_ix321 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_9), .A0 (
          L1_2_L2_1_G1_MINI_ALU_nx469), .A1 (nx4112), .S0 (nx8040)) ;
    inv01 ix4111 (.Y (nx4112), .A (L1_2_L2_1_G1_MINI_ALU_nx316)) ;
    mux21 L1_2_L2_1_G1_MINI_ALU_ix341 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_10), .A0 (
          L1_2_L2_1_G1_MINI_ALU_nx477), .A1 (nx4114), .S0 (nx8040)) ;
    inv01 ix4113 (.Y (nx4114), .A (L1_2_L2_1_G1_MINI_ALU_nx336)) ;
    mux21 L1_2_L2_1_G1_MINI_ALU_ix361 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_11), .A0 (
          L1_2_L2_1_G1_MINI_ALU_nx485), .A1 (nx4116), .S0 (nx8040)) ;
    inv01 ix4115 (.Y (nx4116), .A (L1_2_L2_1_G1_MINI_ALU_nx356)) ;
    mux21 L1_2_L2_1_G1_MINI_ALU_ix381 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_12), .A0 (
          L1_2_L2_1_G1_MINI_ALU_nx493), .A1 (nx4118), .S0 (nx8040)) ;
    inv01 ix4117 (.Y (nx4118), .A (L1_2_L2_1_G1_MINI_ALU_nx376)) ;
    mux21 L1_2_L2_1_G1_MINI_ALU_ix401 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_13), .A0 (
          L1_2_L2_1_G1_MINI_ALU_nx501), .A1 (nx4120), .S0 (nx8040)) ;
    inv01 ix4119 (.Y (nx4120), .A (L1_2_L2_1_G1_MINI_ALU_nx396)) ;
    mux21 L1_2_L2_1_G1_MINI_ALU_ix421 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_14), .A0 (
          L1_2_L2_1_G1_MINI_ALU_nx509), .A1 (nx4122), .S0 (nx8040)) ;
    inv01 ix4121 (.Y (nx4122), .A (L1_2_L2_1_G1_MINI_ALU_nx416)) ;
    mux21 L1_2_L2_1_G1_MINI_ALU_ix441 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_15), .A0 (
          L1_2_L2_1_G1_MINI_ALU_nx517), .A1 (nx4124), .S0 (nx8042)) ;
    inv01 ix4123 (.Y (nx4124), .A (L1_2_L2_1_G1_MINI_ALU_nx436)) ;
    mux21 L1_2_L2_1_G1_MINI_ALU_ix461 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_16), .A0 (nx4126), .A1 (nx4128
          ), .S0 (nx8042)) ;
    inv01 ix4125 (.Y (nx4126), .A (L1_2_L2_1_G1_MINI_ALU_BoothP_16)) ;
    inv01 ix4127 (.Y (nx4128), .A (L1_2_L2_1_G1_MINI_ALU_nx456)) ;
    nor02_2x L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix319 (.Y (
             L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642), .A0 (Start), .A1 (
             CalculatingBooth_dup_1119)) ;
    nor02_2x L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix85 (.Y (
             L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_0), .A0 (nx8052), .A1 (
             nx4130)) ;
    inv01 ix4129 (.Y (nx4130), .A (L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_1)) ;
    mux21 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix125 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_1), .A0 (nx4132), .A1 (
          nx4134), .S0 (nx8052)) ;
    inv01 ix4131 (.Y (nx4132), .A (L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_2)) ;
    inv01 ix4133 (.Y (nx4134), .A (WindowDin_2__1__0)) ;
    mux21 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix133 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_2), .A0 (nx4136), .A1 (
          nx4138), .S0 (nx8052)) ;
    inv01 ix4135 (.Y (nx4136), .A (L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_3)) ;
    inv01 ix4137 (.Y (nx4138), .A (WindowDin_2__1__1)) ;
    mux21 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix141 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_3), .A0 (nx4140), .A1 (
          nx4142), .S0 (nx8052)) ;
    inv01 ix4139 (.Y (nx4140), .A (L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_4)) ;
    inv01 ix4141 (.Y (nx4142), .A (WindowDin_2__1__2)) ;
    mux21 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix149 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_4), .A0 (nx4144), .A1 (
          nx4146), .S0 (nx8052)) ;
    inv01 ix4143 (.Y (nx4144), .A (L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_5)) ;
    inv01 ix4145 (.Y (nx4146), .A (WindowDin_2__1__3)) ;
    mux21 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix157 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_5), .A0 (nx4148), .A1 (
          nx4150), .S0 (nx8052)) ;
    inv01 ix4147 (.Y (nx4148), .A (L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_6)) ;
    inv01 ix4149 (.Y (nx4150), .A (WindowDin_2__1__4)) ;
    mux21 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix165 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_6), .A0 (nx4152), .A1 (
          nx4154), .S0 (nx8052)) ;
    inv01 ix4151 (.Y (nx4152), .A (L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_7)) ;
    inv01 ix4153 (.Y (nx4154), .A (WindowDin_2__1__5)) ;
    mux21 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix173 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_7), .A0 (nx4156), .A1 (
          nx4158), .S0 (nx8054)) ;
    inv01 ix4155 (.Y (nx4156), .A (L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_8)) ;
    inv01 ix4157 (.Y (nx4158), .A (WindowDin_2__1__6)) ;
    mux21 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix181 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_8), .A0 (nx4160), .A1 (
          nx4162), .S0 (nx8054)) ;
    inv01 ix4159 (.Y (nx4160), .A (L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_9)) ;
    inv01 ix4161 (.Y (nx4162), .A (WindowDin_2__1__7)) ;
    nor02_2x L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix89 (.Y (
             L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_9), .A0 (nx8054), .A1 (
             nx4164)) ;
    inv01 ix4163 (.Y (nx4164), .A (L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_10)
          ) ;
    nor02_2x L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix93 (.Y (
             L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_10), .A0 (nx8054), .A1 (
             nx4166)) ;
    inv01 ix4165 (.Y (nx4166), .A (L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_11)
          ) ;
    nor02_2x L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix97 (.Y (
             L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_11), .A0 (nx8054), .A1 (
             nx4168)) ;
    inv01 ix4167 (.Y (nx4168), .A (L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_12)
          ) ;
    nor02_2x L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix101 (.Y (
             L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_12), .A0 (nx8054), .A1 (
             nx4170)) ;
    inv01 ix4169 (.Y (nx4170), .A (L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_13)
          ) ;
    nor02_2x L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix105 (.Y (
             L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_13), .A0 (nx8054), .A1 (
             nx4172)) ;
    inv01 ix4171 (.Y (nx4172), .A (L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_14)
          ) ;
    nor02_2x L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix109 (.Y (
             L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_14), .A0 (nx8056), .A1 (
             nx4174)) ;
    inv01 ix4173 (.Y (nx4174), .A (L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_15)
          ) ;
    nor02_2x L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix113 (.Y (
             L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_15), .A0 (nx8056), .A1 (
             nx4176)) ;
    inv01 ix4175 (.Y (nx4176), .A (L1_2_L2_1_G1_MINI_ALU_BoothPBeforeShift_16)
          ) ;
    nor02_2x L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix117 (.Y (
             L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_16), .A0 (nx8056), .A1 (
             nx4176)) ;
    mux21 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix189 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BoothOperand_0), .A0 (nx4178), .A1 (nx4180), .S0 (
          nx8044)) ;
    inv01 ix4177 (.Y (nx4178), .A (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_0)) ;
    inv01 ix4179 (.Y (nx4180), .A (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_0)) ;
    mux21 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix197 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BoothOperand_1), .A0 (nx4182), .A1 (nx4184), .S0 (
          nx8044)) ;
    inv01 ix4181 (.Y (nx4182), .A (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_1)) ;
    inv01 ix4183 (.Y (nx4184), .A (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_1)) ;
    mux21 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix205 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BoothOperand_2), .A0 (nx4186), .A1 (nx4188), .S0 (
          nx8044)) ;
    inv01 ix4185 (.Y (nx4186), .A (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_2)) ;
    inv01 ix4187 (.Y (nx4188), .A (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_2)) ;
    mux21 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix213 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BoothOperand_3), .A0 (nx4190), .A1 (nx4192), .S0 (
          nx8044)) ;
    inv01 ix4189 (.Y (nx4190), .A (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_3)) ;
    inv01 ix4191 (.Y (nx4192), .A (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_3)) ;
    mux21 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix221 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BoothOperand_4), .A0 (nx4194), .A1 (nx4196), .S0 (
          nx8044)) ;
    inv01 ix4193 (.Y (nx4194), .A (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_4)) ;
    inv01 ix4195 (.Y (nx4196), .A (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_4)) ;
    mux21 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix229 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BoothOperand_5), .A0 (nx4198), .A1 (nx4200), .S0 (
          nx8046)) ;
    inv01 ix4197 (.Y (nx4198), .A (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_5)) ;
    inv01 ix4199 (.Y (nx4200), .A (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_5)) ;
    mux21 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix237 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BoothOperand_6), .A0 (nx4202), .A1 (nx4204), .S0 (
          nx8046)) ;
    inv01 ix4201 (.Y (nx4202), .A (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_6)) ;
    inv01 ix4203 (.Y (nx4204), .A (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_6)) ;
    mux21 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix245 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BoothOperand_7), .A0 (nx4206), .A1 (nx4208), .S0 (
          nx8046)) ;
    inv01 ix4205 (.Y (nx4206), .A (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_7)) ;
    inv01 ix4207 (.Y (nx4208), .A (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_7)) ;
    mux21 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix253 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BoothOperand_8), .A0 (nx4210), .A1 (nx4212), .S0 (
          nx8046)) ;
    inv01 ix4209 (.Y (nx4210), .A (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_8)) ;
    inv01 ix4211 (.Y (nx4212), .A (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_8)) ;
    mux21 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix261 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BoothOperand_9), .A0 (nx4214), .A1 (nx4216), .S0 (
          nx8046)) ;
    inv01 ix4213 (.Y (nx4214), .A (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_9)) ;
    inv01 ix4215 (.Y (nx4216), .A (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_9)) ;
    mux21 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix269 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BoothOperand_10), .A0 (nx4218), .A1 (nx4220), .S0 (
          nx8046)) ;
    inv01 ix4217 (.Y (nx4218), .A (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_10)) ;
    inv01 ix4219 (.Y (nx4220), .A (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_10)) ;
    mux21 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix277 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BoothOperand_11), .A0 (nx4222), .A1 (nx4224), .S0 (
          nx8046)) ;
    inv01 ix4221 (.Y (nx4222), .A (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_11)) ;
    inv01 ix4223 (.Y (nx4224), .A (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_11)) ;
    mux21 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix285 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BoothOperand_12), .A0 (nx4226), .A1 (nx4228), .S0 (
          nx8048)) ;
    inv01 ix4225 (.Y (nx4226), .A (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_12)) ;
    inv01 ix4227 (.Y (nx4228), .A (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_12)) ;
    mux21 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix293 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BoothOperand_13), .A0 (nx4230), .A1 (nx4232), .S0 (
          nx8048)) ;
    inv01 ix4229 (.Y (nx4230), .A (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_13)) ;
    inv01 ix4231 (.Y (nx4232), .A (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_13)) ;
    mux21 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix301 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BoothOperand_14), .A0 (nx4234), .A1 (nx4236), .S0 (
          nx8048)) ;
    inv01 ix4233 (.Y (nx4234), .A (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_14)) ;
    inv01 ix4235 (.Y (nx4236), .A (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_14)) ;
    mux21 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix309 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BoothOperand_15), .A0 (nx4238), .A1 (nx4240), .S0 (
          nx8048)) ;
    inv01 ix4237 (.Y (nx4238), .A (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_15)) ;
    inv01 ix4239 (.Y (nx4240), .A (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_15)) ;
    mux21 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix317 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BoothOperand_16), .A0 (nx4242), .A1 (nx4244), .S0 (
          nx8048)) ;
    inv01 ix4241 (.Y (nx4242), .A (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_16)) ;
    inv01 ix4243 (.Y (nx4244), .A (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_16)) ;
    xnor2 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_ix321 (.Y (
          L1_2_L2_1_G1_MINI_ALU_AddPToBoothOperand), .A0 (nx8048), .A1 (nx4110)
          ) ;
    oai32 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix393 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .A0 (nx8662), .A1 (
          RST), .A2 (nx8058), .B0 (nx4180), .B1 (nx4248)) ;
    oai32 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix403 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .A0 (nx8662), .A1 (
          RST), .A2 (nx8058), .B0 (nx4184), .B1 (nx4248)) ;
    oai32 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix413 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .A0 (nx8662), .A1 (
          RST), .A2 (nx8058), .B0 (nx4188), .B1 (nx4248)) ;
    oai32 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix423 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .A0 (nx8662), .A1 (
          RST), .A2 (nx8058), .B0 (nx4192), .B1 (nx4248)) ;
    oai32 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix433 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .A0 (nx8662), .A1 (
          RST), .A2 (nx8058), .B0 (nx4196), .B1 (nx4248)) ;
    oai32 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix443 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .A0 (nx8662), .A1 (
          RST), .A2 (nx8058), .B0 (nx4200), .B1 (nx4248)) ;
    oai32 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix453 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .A0 (nx8662), .A1 (
          RST), .A2 (nx8060), .B0 (nx4204), .B1 (nx4248)) ;
    oai32 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix463 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .A0 (nx8664), .A1 (
          RST), .A2 (nx8060), .B0 (nx4208), .B1 (nx4250)) ;
    oai32 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix473 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .A0 (nx8664), .A1 (
          RST), .A2 (nx8060), .B0 (nx4212), .B1 (nx4250)) ;
    oai32 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix483 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .A0 (nx4252), .A1 (
          RST), .A2 (nx8060), .B0 (nx4216), .B1 (nx4250)) ;
    inv01 ix4251 (.Y (nx4252), .A (FilterDin_2__1__0)) ;
    oai32 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix493 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .A0 (nx4254), .A1 (
          RST), .A2 (nx8060), .B0 (nx4220), .B1 (nx4250)) ;
    inv01 ix4253 (.Y (nx4254), .A (FilterDin_2__1__1)) ;
    oai32 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix503 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .A0 (nx4256), .A1 (
          RST), .A2 (nx8060), .B0 (nx4224), .B1 (nx4250)) ;
    inv01 ix4255 (.Y (nx4256), .A (FilterDin_2__1__2)) ;
    oai32 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix513 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .A0 (nx4258), .A1 (
          RST), .A2 (nx8060), .B0 (nx4228), .B1 (nx4250)) ;
    inv01 ix4257 (.Y (nx4258), .A (FilterDin_2__1__3)) ;
    oai32 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix523 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .A0 (nx4260), .A1 (
          RST), .A2 (nx8062), .B0 (nx4232), .B1 (nx4250)) ;
    inv01 ix4259 (.Y (nx4260), .A (FilterDin_2__1__4)) ;
    oai32 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix533 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .A0 (nx4262), .A1 (
          RST), .A2 (nx8062), .B0 (nx4236), .B1 (nx4264)) ;
    inv01 ix4261 (.Y (nx4262), .A (FilterDin_2__1__5)) ;
    inv01 ix4263 (.Y (nx4264), .A (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566)) ;
    oai32 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix543 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .A0 (nx4266), .A1 (
          RST), .A2 (nx8062), .B0 (nx4240), .B1 (nx4264)) ;
    inv01 ix4265 (.Y (nx4266), .A (FilterDin_2__1__6)) ;
    oai32 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix553 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .A0 (nx4268), .A1 (
          RST), .A2 (nx8062), .B0 (nx4244), .B1 (nx4264)) ;
    inv01 ix4267 (.Y (nx4268), .A (FilterDin_2__1__7)) ;
    nand02_2x L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix633 (.Y (nx4248), .A0 (
              nx7594), .A1 (nx8062)) ;
    nand02_2x L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix635 (.Y (nx4250), .A0 (
              nx7594), .A1 (nx8062)) ;
    oai32 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix393 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .A0 (nx8664), .A1 (
          RST), .A2 (nx8064), .B0 (nx4178), .B1 (nx4270)) ;
    oai32 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix403 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .A0 (nx8664), .A1 (
          RST), .A2 (nx8064), .B0 (nx4182), .B1 (nx4270)) ;
    oai32 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix413 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .A0 (nx8664), .A1 (
          RST), .A2 (nx8064), .B0 (nx4186), .B1 (nx4270)) ;
    oai32 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix423 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .A0 (nx8664), .A1 (
          RST), .A2 (nx8064), .B0 (nx4190), .B1 (nx4270)) ;
    oai32 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix433 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .A0 (nx8664), .A1 (
          RST), .A2 (nx8064), .B0 (nx4194), .B1 (nx4270)) ;
    oai32 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix443 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .A0 (nx8666), .A1 (
          RST), .A2 (nx8064), .B0 (nx4198), .B1 (nx4270)) ;
    oai32 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix453 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .A0 (nx8666), .A1 (
          RST), .A2 (nx8066), .B0 (nx4202), .B1 (nx4270)) ;
    oai32 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix463 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .A0 (nx8666), .A1 (
          RST), .A2 (nx8066), .B0 (nx4206), .B1 (nx4272)) ;
    oai32 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix473 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .A0 (nx8666), .A1 (
          RST), .A2 (nx8066), .B0 (nx4210), .B1 (nx4272)) ;
    oai32 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix483 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .A0 (nx4252), .A1 (
          RST), .A2 (nx8066), .B0 (nx4214), .B1 (nx4272)) ;
    oai32 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix493 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .A0 (nx4274), .A1 (
          RST), .A2 (nx8066), .B0 (nx4218), .B1 (nx4272)) ;
    inv01 ix4273 (.Y (nx4274), .A (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_10)) ;
    oai32 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix503 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .A0 (nx4276), .A1 (
          RST), .A2 (nx8066), .B0 (nx4222), .B1 (nx4272)) ;
    inv01 ix4275 (.Y (nx4276), .A (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_11)) ;
    oai32 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix513 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .A0 (nx4278), .A1 (
          RST), .A2 (nx8066), .B0 (nx4226), .B1 (nx4272)) ;
    inv01 ix4277 (.Y (nx4278), .A (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_12)) ;
    oai32 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix523 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .A0 (nx4280), .A1 (
          RST), .A2 (nx8068), .B0 (nx4230), .B1 (nx4272)) ;
    inv01 ix4279 (.Y (nx4280), .A (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_13)) ;
    oai32 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix533 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .A0 (nx4282), .A1 (
          RST), .A2 (nx8068), .B0 (nx4234), .B1 (nx4284)) ;
    inv01 ix4281 (.Y (nx4282), .A (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_14)) ;
    inv01 ix4283 (.Y (nx4284), .A (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566)) ;
    oai32 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix543 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .A0 (nx4286), .A1 (
          RST), .A2 (nx8068), .B0 (nx4238), .B1 (nx4284)) ;
    inv01 ix4285 (.Y (nx4286), .A (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_15)) ;
    oai32 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix553 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .A0 (nx4288), .A1 (
          RST), .A2 (nx8068), .B0 (nx4242), .B1 (nx4284)) ;
    inv01 ix4287 (.Y (nx4288), .A (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_16)) ;
    nand02_2x L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix633 (.Y (nx4270), .A0 (
              nx7594), .A1 (nx8068)) ;
    nand02_2x L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix635 (.Y (nx4272), .A0 (
              nx7594), .A1 (nx8068)) ;
    oai32 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix393 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .A0 (nx4290), .A1 (
          RST), .A2 (nx8070), .B0 (L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx384), .B1 (
          nx4292)) ;
    inv01 ix4289 (.Y (nx4290), .A (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_0)) ;
    oai32 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix403 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .A0 (nx4294), .A1 (
          RST), .A2 (nx8070), .B0 (nx4110), .B1 (nx4292)) ;
    inv01 ix4293 (.Y (nx4294), .A (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_1)) ;
    oai32 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix413 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .A0 (nx4296), .A1 (
          RST), .A2 (nx8070), .B0 (L1_2_L2_1_G1_MINI_ALU_nx387), .B1 (nx4292)) ;
    inv01 ix4295 (.Y (nx4296), .A (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_2)) ;
    oai32 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix423 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .A0 (nx4298), .A1 (
          RST), .A2 (nx8070), .B0 (L1_2_L2_1_G1_MINI_ALU_nx399), .B1 (nx4292)) ;
    inv01 ix4297 (.Y (nx4298), .A (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_3)) ;
    oai32 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix433 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .A0 (nx4300), .A1 (
          RST), .A2 (nx8070), .B0 (L1_2_L2_1_G1_MINI_ALU_nx409), .B1 (nx4292)) ;
    inv01 ix4299 (.Y (nx4300), .A (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_4)) ;
    oai32 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix443 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .A0 (nx4302), .A1 (
          RST), .A2 (nx8070), .B0 (L1_2_L2_1_G1_MINI_ALU_nx419), .B1 (nx4292)) ;
    inv01 ix4301 (.Y (nx4302), .A (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_5)) ;
    oai32 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix453 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .A0 (nx4304), .A1 (
          RST), .A2 (nx8070), .B0 (L1_2_L2_1_G1_MINI_ALU_nx429), .B1 (nx4292)) ;
    inv01 ix4303 (.Y (nx4304), .A (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_6)) ;
    oai32 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix463 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .A0 (nx4306), .A1 (
          RST), .A2 (nx8072), .B0 (L1_2_L2_1_G1_MINI_ALU_nx439), .B1 (nx4308)) ;
    inv01 ix4305 (.Y (nx4306), .A (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_7)) ;
    oai32 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix473 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .A0 (nx4310), .A1 (
          RST), .A2 (nx8072), .B0 (L1_2_L2_1_G1_MINI_ALU_nx449), .B1 (nx4308)) ;
    inv01 ix4309 (.Y (nx4310), .A (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_8)) ;
    oai32 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix483 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .A0 (nx4312), .A1 (
          RST), .A2 (nx8072), .B0 (L1_2_L2_1_G1_MINI_ALU_nx469), .B1 (nx4308)) ;
    inv01 ix4311 (.Y (nx4312), .A (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_9)) ;
    oai32 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix493 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .A0 (nx4314), .A1 (
          RST), .A2 (nx8072), .B0 (L1_2_L2_1_G1_MINI_ALU_nx477), .B1 (nx4308)) ;
    inv01 ix4313 (.Y (nx4314), .A (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_10)) ;
    oai32 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix503 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .A0 (nx4316), .A1 (
          RST), .A2 (nx8072), .B0 (L1_2_L2_1_G1_MINI_ALU_nx485), .B1 (nx4308)) ;
    inv01 ix4315 (.Y (nx4316), .A (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_11)) ;
    oai32 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix513 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .A0 (nx4318), .A1 (
          RST), .A2 (nx8072), .B0 (L1_2_L2_1_G1_MINI_ALU_nx493), .B1 (nx4308)) ;
    inv01 ix4317 (.Y (nx4318), .A (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_12)) ;
    oai32 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix523 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .A0 (nx4320), .A1 (
          RST), .A2 (nx8072), .B0 (L1_2_L2_1_G1_MINI_ALU_nx501), .B1 (nx4308)) ;
    inv01 ix4319 (.Y (nx4320), .A (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_13)) ;
    oai32 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix533 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .A0 (nx4322), .A1 (
          RST), .A2 (nx8074), .B0 (L1_2_L2_1_G1_MINI_ALU_nx509), .B1 (nx4324)) ;
    inv01 ix4321 (.Y (nx4322), .A (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_14)) ;
    inv01 ix4323 (.Y (nx4324), .A (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566)) ;
    oai32 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix543 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .A0 (nx4326), .A1 (
          RST), .A2 (nx8074), .B0 (L1_2_L2_1_G1_MINI_ALU_nx517), .B1 (nx4324)) ;
    inv01 ix4325 (.Y (nx4326), .A (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_15)) ;
    oai32 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix553 (.Y (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .A0 (nx4328), .A1 (
          RST), .A2 (nx8074), .B0 (nx4126), .B1 (nx4324)) ;
    inv01 ix4327 (.Y (nx4328), .A (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_16)) ;
    nand02_2x L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix633 (.Y (nx4292), .A0 (
              nx7596), .A1 (nx8074)) ;
    nand02_2x L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix635 (.Y (nx4308), .A0 (
              nx7596), .A1 (nx8074)) ;
    mux21 L1_2_L2_2_G1_MINI_ALU_ix404 (.Y (L1_2_L2_2_G1_MINI_ALU_nx403), .A0 (
          nx4330), .A1 (L1_2_L2_2_G1_MINI_ALU_BoothP_2), .S0 (
          L1_2_L2_2_G1_MINI_ALU_nx395)) ;
    inv01 ix4329 (.Y (nx4330), .A (L1_2_L2_2_G1_MINI_ALU_nx391)) ;
    mux21 L1_2_L2_2_G1_MINI_ALU_ix414 (.Y (L1_2_L2_2_G1_MINI_ALU_nx413), .A0 (
          nx4332), .A1 (L1_2_L2_2_G1_MINI_ALU_BoothP_3), .S0 (
          L1_2_L2_2_G1_MINI_ALU_nx405)) ;
    inv01 ix4331 (.Y (nx4332), .A (L1_2_L2_2_G1_MINI_ALU_nx403)) ;
    mux21 L1_2_L2_2_G1_MINI_ALU_ix424 (.Y (L1_2_L2_2_G1_MINI_ALU_nx423), .A0 (
          nx4334), .A1 (L1_2_L2_2_G1_MINI_ALU_BoothP_4), .S0 (
          L1_2_L2_2_G1_MINI_ALU_nx415)) ;
    inv01 ix4333 (.Y (nx4334), .A (L1_2_L2_2_G1_MINI_ALU_nx413)) ;
    mux21 L1_2_L2_2_G1_MINI_ALU_ix434 (.Y (L1_2_L2_2_G1_MINI_ALU_nx433), .A0 (
          nx4336), .A1 (L1_2_L2_2_G1_MINI_ALU_BoothP_5), .S0 (
          L1_2_L2_2_G1_MINI_ALU_nx425)) ;
    inv01 ix4335 (.Y (nx4336), .A (L1_2_L2_2_G1_MINI_ALU_nx423)) ;
    mux21 L1_2_L2_2_G1_MINI_ALU_ix444 (.Y (L1_2_L2_2_G1_MINI_ALU_nx443), .A0 (
          nx4338), .A1 (L1_2_L2_2_G1_MINI_ALU_BoothP_6), .S0 (
          L1_2_L2_2_G1_MINI_ALU_nx435)) ;
    inv01 ix4337 (.Y (nx4338), .A (L1_2_L2_2_G1_MINI_ALU_nx433)) ;
    mux21 L1_2_L2_2_G1_MINI_ALU_ix454 (.Y (L1_2_L2_2_G1_MINI_ALU_nx453), .A0 (
          nx4340), .A1 (L1_2_L2_2_G1_MINI_ALU_BoothP_7), .S0 (
          L1_2_L2_2_G1_MINI_ALU_nx445)) ;
    inv01 ix4339 (.Y (nx4340), .A (L1_2_L2_2_G1_MINI_ALU_nx443)) ;
    mux21 L1_2_L2_2_G1_MINI_ALU_ix462 (.Y (L1_2_L2_2_G1_MINI_ALU_nx461), .A0 (
          nx4342), .A1 (L1_2_L2_2_G1_MINI_ALU_BoothP_8), .S0 (
          L1_2_L2_2_G1_MINI_ALU_nx455)) ;
    inv01 ix4341 (.Y (nx4342), .A (L1_2_L2_2_G1_MINI_ALU_nx453)) ;
    mux21 L1_2_L2_2_G1_MINI_ALU_ix468 (.Y (L1_2_L2_2_G1_MINI_ALU_nx467), .A0 (
          nx4344), .A1 (L1_2_L2_2_G1_MINI_ALU_BoothP_9), .S0 (
          L1_2_L2_2_G1_MINI_ALU_nx463)) ;
    inv01 ix4343 (.Y (nx4344), .A (L1_2_L2_2_G1_MINI_ALU_nx461)) ;
    mux21 L1_2_L2_2_G1_MINI_ALU_ix476 (.Y (L1_2_L2_2_G1_MINI_ALU_nx475), .A0 (
          nx4346), .A1 (L1_2_L2_2_G1_MINI_ALU_BoothP_10), .S0 (
          L1_2_L2_2_G1_MINI_ALU_nx471)) ;
    inv01 ix4345 (.Y (nx4346), .A (L1_2_L2_2_G1_MINI_ALU_nx467)) ;
    mux21 L1_2_L2_2_G1_MINI_ALU_ix484 (.Y (L1_2_L2_2_G1_MINI_ALU_nx483), .A0 (
          nx4348), .A1 (L1_2_L2_2_G1_MINI_ALU_BoothP_11), .S0 (
          L1_2_L2_2_G1_MINI_ALU_nx479)) ;
    inv01 ix4347 (.Y (nx4348), .A (L1_2_L2_2_G1_MINI_ALU_nx475)) ;
    mux21 L1_2_L2_2_G1_MINI_ALU_ix492 (.Y (L1_2_L2_2_G1_MINI_ALU_nx491), .A0 (
          nx4350), .A1 (L1_2_L2_2_G1_MINI_ALU_BoothP_12), .S0 (
          L1_2_L2_2_G1_MINI_ALU_nx487)) ;
    inv01 ix4349 (.Y (nx4350), .A (L1_2_L2_2_G1_MINI_ALU_nx483)) ;
    mux21 L1_2_L2_2_G1_MINI_ALU_ix500 (.Y (L1_2_L2_2_G1_MINI_ALU_nx499), .A0 (
          nx4352), .A1 (L1_2_L2_2_G1_MINI_ALU_BoothP_13), .S0 (
          L1_2_L2_2_G1_MINI_ALU_nx495)) ;
    inv01 ix4351 (.Y (nx4352), .A (L1_2_L2_2_G1_MINI_ALU_nx491)) ;
    mux21 L1_2_L2_2_G1_MINI_ALU_ix508 (.Y (L1_2_L2_2_G1_MINI_ALU_nx507), .A0 (
          nx4354), .A1 (L1_2_L2_2_G1_MINI_ALU_BoothP_14), .S0 (
          L1_2_L2_2_G1_MINI_ALU_nx503)) ;
    inv01 ix4353 (.Y (nx4354), .A (L1_2_L2_2_G1_MINI_ALU_nx499)) ;
    mux21 L1_2_L2_2_G1_MINI_ALU_ix516 (.Y (L1_2_L2_2_G1_MINI_ALU_nx515), .A0 (
          nx4356), .A1 (L1_2_L2_2_G1_MINI_ALU_BoothP_15), .S0 (
          L1_2_L2_2_G1_MINI_ALU_nx511)) ;
    inv01 ix4355 (.Y (nx4356), .A (L1_2_L2_2_G1_MINI_ALU_nx507)) ;
    mux21 L1_2_L2_2_G1_MINI_ALU_ix161 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_1), .A0 (nx4358), .A1 (
          L1_2_L2_2_G1_MINI_ALU_nx379), .S0 (nx8078)) ;
    inv01 ix4357 (.Y (nx4358), .A (L1_2_L2_2_G1_MINI_ALU_BoothP_1)) ;
    mux21 L1_2_L2_2_G1_MINI_ALU_ix181 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_2), .A0 (
          L1_2_L2_2_G1_MINI_ALU_nx387), .A1 (L1_2_L2_2_G1_MINI_ALU_nx389), .S0 (
          nx8078)) ;
    mux21 L1_2_L2_2_G1_MINI_ALU_ix201 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_3), .A0 (
          L1_2_L2_2_G1_MINI_ALU_nx399), .A1 (L1_2_L2_2_G1_MINI_ALU_nx401), .S0 (
          nx8078)) ;
    mux21 L1_2_L2_2_G1_MINI_ALU_ix221 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_4), .A0 (
          L1_2_L2_2_G1_MINI_ALU_nx409), .A1 (L1_2_L2_2_G1_MINI_ALU_nx411), .S0 (
          nx8078)) ;
    mux21 L1_2_L2_2_G1_MINI_ALU_ix241 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_5), .A0 (
          L1_2_L2_2_G1_MINI_ALU_nx419), .A1 (L1_2_L2_2_G1_MINI_ALU_nx421), .S0 (
          nx8078)) ;
    mux21 L1_2_L2_2_G1_MINI_ALU_ix261 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_6), .A0 (
          L1_2_L2_2_G1_MINI_ALU_nx429), .A1 (L1_2_L2_2_G1_MINI_ALU_nx431), .S0 (
          nx8078)) ;
    mux21 L1_2_L2_2_G1_MINI_ALU_ix281 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_7), .A0 (
          L1_2_L2_2_G1_MINI_ALU_nx439), .A1 (L1_2_L2_2_G1_MINI_ALU_nx441), .S0 (
          nx8078)) ;
    mux21 L1_2_L2_2_G1_MINI_ALU_ix301 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_8), .A0 (
          L1_2_L2_2_G1_MINI_ALU_nx449), .A1 (L1_2_L2_2_G1_MINI_ALU_nx451), .S0 (
          nx8080)) ;
    mux21 L1_2_L2_2_G1_MINI_ALU_ix321 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_9), .A0 (
          L1_2_L2_2_G1_MINI_ALU_nx469), .A1 (nx4360), .S0 (nx8080)) ;
    inv01 ix4359 (.Y (nx4360), .A (L1_2_L2_2_G1_MINI_ALU_nx316)) ;
    mux21 L1_2_L2_2_G1_MINI_ALU_ix341 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_10), .A0 (
          L1_2_L2_2_G1_MINI_ALU_nx477), .A1 (nx4362), .S0 (nx8080)) ;
    inv01 ix4361 (.Y (nx4362), .A (L1_2_L2_2_G1_MINI_ALU_nx336)) ;
    mux21 L1_2_L2_2_G1_MINI_ALU_ix361 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_11), .A0 (
          L1_2_L2_2_G1_MINI_ALU_nx485), .A1 (nx4364), .S0 (nx8080)) ;
    inv01 ix4363 (.Y (nx4364), .A (L1_2_L2_2_G1_MINI_ALU_nx356)) ;
    mux21 L1_2_L2_2_G1_MINI_ALU_ix381 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_12), .A0 (
          L1_2_L2_2_G1_MINI_ALU_nx493), .A1 (nx4366), .S0 (nx8080)) ;
    inv01 ix4365 (.Y (nx4366), .A (L1_2_L2_2_G1_MINI_ALU_nx376)) ;
    mux21 L1_2_L2_2_G1_MINI_ALU_ix401 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_13), .A0 (
          L1_2_L2_2_G1_MINI_ALU_nx501), .A1 (nx4368), .S0 (nx8080)) ;
    inv01 ix4367 (.Y (nx4368), .A (L1_2_L2_2_G1_MINI_ALU_nx396)) ;
    mux21 L1_2_L2_2_G1_MINI_ALU_ix421 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_14), .A0 (
          L1_2_L2_2_G1_MINI_ALU_nx509), .A1 (nx4370), .S0 (nx8080)) ;
    inv01 ix4369 (.Y (nx4370), .A (L1_2_L2_2_G1_MINI_ALU_nx416)) ;
    mux21 L1_2_L2_2_G1_MINI_ALU_ix441 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_15), .A0 (
          L1_2_L2_2_G1_MINI_ALU_nx517), .A1 (nx4372), .S0 (nx8082)) ;
    inv01 ix4371 (.Y (nx4372), .A (L1_2_L2_2_G1_MINI_ALU_nx436)) ;
    mux21 L1_2_L2_2_G1_MINI_ALU_ix461 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_16), .A0 (nx4374), .A1 (nx4376
          ), .S0 (nx8082)) ;
    inv01 ix4373 (.Y (nx4374), .A (L1_2_L2_2_G1_MINI_ALU_BoothP_16)) ;
    inv01 ix4375 (.Y (nx4376), .A (L1_2_L2_2_G1_MINI_ALU_nx456)) ;
    nor02_2x L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix319 (.Y (
             L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642), .A0 (Start), .A1 (
             CalculatingBooth_dup_1119)) ;
    nor02_2x L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix85 (.Y (
             L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_0), .A0 (nx8092), .A1 (
             nx4378)) ;
    inv01 ix4377 (.Y (nx4378), .A (L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_1)) ;
    mux21 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix125 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_1), .A0 (nx4380), .A1 (
          nx4382), .S0 (nx8092)) ;
    inv01 ix4379 (.Y (nx4380), .A (L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_2)) ;
    inv01 ix4381 (.Y (nx4382), .A (WindowDin_2__2__0)) ;
    mux21 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix133 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_2), .A0 (nx4384), .A1 (
          nx4386), .S0 (nx8092)) ;
    inv01 ix4383 (.Y (nx4384), .A (L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_3)) ;
    inv01 ix4385 (.Y (nx4386), .A (WindowDin_2__2__1)) ;
    mux21 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix141 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_3), .A0 (nx4388), .A1 (
          nx4390), .S0 (nx8092)) ;
    inv01 ix4387 (.Y (nx4388), .A (L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_4)) ;
    inv01 ix4389 (.Y (nx4390), .A (WindowDin_2__2__2)) ;
    mux21 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix149 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_4), .A0 (nx4392), .A1 (
          nx4394), .S0 (nx8092)) ;
    inv01 ix4391 (.Y (nx4392), .A (L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_5)) ;
    inv01 ix4393 (.Y (nx4394), .A (WindowDin_2__2__3)) ;
    mux21 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix157 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_5), .A0 (nx4396), .A1 (
          nx4398), .S0 (nx8092)) ;
    inv01 ix4395 (.Y (nx4396), .A (L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_6)) ;
    inv01 ix4397 (.Y (nx4398), .A (WindowDin_2__2__4)) ;
    mux21 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix165 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_6), .A0 (nx4400), .A1 (
          nx4402), .S0 (nx8092)) ;
    inv01 ix4399 (.Y (nx4400), .A (L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_7)) ;
    inv01 ix4401 (.Y (nx4402), .A (WindowDin_2__2__5)) ;
    mux21 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix173 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_7), .A0 (nx4404), .A1 (
          nx4406), .S0 (nx8094)) ;
    inv01 ix4403 (.Y (nx4404), .A (L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_8)) ;
    inv01 ix4405 (.Y (nx4406), .A (WindowDin_2__2__6)) ;
    mux21 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix181 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_8), .A0 (nx4408), .A1 (
          nx4410), .S0 (nx8094)) ;
    inv01 ix4407 (.Y (nx4408), .A (L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_9)) ;
    inv01 ix4409 (.Y (nx4410), .A (WindowDin_2__2__7)) ;
    nor02_2x L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix89 (.Y (
             L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_9), .A0 (nx8094), .A1 (
             nx4412)) ;
    inv01 ix4411 (.Y (nx4412), .A (L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_10)
          ) ;
    nor02_2x L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix93 (.Y (
             L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_10), .A0 (nx8094), .A1 (
             nx4414)) ;
    inv01 ix4413 (.Y (nx4414), .A (L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_11)
          ) ;
    nor02_2x L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix97 (.Y (
             L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_11), .A0 (nx8094), .A1 (
             nx4416)) ;
    inv01 ix4415 (.Y (nx4416), .A (L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_12)
          ) ;
    nor02_2x L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix101 (.Y (
             L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_12), .A0 (nx8094), .A1 (
             nx4418)) ;
    inv01 ix4417 (.Y (nx4418), .A (L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_13)
          ) ;
    nor02_2x L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix105 (.Y (
             L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_13), .A0 (nx8094), .A1 (
             nx4420)) ;
    inv01 ix4419 (.Y (nx4420), .A (L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_14)
          ) ;
    nor02_2x L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix109 (.Y (
             L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_14), .A0 (nx8096), .A1 (
             nx4422)) ;
    inv01 ix4421 (.Y (nx4422), .A (L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_15)
          ) ;
    nor02_2x L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix113 (.Y (
             L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_15), .A0 (nx8096), .A1 (
             nx4424)) ;
    inv01 ix4423 (.Y (nx4424), .A (L1_2_L2_2_G1_MINI_ALU_BoothPBeforeShift_16)
          ) ;
    nor02_2x L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix117 (.Y (
             L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_16), .A0 (nx8096), .A1 (
             nx4424)) ;
    mux21 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix189 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BoothOperand_0), .A0 (nx4426), .A1 (nx4428), .S0 (
          nx8084)) ;
    inv01 ix4425 (.Y (nx4426), .A (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_0)) ;
    inv01 ix4427 (.Y (nx4428), .A (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_0)) ;
    mux21 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix197 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BoothOperand_1), .A0 (nx4430), .A1 (nx4432), .S0 (
          nx8084)) ;
    inv01 ix4429 (.Y (nx4430), .A (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_1)) ;
    inv01 ix4431 (.Y (nx4432), .A (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_1)) ;
    mux21 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix205 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BoothOperand_2), .A0 (nx4434), .A1 (nx4436), .S0 (
          nx8084)) ;
    inv01 ix4433 (.Y (nx4434), .A (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_2)) ;
    inv01 ix4435 (.Y (nx4436), .A (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_2)) ;
    mux21 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix213 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BoothOperand_3), .A0 (nx4438), .A1 (nx4440), .S0 (
          nx8084)) ;
    inv01 ix4437 (.Y (nx4438), .A (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_3)) ;
    inv01 ix4439 (.Y (nx4440), .A (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_3)) ;
    mux21 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix221 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BoothOperand_4), .A0 (nx4442), .A1 (nx4444), .S0 (
          nx8084)) ;
    inv01 ix4441 (.Y (nx4442), .A (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_4)) ;
    inv01 ix4443 (.Y (nx4444), .A (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_4)) ;
    mux21 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix229 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BoothOperand_5), .A0 (nx4446), .A1 (nx4448), .S0 (
          nx8086)) ;
    inv01 ix4445 (.Y (nx4446), .A (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_5)) ;
    inv01 ix4447 (.Y (nx4448), .A (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_5)) ;
    mux21 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix237 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BoothOperand_6), .A0 (nx4450), .A1 (nx4452), .S0 (
          nx8086)) ;
    inv01 ix4449 (.Y (nx4450), .A (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_6)) ;
    inv01 ix4451 (.Y (nx4452), .A (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_6)) ;
    mux21 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix245 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BoothOperand_7), .A0 (nx4454), .A1 (nx4456), .S0 (
          nx8086)) ;
    inv01 ix4453 (.Y (nx4454), .A (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_7)) ;
    inv01 ix4455 (.Y (nx4456), .A (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_7)) ;
    mux21 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix253 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BoothOperand_8), .A0 (nx4458), .A1 (nx4460), .S0 (
          nx8086)) ;
    inv01 ix4457 (.Y (nx4458), .A (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_8)) ;
    inv01 ix4459 (.Y (nx4460), .A (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_8)) ;
    mux21 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix261 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BoothOperand_9), .A0 (nx4462), .A1 (nx4464), .S0 (
          nx8086)) ;
    inv01 ix4461 (.Y (nx4462), .A (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_9)) ;
    inv01 ix4463 (.Y (nx4464), .A (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_9)) ;
    mux21 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix269 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BoothOperand_10), .A0 (nx4466), .A1 (nx4468), .S0 (
          nx8086)) ;
    inv01 ix4465 (.Y (nx4466), .A (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_10)) ;
    inv01 ix4467 (.Y (nx4468), .A (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_10)) ;
    mux21 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix277 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BoothOperand_11), .A0 (nx4470), .A1 (nx4472), .S0 (
          nx8086)) ;
    inv01 ix4469 (.Y (nx4470), .A (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_11)) ;
    inv01 ix4471 (.Y (nx4472), .A (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_11)) ;
    mux21 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix285 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BoothOperand_12), .A0 (nx4474), .A1 (nx4476), .S0 (
          nx8088)) ;
    inv01 ix4473 (.Y (nx4474), .A (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_12)) ;
    inv01 ix4475 (.Y (nx4476), .A (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_12)) ;
    mux21 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix293 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BoothOperand_13), .A0 (nx4478), .A1 (nx4480), .S0 (
          nx8088)) ;
    inv01 ix4477 (.Y (nx4478), .A (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_13)) ;
    inv01 ix4479 (.Y (nx4480), .A (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_13)) ;
    mux21 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix301 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BoothOperand_14), .A0 (nx4482), .A1 (nx4484), .S0 (
          nx8088)) ;
    inv01 ix4481 (.Y (nx4482), .A (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_14)) ;
    inv01 ix4483 (.Y (nx4484), .A (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_14)) ;
    mux21 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix309 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BoothOperand_15), .A0 (nx4486), .A1 (nx4488), .S0 (
          nx8088)) ;
    inv01 ix4485 (.Y (nx4486), .A (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_15)) ;
    inv01 ix4487 (.Y (nx4488), .A (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_15)) ;
    mux21 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix317 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BoothOperand_16), .A0 (nx4490), .A1 (nx4492), .S0 (
          nx8088)) ;
    inv01 ix4489 (.Y (nx4490), .A (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDout_16)) ;
    inv01 ix4491 (.Y (nx4492), .A (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterADout_16)) ;
    xnor2 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_ix321 (.Y (
          L1_2_L2_2_G1_MINI_ALU_AddPToBoothOperand), .A0 (nx8088), .A1 (nx4358)
          ) ;
    oai32 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix393 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .A0 (nx8668), .A1 (
          RST), .A2 (nx8098), .B0 (nx4428), .B1 (nx4496)) ;
    oai32 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix403 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .A0 (nx8668), .A1 (
          RST), .A2 (nx8098), .B0 (nx4432), .B1 (nx4496)) ;
    oai32 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix413 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .A0 (nx8668), .A1 (
          RST), .A2 (nx8098), .B0 (nx4436), .B1 (nx4496)) ;
    oai32 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix423 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .A0 (nx8668), .A1 (
          RST), .A2 (nx8098), .B0 (nx4440), .B1 (nx4496)) ;
    oai32 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix433 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .A0 (nx8668), .A1 (
          RST), .A2 (nx8098), .B0 (nx4444), .B1 (nx4496)) ;
    oai32 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix443 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .A0 (nx8668), .A1 (
          RST), .A2 (nx8098), .B0 (nx4448), .B1 (nx4496)) ;
    oai32 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix453 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .A0 (nx8668), .A1 (
          RST), .A2 (nx8100), .B0 (nx4452), .B1 (nx4496)) ;
    oai32 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix463 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .A0 (nx8670), .A1 (
          RST), .A2 (nx8100), .B0 (nx4456), .B1 (nx4498)) ;
    oai32 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix473 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .A0 (nx8670), .A1 (
          RST), .A2 (nx8100), .B0 (nx4460), .B1 (nx4498)) ;
    oai32 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix483 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .A0 (nx4500), .A1 (
          RST), .A2 (nx8100), .B0 (nx4464), .B1 (nx4498)) ;
    inv01 ix4499 (.Y (nx4500), .A (FilterDin_2__2__0)) ;
    oai32 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix493 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .A0 (nx4502), .A1 (
          RST), .A2 (nx8100), .B0 (nx4468), .B1 (nx4498)) ;
    inv01 ix4501 (.Y (nx4502), .A (FilterDin_2__2__1)) ;
    oai32 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix503 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .A0 (nx4504), .A1 (
          RST), .A2 (nx8100), .B0 (nx4472), .B1 (nx4498)) ;
    inv01 ix4503 (.Y (nx4504), .A (FilterDin_2__2__2)) ;
    oai32 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix513 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .A0 (nx4506), .A1 (
          RST), .A2 (nx8100), .B0 (nx4476), .B1 (nx4498)) ;
    inv01 ix4505 (.Y (nx4506), .A (FilterDin_2__2__3)) ;
    oai32 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix523 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .A0 (nx4508), .A1 (
          RST), .A2 (nx8102), .B0 (nx4480), .B1 (nx4498)) ;
    inv01 ix4507 (.Y (nx4508), .A (FilterDin_2__2__4)) ;
    oai32 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix533 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .A0 (nx4510), .A1 (
          RST), .A2 (nx8102), .B0 (nx4484), .B1 (nx4512)) ;
    inv01 ix4509 (.Y (nx4510), .A (FilterDin_2__2__5)) ;
    inv01 ix4511 (.Y (nx4512), .A (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566)) ;
    oai32 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix543 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .A0 (nx4514), .A1 (
          RST), .A2 (nx8102), .B0 (nx4488), .B1 (nx4512)) ;
    inv01 ix4513 (.Y (nx4514), .A (FilterDin_2__2__6)) ;
    oai32 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix553 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .A0 (nx4516), .A1 (
          RST), .A2 (nx8102), .B0 (nx4492), .B1 (nx4512)) ;
    inv01 ix4515 (.Y (nx4516), .A (FilterDin_2__2__7)) ;
    nand02_2x L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix633 (.Y (nx4496), .A0 (
              nx7596), .A1 (nx8102)) ;
    nand02_2x L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix635 (.Y (nx4498), .A0 (
              nx7596), .A1 (nx8102)) ;
    oai32 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix393 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .A0 (nx8670), .A1 (
          RST), .A2 (nx8104), .B0 (nx4426), .B1 (nx4518)) ;
    oai32 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix403 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .A0 (nx8670), .A1 (
          RST), .A2 (nx8104), .B0 (nx4430), .B1 (nx4518)) ;
    oai32 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix413 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .A0 (nx8670), .A1 (
          RST), .A2 (nx8104), .B0 (nx4434), .B1 (nx4518)) ;
    oai32 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix423 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .A0 (nx8670), .A1 (
          RST), .A2 (nx8104), .B0 (nx4438), .B1 (nx4518)) ;
    oai32 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix433 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .A0 (nx8670), .A1 (
          RST), .A2 (nx8104), .B0 (nx4442), .B1 (nx4518)) ;
    oai32 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix443 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .A0 (nx8672), .A1 (
          RST), .A2 (nx8104), .B0 (nx4446), .B1 (nx4518)) ;
    oai32 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix453 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .A0 (nx8672), .A1 (
          RST), .A2 (nx8106), .B0 (nx4450), .B1 (nx4518)) ;
    oai32 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix463 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .A0 (nx8672), .A1 (
          RST), .A2 (nx8106), .B0 (nx4454), .B1 (nx4520)) ;
    oai32 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix473 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .A0 (nx8672), .A1 (
          RST), .A2 (nx8106), .B0 (nx4458), .B1 (nx4520)) ;
    oai32 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix483 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .A0 (nx4500), .A1 (
          RST), .A2 (nx8106), .B0 (nx4462), .B1 (nx4520)) ;
    oai32 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix493 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .A0 (nx4522), .A1 (
          RST), .A2 (nx8106), .B0 (nx4466), .B1 (nx4520)) ;
    inv01 ix4521 (.Y (nx4522), .A (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_10)) ;
    oai32 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix503 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .A0 (nx4524), .A1 (
          RST), .A2 (nx8106), .B0 (nx4470), .B1 (nx4520)) ;
    inv01 ix4523 (.Y (nx4524), .A (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_11)) ;
    oai32 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix513 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .A0 (nx4526), .A1 (
          RST), .A2 (nx8106), .B0 (nx4474), .B1 (nx4520)) ;
    inv01 ix4525 (.Y (nx4526), .A (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_12)) ;
    oai32 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix523 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .A0 (nx4528), .A1 (
          RST), .A2 (nx8108), .B0 (nx4478), .B1 (nx4520)) ;
    inv01 ix4527 (.Y (nx4528), .A (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_13)) ;
    oai32 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix533 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .A0 (nx4530), .A1 (
          RST), .A2 (nx8108), .B0 (nx4482), .B1 (nx4532)) ;
    inv01 ix4529 (.Y (nx4530), .A (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_14)) ;
    inv01 ix4531 (.Y (nx4532), .A (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566)) ;
    oai32 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix543 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .A0 (nx4534), .A1 (
          RST), .A2 (nx8108), .B0 (nx4486), .B1 (nx4532)) ;
    inv01 ix4533 (.Y (nx4534), .A (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_15)) ;
    oai32 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix553 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .A0 (nx4536), .A1 (
          RST), .A2 (nx8108), .B0 (nx4490), .B1 (nx4532)) ;
    inv01 ix4535 (.Y (nx4536), .A (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterSDin_16)) ;
    nand02_2x L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix633 (.Y (nx4518), .A0 (
              nx7596), .A1 (nx8108)) ;
    nand02_2x L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix635 (.Y (nx4520), .A0 (
              nx7596), .A1 (nx8108)) ;
    oai32 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix393 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .A0 (nx4538), .A1 (
          RST), .A2 (nx8110), .B0 (L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx384), .B1 (
          nx4540)) ;
    inv01 ix4537 (.Y (nx4538), .A (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_0)) ;
    oai32 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix403 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .A0 (nx4542), .A1 (
          RST), .A2 (nx8110), .B0 (nx4358), .B1 (nx4540)) ;
    inv01 ix4541 (.Y (nx4542), .A (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_1)) ;
    oai32 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix413 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .A0 (nx4544), .A1 (
          RST), .A2 (nx8110), .B0 (L1_2_L2_2_G1_MINI_ALU_nx387), .B1 (nx4540)) ;
    inv01 ix4543 (.Y (nx4544), .A (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_2)) ;
    oai32 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix423 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .A0 (nx4546), .A1 (
          RST), .A2 (nx8110), .B0 (L1_2_L2_2_G1_MINI_ALU_nx399), .B1 (nx4540)) ;
    inv01 ix4545 (.Y (nx4546), .A (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_3)) ;
    oai32 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix433 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .A0 (nx4548), .A1 (
          RST), .A2 (nx8110), .B0 (L1_2_L2_2_G1_MINI_ALU_nx409), .B1 (nx4540)) ;
    inv01 ix4547 (.Y (nx4548), .A (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_4)) ;
    oai32 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix443 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .A0 (nx4550), .A1 (
          RST), .A2 (nx8110), .B0 (L1_2_L2_2_G1_MINI_ALU_nx419), .B1 (nx4540)) ;
    inv01 ix4549 (.Y (nx4550), .A (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_5)) ;
    oai32 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix453 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .A0 (nx4552), .A1 (
          RST), .A2 (nx8110), .B0 (L1_2_L2_2_G1_MINI_ALU_nx429), .B1 (nx4540)) ;
    inv01 ix4551 (.Y (nx4552), .A (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_6)) ;
    oai32 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix463 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .A0 (nx4554), .A1 (
          RST), .A2 (nx8112), .B0 (L1_2_L2_2_G1_MINI_ALU_nx439), .B1 (nx4556)) ;
    inv01 ix4553 (.Y (nx4554), .A (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_7)) ;
    oai32 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix473 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .A0 (nx4558), .A1 (
          RST), .A2 (nx8112), .B0 (L1_2_L2_2_G1_MINI_ALU_nx449), .B1 (nx4556)) ;
    inv01 ix4557 (.Y (nx4558), .A (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_8)) ;
    oai32 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix483 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .A0 (nx4560), .A1 (
          RST), .A2 (nx8112), .B0 (L1_2_L2_2_G1_MINI_ALU_nx469), .B1 (nx4556)) ;
    inv01 ix4559 (.Y (nx4560), .A (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_9)) ;
    oai32 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix493 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .A0 (nx4562), .A1 (
          RST), .A2 (nx8112), .B0 (L1_2_L2_2_G1_MINI_ALU_nx477), .B1 (nx4556)) ;
    inv01 ix4561 (.Y (nx4562), .A (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_10)) ;
    oai32 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix503 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .A0 (nx4564), .A1 (
          RST), .A2 (nx8112), .B0 (L1_2_L2_2_G1_MINI_ALU_nx485), .B1 (nx4556)) ;
    inv01 ix4563 (.Y (nx4564), .A (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_11)) ;
    oai32 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix513 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .A0 (nx4566), .A1 (
          RST), .A2 (nx8112), .B0 (L1_2_L2_2_G1_MINI_ALU_nx493), .B1 (nx4556)) ;
    inv01 ix4565 (.Y (nx4566), .A (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_12)) ;
    oai32 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix523 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .A0 (nx4568), .A1 (
          RST), .A2 (nx8112), .B0 (L1_2_L2_2_G1_MINI_ALU_nx501), .B1 (nx4556)) ;
    inv01 ix4567 (.Y (nx4568), .A (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_13)) ;
    oai32 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix533 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .A0 (nx4570), .A1 (
          RST), .A2 (nx8114), .B0 (L1_2_L2_2_G1_MINI_ALU_nx509), .B1 (nx4572)) ;
    inv01 ix4569 (.Y (nx4570), .A (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_14)) ;
    inv01 ix4571 (.Y (nx4572), .A (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566)) ;
    oai32 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix543 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .A0 (nx4574), .A1 (
          RST), .A2 (nx8114), .B0 (L1_2_L2_2_G1_MINI_ALU_nx517), .B1 (nx4572)) ;
    inv01 ix4573 (.Y (nx4574), .A (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_15)) ;
    oai32 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix553 (.Y (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .A0 (nx4576), .A1 (
          RST), .A2 (nx8114), .B0 (nx4374), .B1 (nx4572)) ;
    inv01 ix4575 (.Y (nx4576), .A (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_RegisterPDin_16)) ;
    nand02_2x L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix633 (.Y (nx4540), .A0 (
              nx7596), .A1 (nx8114)) ;
    nand02_2x L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix635 (.Y (nx4556), .A0 (
              nx7598), .A1 (nx8114)) ;
    mux21 L1_2_L2_3_G2_MINI_ALU_ix404 (.Y (L1_2_L2_3_G2_MINI_ALU_nx403), .A0 (
          nx4578), .A1 (L1_2_L2_3_G2_MINI_ALU_BoothP_2), .S0 (
          L1_2_L2_3_G2_MINI_ALU_nx395)) ;
    inv01 ix4577 (.Y (nx4578), .A (L1_2_L2_3_G2_MINI_ALU_nx391)) ;
    mux21 L1_2_L2_3_G2_MINI_ALU_ix414 (.Y (L1_2_L2_3_G2_MINI_ALU_nx413), .A0 (
          nx4580), .A1 (L1_2_L2_3_G2_MINI_ALU_BoothP_3), .S0 (
          L1_2_L2_3_G2_MINI_ALU_nx405)) ;
    inv01 ix4579 (.Y (nx4580), .A (L1_2_L2_3_G2_MINI_ALU_nx403)) ;
    mux21 L1_2_L2_3_G2_MINI_ALU_ix424 (.Y (L1_2_L2_3_G2_MINI_ALU_nx423), .A0 (
          nx4582), .A1 (L1_2_L2_3_G2_MINI_ALU_BoothP_4), .S0 (
          L1_2_L2_3_G2_MINI_ALU_nx415)) ;
    inv01 ix4581 (.Y (nx4582), .A (L1_2_L2_3_G2_MINI_ALU_nx413)) ;
    mux21 L1_2_L2_3_G2_MINI_ALU_ix434 (.Y (L1_2_L2_3_G2_MINI_ALU_nx433), .A0 (
          nx4584), .A1 (L1_2_L2_3_G2_MINI_ALU_BoothP_5), .S0 (
          L1_2_L2_3_G2_MINI_ALU_nx425)) ;
    inv01 ix4583 (.Y (nx4584), .A (L1_2_L2_3_G2_MINI_ALU_nx423)) ;
    mux21 L1_2_L2_3_G2_MINI_ALU_ix444 (.Y (L1_2_L2_3_G2_MINI_ALU_nx443), .A0 (
          nx4586), .A1 (L1_2_L2_3_G2_MINI_ALU_BoothP_6), .S0 (
          L1_2_L2_3_G2_MINI_ALU_nx435)) ;
    inv01 ix4585 (.Y (nx4586), .A (L1_2_L2_3_G2_MINI_ALU_nx433)) ;
    mux21 L1_2_L2_3_G2_MINI_ALU_ix454 (.Y (L1_2_L2_3_G2_MINI_ALU_nx453), .A0 (
          nx4588), .A1 (L1_2_L2_3_G2_MINI_ALU_BoothP_7), .S0 (
          L1_2_L2_3_G2_MINI_ALU_nx445)) ;
    inv01 ix4587 (.Y (nx4588), .A (L1_2_L2_3_G2_MINI_ALU_nx443)) ;
    mux21 L1_2_L2_3_G2_MINI_ALU_ix462 (.Y (L1_2_L2_3_G2_MINI_ALU_nx461), .A0 (
          nx4590), .A1 (L1_2_L2_3_G2_MINI_ALU_BoothP_8), .S0 (
          L1_2_L2_3_G2_MINI_ALU_nx455)) ;
    inv01 ix4589 (.Y (nx4590), .A (L1_2_L2_3_G2_MINI_ALU_nx453)) ;
    mux21 L1_2_L2_3_G2_MINI_ALU_ix468 (.Y (L1_2_L2_3_G2_MINI_ALU_nx467), .A0 (
          nx4592), .A1 (L1_2_L2_3_G2_MINI_ALU_BoothP_9), .S0 (
          L1_2_L2_3_G2_MINI_ALU_nx463)) ;
    inv01 ix4591 (.Y (nx4592), .A (L1_2_L2_3_G2_MINI_ALU_nx461)) ;
    mux21 L1_2_L2_3_G2_MINI_ALU_ix476 (.Y (L1_2_L2_3_G2_MINI_ALU_nx475), .A0 (
          nx4594), .A1 (L1_2_L2_3_G2_MINI_ALU_BoothP_10), .S0 (
          L1_2_L2_3_G2_MINI_ALU_nx471)) ;
    inv01 ix4593 (.Y (nx4594), .A (L1_2_L2_3_G2_MINI_ALU_nx467)) ;
    mux21 L1_2_L2_3_G2_MINI_ALU_ix484 (.Y (L1_2_L2_3_G2_MINI_ALU_nx483), .A0 (
          nx4596), .A1 (L1_2_L2_3_G2_MINI_ALU_BoothP_11), .S0 (
          L1_2_L2_3_G2_MINI_ALU_nx479)) ;
    inv01 ix4595 (.Y (nx4596), .A (L1_2_L2_3_G2_MINI_ALU_nx475)) ;
    mux21 L1_2_L2_3_G2_MINI_ALU_ix492 (.Y (L1_2_L2_3_G2_MINI_ALU_nx491), .A0 (
          nx4598), .A1 (L1_2_L2_3_G2_MINI_ALU_BoothP_12), .S0 (
          L1_2_L2_3_G2_MINI_ALU_nx487)) ;
    inv01 ix4597 (.Y (nx4598), .A (L1_2_L2_3_G2_MINI_ALU_nx483)) ;
    mux21 L1_2_L2_3_G2_MINI_ALU_ix500 (.Y (L1_2_L2_3_G2_MINI_ALU_nx499), .A0 (
          nx4600), .A1 (L1_2_L2_3_G2_MINI_ALU_BoothP_13), .S0 (
          L1_2_L2_3_G2_MINI_ALU_nx495)) ;
    inv01 ix4599 (.Y (nx4600), .A (L1_2_L2_3_G2_MINI_ALU_nx491)) ;
    mux21 L1_2_L2_3_G2_MINI_ALU_ix508 (.Y (L1_2_L2_3_G2_MINI_ALU_nx507), .A0 (
          nx4602), .A1 (L1_2_L2_3_G2_MINI_ALU_BoothP_14), .S0 (
          L1_2_L2_3_G2_MINI_ALU_nx503)) ;
    inv01 ix4601 (.Y (nx4602), .A (L1_2_L2_3_G2_MINI_ALU_nx499)) ;
    mux21 L1_2_L2_3_G2_MINI_ALU_ix516 (.Y (L1_2_L2_3_G2_MINI_ALU_nx515), .A0 (
          nx4604), .A1 (L1_2_L2_3_G2_MINI_ALU_BoothP_15), .S0 (
          L1_2_L2_3_G2_MINI_ALU_nx511)) ;
    inv01 ix4603 (.Y (nx4604), .A (L1_2_L2_3_G2_MINI_ALU_nx507)) ;
    mux21 L1_2_L2_3_G2_MINI_ALU_ix161 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_1), .A0 (nx4606), .A1 (
          L1_2_L2_3_G2_MINI_ALU_nx379), .S0 (nx8118)) ;
    inv01 ix4605 (.Y (nx4606), .A (L1_2_L2_3_G2_MINI_ALU_BoothP_1)) ;
    mux21 L1_2_L2_3_G2_MINI_ALU_ix181 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_2), .A0 (
          L1_2_L2_3_G2_MINI_ALU_nx387), .A1 (L1_2_L2_3_G2_MINI_ALU_nx389), .S0 (
          nx8118)) ;
    mux21 L1_2_L2_3_G2_MINI_ALU_ix201 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_3), .A0 (
          L1_2_L2_3_G2_MINI_ALU_nx399), .A1 (L1_2_L2_3_G2_MINI_ALU_nx401), .S0 (
          nx8118)) ;
    mux21 L1_2_L2_3_G2_MINI_ALU_ix221 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_4), .A0 (
          L1_2_L2_3_G2_MINI_ALU_nx409), .A1 (L1_2_L2_3_G2_MINI_ALU_nx411), .S0 (
          nx8118)) ;
    mux21 L1_2_L2_3_G2_MINI_ALU_ix241 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_5), .A0 (
          L1_2_L2_3_G2_MINI_ALU_nx419), .A1 (L1_2_L2_3_G2_MINI_ALU_nx421), .S0 (
          nx8118)) ;
    mux21 L1_2_L2_3_G2_MINI_ALU_ix261 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_6), .A0 (
          L1_2_L2_3_G2_MINI_ALU_nx429), .A1 (L1_2_L2_3_G2_MINI_ALU_nx431), .S0 (
          nx8118)) ;
    mux21 L1_2_L2_3_G2_MINI_ALU_ix281 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_7), .A0 (
          L1_2_L2_3_G2_MINI_ALU_nx439), .A1 (L1_2_L2_3_G2_MINI_ALU_nx441), .S0 (
          nx8118)) ;
    mux21 L1_2_L2_3_G2_MINI_ALU_ix301 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_8), .A0 (
          L1_2_L2_3_G2_MINI_ALU_nx449), .A1 (L1_2_L2_3_G2_MINI_ALU_nx451), .S0 (
          nx8120)) ;
    mux21 L1_2_L2_3_G2_MINI_ALU_ix321 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_9), .A0 (
          L1_2_L2_3_G2_MINI_ALU_nx469), .A1 (nx4608), .S0 (nx8120)) ;
    inv01 ix4607 (.Y (nx4608), .A (L1_2_L2_3_G2_MINI_ALU_nx316)) ;
    mux21 L1_2_L2_3_G2_MINI_ALU_ix341 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_10), .A0 (
          L1_2_L2_3_G2_MINI_ALU_nx477), .A1 (nx4610), .S0 (nx8120)) ;
    inv01 ix4609 (.Y (nx4610), .A (L1_2_L2_3_G2_MINI_ALU_nx336)) ;
    mux21 L1_2_L2_3_G2_MINI_ALU_ix361 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_11), .A0 (
          L1_2_L2_3_G2_MINI_ALU_nx485), .A1 (nx4612), .S0 (nx8120)) ;
    inv01 ix4611 (.Y (nx4612), .A (L1_2_L2_3_G2_MINI_ALU_nx356)) ;
    mux21 L1_2_L2_3_G2_MINI_ALU_ix381 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_12), .A0 (
          L1_2_L2_3_G2_MINI_ALU_nx493), .A1 (nx4614), .S0 (nx8120)) ;
    inv01 ix4613 (.Y (nx4614), .A (L1_2_L2_3_G2_MINI_ALU_nx376)) ;
    mux21 L1_2_L2_3_G2_MINI_ALU_ix401 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_13), .A0 (
          L1_2_L2_3_G2_MINI_ALU_nx501), .A1 (nx4616), .S0 (nx8120)) ;
    inv01 ix4615 (.Y (nx4616), .A (L1_2_L2_3_G2_MINI_ALU_nx396)) ;
    mux21 L1_2_L2_3_G2_MINI_ALU_ix421 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_14), .A0 (
          L1_2_L2_3_G2_MINI_ALU_nx509), .A1 (nx4618), .S0 (nx8120)) ;
    inv01 ix4617 (.Y (nx4618), .A (L1_2_L2_3_G2_MINI_ALU_nx416)) ;
    mux21 L1_2_L2_3_G2_MINI_ALU_ix441 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_15), .A0 (
          L1_2_L2_3_G2_MINI_ALU_nx517), .A1 (nx4620), .S0 (nx8122)) ;
    inv01 ix4619 (.Y (nx4620), .A (L1_2_L2_3_G2_MINI_ALU_nx436)) ;
    mux21 L1_2_L2_3_G2_MINI_ALU_ix461 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_16), .A0 (nx4622), .A1 (nx4624
          ), .S0 (nx8122)) ;
    inv01 ix4621 (.Y (nx4622), .A (L1_2_L2_3_G2_MINI_ALU_BoothP_16)) ;
    inv01 ix4623 (.Y (nx4624), .A (L1_2_L2_3_G2_MINI_ALU_nx456)) ;
    nor02_2x L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix319 (.Y (
             L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642), .A0 (Start), .A1 (
             CalculatingBooth_dup_1119)) ;
    nor02_2x L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix85 (.Y (
             L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_0), .A0 (nx8132), .A1 (
             nx4626)) ;
    inv01 ix4625 (.Y (nx4626), .A (L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_1)) ;
    mux21 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix125 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_1), .A0 (nx4628), .A1 (
          nx4630), .S0 (nx8132)) ;
    inv01 ix4627 (.Y (nx4628), .A (L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_2)) ;
    inv01 ix4629 (.Y (nx4630), .A (WindowDin_2__3__0)) ;
    mux21 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix133 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_2), .A0 (nx4632), .A1 (
          nx4634), .S0 (nx8132)) ;
    inv01 ix4631 (.Y (nx4632), .A (L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_3)) ;
    inv01 ix4633 (.Y (nx4634), .A (WindowDin_2__3__1)) ;
    mux21 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix141 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_3), .A0 (nx4636), .A1 (
          nx4638), .S0 (nx8132)) ;
    inv01 ix4635 (.Y (nx4636), .A (L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_4)) ;
    inv01 ix4637 (.Y (nx4638), .A (WindowDin_2__3__2)) ;
    mux21 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix149 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_4), .A0 (nx4640), .A1 (
          nx4642), .S0 (nx8132)) ;
    inv01 ix4639 (.Y (nx4640), .A (L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_5)) ;
    inv01 ix4641 (.Y (nx4642), .A (WindowDin_2__3__3)) ;
    mux21 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix157 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_5), .A0 (nx4644), .A1 (
          nx4646), .S0 (nx8132)) ;
    inv01 ix4643 (.Y (nx4644), .A (L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_6)) ;
    inv01 ix4645 (.Y (nx4646), .A (WindowDin_2__3__4)) ;
    mux21 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix165 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_6), .A0 (nx4648), .A1 (
          nx4650), .S0 (nx8132)) ;
    inv01 ix4647 (.Y (nx4648), .A (L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_7)) ;
    inv01 ix4649 (.Y (nx4650), .A (WindowDin_2__3__5)) ;
    mux21 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix173 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_7), .A0 (nx4652), .A1 (
          nx4654), .S0 (nx8134)) ;
    inv01 ix4651 (.Y (nx4652), .A (L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_8)) ;
    inv01 ix4653 (.Y (nx4654), .A (WindowDin_2__3__6)) ;
    mux21 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix181 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_8), .A0 (nx4656), .A1 (
          nx4658), .S0 (nx8134)) ;
    inv01 ix4655 (.Y (nx4656), .A (L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_9)) ;
    inv01 ix4657 (.Y (nx4658), .A (WindowDin_2__3__7)) ;
    nor02_2x L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix89 (.Y (
             L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_9), .A0 (nx8134), .A1 (
             nx4660)) ;
    inv01 ix4659 (.Y (nx4660), .A (L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_10)
          ) ;
    nor02_2x L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix93 (.Y (
             L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_10), .A0 (nx8134), .A1 (
             nx4662)) ;
    inv01 ix4661 (.Y (nx4662), .A (L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_11)
          ) ;
    nor02_2x L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix97 (.Y (
             L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_11), .A0 (nx8134), .A1 (
             nx4664)) ;
    inv01 ix4663 (.Y (nx4664), .A (L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_12)
          ) ;
    nor02_2x L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix101 (.Y (
             L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_12), .A0 (nx8134), .A1 (
             nx4666)) ;
    inv01 ix4665 (.Y (nx4666), .A (L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_13)
          ) ;
    nor02_2x L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix105 (.Y (
             L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_13), .A0 (nx8134), .A1 (
             nx4668)) ;
    inv01 ix4667 (.Y (nx4668), .A (L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_14)
          ) ;
    nor02_2x L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix109 (.Y (
             L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_14), .A0 (nx8136), .A1 (
             nx4670)) ;
    inv01 ix4669 (.Y (nx4670), .A (L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_15)
          ) ;
    nor02_2x L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix113 (.Y (
             L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_15), .A0 (nx8136), .A1 (
             nx4672)) ;
    inv01 ix4671 (.Y (nx4672), .A (L1_2_L2_3_G2_MINI_ALU_BoothPBeforeShift_16)
          ) ;
    nor02_2x L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix117 (.Y (
             L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_16), .A0 (nx8136), .A1 (
             nx4672)) ;
    mux21 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix189 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BoothOperand_0), .A0 (nx4674), .A1 (nx4676), .S0 (
          nx8124)) ;
    inv01 ix4673 (.Y (nx4674), .A (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_0)) ;
    inv01 ix4675 (.Y (nx4676), .A (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_0)) ;
    mux21 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix197 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BoothOperand_1), .A0 (nx4678), .A1 (nx4680), .S0 (
          nx8124)) ;
    inv01 ix4677 (.Y (nx4678), .A (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_1)) ;
    inv01 ix4679 (.Y (nx4680), .A (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_1)) ;
    mux21 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix205 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BoothOperand_2), .A0 (nx4682), .A1 (nx4684), .S0 (
          nx8124)) ;
    inv01 ix4681 (.Y (nx4682), .A (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_2)) ;
    inv01 ix4683 (.Y (nx4684), .A (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_2)) ;
    mux21 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix213 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BoothOperand_3), .A0 (nx4686), .A1 (nx4688), .S0 (
          nx8124)) ;
    inv01 ix4685 (.Y (nx4686), .A (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_3)) ;
    inv01 ix4687 (.Y (nx4688), .A (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_3)) ;
    mux21 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix221 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BoothOperand_4), .A0 (nx4690), .A1 (nx4692), .S0 (
          nx8124)) ;
    inv01 ix4689 (.Y (nx4690), .A (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_4)) ;
    inv01 ix4691 (.Y (nx4692), .A (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_4)) ;
    mux21 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix229 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BoothOperand_5), .A0 (nx4694), .A1 (nx4696), .S0 (
          nx8126)) ;
    inv01 ix4693 (.Y (nx4694), .A (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_5)) ;
    inv01 ix4695 (.Y (nx4696), .A (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_5)) ;
    mux21 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix237 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BoothOperand_6), .A0 (nx4698), .A1 (nx4700), .S0 (
          nx8126)) ;
    inv01 ix4697 (.Y (nx4698), .A (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_6)) ;
    inv01 ix4699 (.Y (nx4700), .A (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_6)) ;
    mux21 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix245 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BoothOperand_7), .A0 (nx4702), .A1 (nx4704), .S0 (
          nx8126)) ;
    inv01 ix4701 (.Y (nx4702), .A (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_7)) ;
    inv01 ix4703 (.Y (nx4704), .A (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_7)) ;
    mux21 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix253 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BoothOperand_8), .A0 (nx4706), .A1 (nx4708), .S0 (
          nx8126)) ;
    inv01 ix4705 (.Y (nx4706), .A (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_8)) ;
    inv01 ix4707 (.Y (nx4708), .A (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_8)) ;
    mux21 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix261 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BoothOperand_9), .A0 (nx4710), .A1 (nx4712), .S0 (
          nx8126)) ;
    inv01 ix4709 (.Y (nx4710), .A (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_9)) ;
    inv01 ix4711 (.Y (nx4712), .A (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_9)) ;
    mux21 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix269 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BoothOperand_10), .A0 (nx4714), .A1 (nx4716), .S0 (
          nx8126)) ;
    inv01 ix4713 (.Y (nx4714), .A (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_10)) ;
    inv01 ix4715 (.Y (nx4716), .A (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_10)) ;
    mux21 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix277 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BoothOperand_11), .A0 (nx4718), .A1 (nx4720), .S0 (
          nx8126)) ;
    inv01 ix4717 (.Y (nx4718), .A (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_11)) ;
    inv01 ix4719 (.Y (nx4720), .A (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_11)) ;
    mux21 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix285 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BoothOperand_12), .A0 (nx4722), .A1 (nx4724), .S0 (
          nx8128)) ;
    inv01 ix4721 (.Y (nx4722), .A (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_12)) ;
    inv01 ix4723 (.Y (nx4724), .A (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_12)) ;
    mux21 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix293 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BoothOperand_13), .A0 (nx4726), .A1 (nx4728), .S0 (
          nx8128)) ;
    inv01 ix4725 (.Y (nx4726), .A (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_13)) ;
    inv01 ix4727 (.Y (nx4728), .A (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_13)) ;
    mux21 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix301 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BoothOperand_14), .A0 (nx4730), .A1 (nx4732), .S0 (
          nx8128)) ;
    inv01 ix4729 (.Y (nx4730), .A (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_14)) ;
    inv01 ix4731 (.Y (nx4732), .A (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_14)) ;
    mux21 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix309 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BoothOperand_15), .A0 (nx4734), .A1 (nx4736), .S0 (
          nx8128)) ;
    inv01 ix4733 (.Y (nx4734), .A (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_15)) ;
    inv01 ix4735 (.Y (nx4736), .A (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_15)) ;
    mux21 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix317 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BoothOperand_16), .A0 (nx4738), .A1 (nx4740), .S0 (
          nx8128)) ;
    inv01 ix4737 (.Y (nx4738), .A (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_16)) ;
    inv01 ix4739 (.Y (nx4740), .A (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_16)) ;
    xnor2 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix321 (.Y (
          L1_2_L2_3_G2_MINI_ALU_AddPToBoothOperand), .A0 (nx8128), .A1 (nx4606)
          ) ;
    oai32 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix393 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .A0 (nx8674), .A1 (
          RST), .A2 (nx8138), .B0 (nx4676), .B1 (nx4744)) ;
    oai32 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix403 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .A0 (nx8674), .A1 (
          RST), .A2 (nx8138), .B0 (nx4680), .B1 (nx4744)) ;
    oai32 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix413 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .A0 (nx8674), .A1 (
          RST), .A2 (nx8138), .B0 (nx4684), .B1 (nx4744)) ;
    oai32 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix423 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .A0 (nx8674), .A1 (
          RST), .A2 (nx8138), .B0 (nx4688), .B1 (nx4744)) ;
    oai32 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix433 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .A0 (nx8674), .A1 (
          RST), .A2 (nx8138), .B0 (nx4692), .B1 (nx4744)) ;
    oai32 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix443 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .A0 (nx8674), .A1 (
          RST), .A2 (nx8138), .B0 (nx4696), .B1 (nx4744)) ;
    oai32 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix453 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .A0 (nx8674), .A1 (
          RST), .A2 (nx8140), .B0 (nx4700), .B1 (nx4744)) ;
    oai32 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix463 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .A0 (nx8676), .A1 (
          RST), .A2 (nx8140), .B0 (nx4704), .B1 (nx4746)) ;
    oai32 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix473 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .A0 (nx8676), .A1 (
          RST), .A2 (nx8140), .B0 (nx4708), .B1 (nx4746)) ;
    oai32 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix483 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .A0 (nx4748), .A1 (
          RST), .A2 (nx8140), .B0 (nx4712), .B1 (nx4746)) ;
    inv01 ix4747 (.Y (nx4748), .A (FilterDin_2__3__0)) ;
    oai32 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix493 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .A0 (nx4750), .A1 (
          RST), .A2 (nx8140), .B0 (nx4716), .B1 (nx4746)) ;
    inv01 ix4749 (.Y (nx4750), .A (FilterDin_2__3__1)) ;
    oai32 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix503 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .A0 (nx4752), .A1 (
          RST), .A2 (nx8140), .B0 (nx4720), .B1 (nx4746)) ;
    inv01 ix4751 (.Y (nx4752), .A (FilterDin_2__3__2)) ;
    oai32 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix513 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .A0 (nx4754), .A1 (
          RST), .A2 (nx8140), .B0 (nx4724), .B1 (nx4746)) ;
    inv01 ix4753 (.Y (nx4754), .A (FilterDin_2__3__3)) ;
    oai32 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix523 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .A0 (nx4756), .A1 (
          RST), .A2 (nx8142), .B0 (nx4728), .B1 (nx4746)) ;
    inv01 ix4755 (.Y (nx4756), .A (FilterDin_2__3__4)) ;
    oai32 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix533 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .A0 (nx4758), .A1 (
          RST), .A2 (nx8142), .B0 (nx4732), .B1 (nx4760)) ;
    inv01 ix4757 (.Y (nx4758), .A (FilterDin_2__3__5)) ;
    inv01 ix4759 (.Y (nx4760), .A (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566)) ;
    oai32 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix543 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .A0 (nx4762), .A1 (
          RST), .A2 (nx8142), .B0 (nx4736), .B1 (nx4760)) ;
    inv01 ix4761 (.Y (nx4762), .A (FilterDin_2__3__6)) ;
    oai32 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix553 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .A0 (nx4764), .A1 (
          RST), .A2 (nx8142), .B0 (nx4740), .B1 (nx4760)) ;
    inv01 ix4763 (.Y (nx4764), .A (FilterDin_2__3__7)) ;
    nand02_2x L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix633 (.Y (nx4744), .A0 (
              nx7598), .A1 (nx8142)) ;
    nand02_2x L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix635 (.Y (nx4746), .A0 (
              nx7598), .A1 (nx8142)) ;
    oai32 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix393 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .A0 (nx8676), .A1 (
          RST), .A2 (nx8144), .B0 (nx4674), .B1 (nx4766)) ;
    oai32 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix403 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .A0 (nx8676), .A1 (
          RST), .A2 (nx8144), .B0 (nx4678), .B1 (nx4766)) ;
    oai32 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix413 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .A0 (nx8676), .A1 (
          RST), .A2 (nx8144), .B0 (nx4682), .B1 (nx4766)) ;
    oai32 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix423 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .A0 (nx8676), .A1 (
          RST), .A2 (nx8144), .B0 (nx4686), .B1 (nx4766)) ;
    oai32 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix433 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .A0 (nx8676), .A1 (
          RST), .A2 (nx8144), .B0 (nx4690), .B1 (nx4766)) ;
    oai32 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix443 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .A0 (nx8678), .A1 (
          RST), .A2 (nx8144), .B0 (nx4694), .B1 (nx4766)) ;
    oai32 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix453 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .A0 (nx8678), .A1 (
          RST), .A2 (nx8146), .B0 (nx4698), .B1 (nx4766)) ;
    oai32 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix463 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .A0 (nx8678), .A1 (
          RST), .A2 (nx8146), .B0 (nx4702), .B1 (nx4768)) ;
    oai32 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix473 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .A0 (nx8678), .A1 (
          RST), .A2 (nx8146), .B0 (nx4706), .B1 (nx4768)) ;
    oai32 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix483 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .A0 (nx4748), .A1 (
          RST), .A2 (nx8146), .B0 (nx4710), .B1 (nx4768)) ;
    oai32 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix493 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .A0 (nx4770), .A1 (
          RST), .A2 (nx8146), .B0 (nx4714), .B1 (nx4768)) ;
    inv01 ix4769 (.Y (nx4770), .A (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_10)) ;
    oai32 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix503 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .A0 (nx4772), .A1 (
          RST), .A2 (nx8146), .B0 (nx4718), .B1 (nx4768)) ;
    inv01 ix4771 (.Y (nx4772), .A (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_11)) ;
    oai32 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix513 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .A0 (nx4774), .A1 (
          RST), .A2 (nx8146), .B0 (nx4722), .B1 (nx4768)) ;
    inv01 ix4773 (.Y (nx4774), .A (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_12)) ;
    oai32 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix523 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .A0 (nx4776), .A1 (
          RST), .A2 (nx8148), .B0 (nx4726), .B1 (nx4768)) ;
    inv01 ix4775 (.Y (nx4776), .A (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_13)) ;
    oai32 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix533 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .A0 (nx4778), .A1 (
          RST), .A2 (nx8148), .B0 (nx4730), .B1 (nx4780)) ;
    inv01 ix4777 (.Y (nx4778), .A (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_14)) ;
    inv01 ix4779 (.Y (nx4780), .A (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566)) ;
    oai32 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix543 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .A0 (nx4782), .A1 (
          RST), .A2 (nx8148), .B0 (nx4734), .B1 (nx4780)) ;
    inv01 ix4781 (.Y (nx4782), .A (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_15)) ;
    oai32 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix553 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .A0 (nx4784), .A1 (
          RST), .A2 (nx8148), .B0 (nx4738), .B1 (nx4780)) ;
    inv01 ix4783 (.Y (nx4784), .A (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_16)) ;
    nand02_2x L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix633 (.Y (nx4766), .A0 (
              nx7598), .A1 (nx8148)) ;
    nand02_2x L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix635 (.Y (nx4768), .A0 (
              nx7598), .A1 (nx8148)) ;
    oai32 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix393 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .A0 (nx4786), .A1 (
          RST), .A2 (nx8150), .B0 (L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx384), .B1 (
          nx4788)) ;
    inv01 ix4785 (.Y (nx4786), .A (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_0)) ;
    oai32 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix403 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .A0 (nx4790), .A1 (
          RST), .A2 (nx8150), .B0 (nx4606), .B1 (nx4788)) ;
    inv01 ix4789 (.Y (nx4790), .A (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_1)) ;
    oai32 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix413 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .A0 (nx4792), .A1 (
          RST), .A2 (nx8150), .B0 (L1_2_L2_3_G2_MINI_ALU_nx387), .B1 (nx4788)) ;
    inv01 ix4791 (.Y (nx4792), .A (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_2)) ;
    oai32 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix423 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .A0 (nx4794), .A1 (
          RST), .A2 (nx8150), .B0 (L1_2_L2_3_G2_MINI_ALU_nx399), .B1 (nx4788)) ;
    inv01 ix4793 (.Y (nx4794), .A (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_3)) ;
    oai32 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix433 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .A0 (nx4796), .A1 (
          RST), .A2 (nx8150), .B0 (L1_2_L2_3_G2_MINI_ALU_nx409), .B1 (nx4788)) ;
    inv01 ix4795 (.Y (nx4796), .A (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_4)) ;
    oai32 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix443 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .A0 (nx4798), .A1 (
          RST), .A2 (nx8150), .B0 (L1_2_L2_3_G2_MINI_ALU_nx419), .B1 (nx4788)) ;
    inv01 ix4797 (.Y (nx4798), .A (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_5)) ;
    oai32 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix453 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .A0 (nx4800), .A1 (
          RST), .A2 (nx8150), .B0 (L1_2_L2_3_G2_MINI_ALU_nx429), .B1 (nx4788)) ;
    inv01 ix4799 (.Y (nx4800), .A (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_6)) ;
    oai32 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix463 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .A0 (nx4802), .A1 (
          RST), .A2 (nx8152), .B0 (L1_2_L2_3_G2_MINI_ALU_nx439), .B1 (nx4804)) ;
    inv01 ix4801 (.Y (nx4802), .A (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_7)) ;
    oai32 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix473 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .A0 (nx4806), .A1 (
          RST), .A2 (nx8152), .B0 (L1_2_L2_3_G2_MINI_ALU_nx449), .B1 (nx4804)) ;
    inv01 ix4805 (.Y (nx4806), .A (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_8)) ;
    oai32 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix483 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .A0 (nx4808), .A1 (
          RST), .A2 (nx8152), .B0 (L1_2_L2_3_G2_MINI_ALU_nx469), .B1 (nx4804)) ;
    inv01 ix4807 (.Y (nx4808), .A (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_9)) ;
    oai32 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix493 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .A0 (nx4810), .A1 (
          RST), .A2 (nx8152), .B0 (L1_2_L2_3_G2_MINI_ALU_nx477), .B1 (nx4804)) ;
    inv01 ix4809 (.Y (nx4810), .A (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_10)) ;
    oai32 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix503 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .A0 (nx4812), .A1 (
          RST), .A2 (nx8152), .B0 (L1_2_L2_3_G2_MINI_ALU_nx485), .B1 (nx4804)) ;
    inv01 ix4811 (.Y (nx4812), .A (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_11)) ;
    oai32 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix513 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .A0 (nx4814), .A1 (
          RST), .A2 (nx8152), .B0 (L1_2_L2_3_G2_MINI_ALU_nx493), .B1 (nx4804)) ;
    inv01 ix4813 (.Y (nx4814), .A (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_12)) ;
    oai32 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix523 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .A0 (nx4816), .A1 (
          RST), .A2 (nx8152), .B0 (L1_2_L2_3_G2_MINI_ALU_nx501), .B1 (nx4804)) ;
    inv01 ix4815 (.Y (nx4816), .A (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_13)) ;
    oai32 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix533 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .A0 (nx4818), .A1 (
          RST), .A2 (nx8154), .B0 (L1_2_L2_3_G2_MINI_ALU_nx509), .B1 (nx4820)) ;
    inv01 ix4817 (.Y (nx4818), .A (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_14)) ;
    inv01 ix4819 (.Y (nx4820), .A (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566)) ;
    oai32 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix543 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .A0 (nx4822), .A1 (
          RST), .A2 (nx8154), .B0 (L1_2_L2_3_G2_MINI_ALU_nx517), .B1 (nx4820)) ;
    inv01 ix4821 (.Y (nx4822), .A (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_15)) ;
    oai32 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix553 (.Y (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .A0 (nx4824), .A1 (
          RST), .A2 (nx8154), .B0 (nx4622), .B1 (nx4820)) ;
    inv01 ix4823 (.Y (nx4824), .A (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_16)) ;
    nand02_2x L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix633 (.Y (nx4788), .A0 (
              nx7598), .A1 (nx8154)) ;
    nand02_2x L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix635 (.Y (nx4804), .A0 (
              nx7598), .A1 (nx8154)) ;
    mux21 L1_2_L2_4_G2_MINI_ALU_ix404 (.Y (L1_2_L2_4_G2_MINI_ALU_nx403), .A0 (
          nx4826), .A1 (L1_2_L2_4_G2_MINI_ALU_BoothP_2), .S0 (
          L1_2_L2_4_G2_MINI_ALU_nx395)) ;
    inv01 ix4825 (.Y (nx4826), .A (L1_2_L2_4_G2_MINI_ALU_nx391)) ;
    mux21 L1_2_L2_4_G2_MINI_ALU_ix414 (.Y (L1_2_L2_4_G2_MINI_ALU_nx413), .A0 (
          nx4828), .A1 (L1_2_L2_4_G2_MINI_ALU_BoothP_3), .S0 (
          L1_2_L2_4_G2_MINI_ALU_nx405)) ;
    inv01 ix4827 (.Y (nx4828), .A (L1_2_L2_4_G2_MINI_ALU_nx403)) ;
    mux21 L1_2_L2_4_G2_MINI_ALU_ix424 (.Y (L1_2_L2_4_G2_MINI_ALU_nx423), .A0 (
          nx4830), .A1 (L1_2_L2_4_G2_MINI_ALU_BoothP_4), .S0 (
          L1_2_L2_4_G2_MINI_ALU_nx415)) ;
    inv01 ix4829 (.Y (nx4830), .A (L1_2_L2_4_G2_MINI_ALU_nx413)) ;
    mux21 L1_2_L2_4_G2_MINI_ALU_ix434 (.Y (L1_2_L2_4_G2_MINI_ALU_nx433), .A0 (
          nx4832), .A1 (L1_2_L2_4_G2_MINI_ALU_BoothP_5), .S0 (
          L1_2_L2_4_G2_MINI_ALU_nx425)) ;
    inv01 ix4831 (.Y (nx4832), .A (L1_2_L2_4_G2_MINI_ALU_nx423)) ;
    mux21 L1_2_L2_4_G2_MINI_ALU_ix444 (.Y (L1_2_L2_4_G2_MINI_ALU_nx443), .A0 (
          nx4834), .A1 (L1_2_L2_4_G2_MINI_ALU_BoothP_6), .S0 (
          L1_2_L2_4_G2_MINI_ALU_nx435)) ;
    inv01 ix4833 (.Y (nx4834), .A (L1_2_L2_4_G2_MINI_ALU_nx433)) ;
    mux21 L1_2_L2_4_G2_MINI_ALU_ix454 (.Y (L1_2_L2_4_G2_MINI_ALU_nx453), .A0 (
          nx4836), .A1 (L1_2_L2_4_G2_MINI_ALU_BoothP_7), .S0 (
          L1_2_L2_4_G2_MINI_ALU_nx445)) ;
    inv01 ix4835 (.Y (nx4836), .A (L1_2_L2_4_G2_MINI_ALU_nx443)) ;
    mux21 L1_2_L2_4_G2_MINI_ALU_ix462 (.Y (L1_2_L2_4_G2_MINI_ALU_nx461), .A0 (
          nx4838), .A1 (L1_2_L2_4_G2_MINI_ALU_BoothP_8), .S0 (
          L1_2_L2_4_G2_MINI_ALU_nx455)) ;
    inv01 ix4837 (.Y (nx4838), .A (L1_2_L2_4_G2_MINI_ALU_nx453)) ;
    mux21 L1_2_L2_4_G2_MINI_ALU_ix468 (.Y (L1_2_L2_4_G2_MINI_ALU_nx467), .A0 (
          nx4840), .A1 (L1_2_L2_4_G2_MINI_ALU_BoothP_9), .S0 (
          L1_2_L2_4_G2_MINI_ALU_nx463)) ;
    inv01 ix4839 (.Y (nx4840), .A (L1_2_L2_4_G2_MINI_ALU_nx461)) ;
    mux21 L1_2_L2_4_G2_MINI_ALU_ix476 (.Y (L1_2_L2_4_G2_MINI_ALU_nx475), .A0 (
          nx4842), .A1 (L1_2_L2_4_G2_MINI_ALU_BoothP_10), .S0 (
          L1_2_L2_4_G2_MINI_ALU_nx471)) ;
    inv01 ix4841 (.Y (nx4842), .A (L1_2_L2_4_G2_MINI_ALU_nx467)) ;
    mux21 L1_2_L2_4_G2_MINI_ALU_ix484 (.Y (L1_2_L2_4_G2_MINI_ALU_nx483), .A0 (
          nx4844), .A1 (L1_2_L2_4_G2_MINI_ALU_BoothP_11), .S0 (
          L1_2_L2_4_G2_MINI_ALU_nx479)) ;
    inv01 ix4843 (.Y (nx4844), .A (L1_2_L2_4_G2_MINI_ALU_nx475)) ;
    mux21 L1_2_L2_4_G2_MINI_ALU_ix492 (.Y (L1_2_L2_4_G2_MINI_ALU_nx491), .A0 (
          nx4846), .A1 (L1_2_L2_4_G2_MINI_ALU_BoothP_12), .S0 (
          L1_2_L2_4_G2_MINI_ALU_nx487)) ;
    inv01 ix4845 (.Y (nx4846), .A (L1_2_L2_4_G2_MINI_ALU_nx483)) ;
    mux21 L1_2_L2_4_G2_MINI_ALU_ix500 (.Y (L1_2_L2_4_G2_MINI_ALU_nx499), .A0 (
          nx4848), .A1 (L1_2_L2_4_G2_MINI_ALU_BoothP_13), .S0 (
          L1_2_L2_4_G2_MINI_ALU_nx495)) ;
    inv01 ix4847 (.Y (nx4848), .A (L1_2_L2_4_G2_MINI_ALU_nx491)) ;
    mux21 L1_2_L2_4_G2_MINI_ALU_ix508 (.Y (L1_2_L2_4_G2_MINI_ALU_nx507), .A0 (
          nx4850), .A1 (L1_2_L2_4_G2_MINI_ALU_BoothP_14), .S0 (
          L1_2_L2_4_G2_MINI_ALU_nx503)) ;
    inv01 ix4849 (.Y (nx4850), .A (L1_2_L2_4_G2_MINI_ALU_nx499)) ;
    mux21 L1_2_L2_4_G2_MINI_ALU_ix516 (.Y (L1_2_L2_4_G2_MINI_ALU_nx515), .A0 (
          nx4852), .A1 (L1_2_L2_4_G2_MINI_ALU_BoothP_15), .S0 (
          L1_2_L2_4_G2_MINI_ALU_nx511)) ;
    inv01 ix4851 (.Y (nx4852), .A (L1_2_L2_4_G2_MINI_ALU_nx507)) ;
    mux21 L1_2_L2_4_G2_MINI_ALU_ix161 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_1), .A0 (nx4854), .A1 (
          L1_2_L2_4_G2_MINI_ALU_nx379), .S0 (nx8158)) ;
    inv01 ix4853 (.Y (nx4854), .A (L1_2_L2_4_G2_MINI_ALU_BoothP_1)) ;
    mux21 L1_2_L2_4_G2_MINI_ALU_ix181 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_2), .A0 (
          L1_2_L2_4_G2_MINI_ALU_nx387), .A1 (L1_2_L2_4_G2_MINI_ALU_nx389), .S0 (
          nx8158)) ;
    mux21 L1_2_L2_4_G2_MINI_ALU_ix201 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_3), .A0 (
          L1_2_L2_4_G2_MINI_ALU_nx399), .A1 (L1_2_L2_4_G2_MINI_ALU_nx401), .S0 (
          nx8158)) ;
    mux21 L1_2_L2_4_G2_MINI_ALU_ix221 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_4), .A0 (
          L1_2_L2_4_G2_MINI_ALU_nx409), .A1 (L1_2_L2_4_G2_MINI_ALU_nx411), .S0 (
          nx8158)) ;
    mux21 L1_2_L2_4_G2_MINI_ALU_ix241 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_5), .A0 (
          L1_2_L2_4_G2_MINI_ALU_nx419), .A1 (L1_2_L2_4_G2_MINI_ALU_nx421), .S0 (
          nx8158)) ;
    mux21 L1_2_L2_4_G2_MINI_ALU_ix261 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_6), .A0 (
          L1_2_L2_4_G2_MINI_ALU_nx429), .A1 (L1_2_L2_4_G2_MINI_ALU_nx431), .S0 (
          nx8158)) ;
    mux21 L1_2_L2_4_G2_MINI_ALU_ix281 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_7), .A0 (
          L1_2_L2_4_G2_MINI_ALU_nx439), .A1 (L1_2_L2_4_G2_MINI_ALU_nx441), .S0 (
          nx8158)) ;
    mux21 L1_2_L2_4_G2_MINI_ALU_ix301 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_8), .A0 (
          L1_2_L2_4_G2_MINI_ALU_nx449), .A1 (L1_2_L2_4_G2_MINI_ALU_nx451), .S0 (
          nx8160)) ;
    mux21 L1_2_L2_4_G2_MINI_ALU_ix321 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_9), .A0 (
          L1_2_L2_4_G2_MINI_ALU_nx469), .A1 (nx4856), .S0 (nx8160)) ;
    inv01 ix4855 (.Y (nx4856), .A (L1_2_L2_4_G2_MINI_ALU_nx316)) ;
    mux21 L1_2_L2_4_G2_MINI_ALU_ix341 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_10), .A0 (
          L1_2_L2_4_G2_MINI_ALU_nx477), .A1 (nx4858), .S0 (nx8160)) ;
    inv01 ix4857 (.Y (nx4858), .A (L1_2_L2_4_G2_MINI_ALU_nx336)) ;
    mux21 L1_2_L2_4_G2_MINI_ALU_ix361 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_11), .A0 (
          L1_2_L2_4_G2_MINI_ALU_nx485), .A1 (nx4860), .S0 (nx8160)) ;
    inv01 ix4859 (.Y (nx4860), .A (L1_2_L2_4_G2_MINI_ALU_nx356)) ;
    mux21 L1_2_L2_4_G2_MINI_ALU_ix381 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_12), .A0 (
          L1_2_L2_4_G2_MINI_ALU_nx493), .A1 (nx4862), .S0 (nx8160)) ;
    inv01 ix4861 (.Y (nx4862), .A (L1_2_L2_4_G2_MINI_ALU_nx376)) ;
    mux21 L1_2_L2_4_G2_MINI_ALU_ix401 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_13), .A0 (
          L1_2_L2_4_G2_MINI_ALU_nx501), .A1 (nx4864), .S0 (nx8160)) ;
    inv01 ix4863 (.Y (nx4864), .A (L1_2_L2_4_G2_MINI_ALU_nx396)) ;
    mux21 L1_2_L2_4_G2_MINI_ALU_ix421 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_14), .A0 (
          L1_2_L2_4_G2_MINI_ALU_nx509), .A1 (nx4866), .S0 (nx8160)) ;
    inv01 ix4865 (.Y (nx4866), .A (L1_2_L2_4_G2_MINI_ALU_nx416)) ;
    mux21 L1_2_L2_4_G2_MINI_ALU_ix441 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_15), .A0 (
          L1_2_L2_4_G2_MINI_ALU_nx517), .A1 (nx4868), .S0 (nx8162)) ;
    inv01 ix4867 (.Y (nx4868), .A (L1_2_L2_4_G2_MINI_ALU_nx436)) ;
    mux21 L1_2_L2_4_G2_MINI_ALU_ix461 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_16), .A0 (nx4870), .A1 (nx4872
          ), .S0 (nx8162)) ;
    inv01 ix4869 (.Y (nx4870), .A (L1_2_L2_4_G2_MINI_ALU_BoothP_16)) ;
    inv01 ix4871 (.Y (nx4872), .A (L1_2_L2_4_G2_MINI_ALU_nx456)) ;
    nor02_2x L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix319 (.Y (
             L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642), .A0 (Start), .A1 (
             CalculatingBooth_dup_1162)) ;
    nor02_2x L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix85 (.Y (
             L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_0), .A0 (nx8172), .A1 (
             nx4874)) ;
    inv01 ix4873 (.Y (nx4874), .A (L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_1)) ;
    mux21 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix125 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_1), .A0 (nx4876), .A1 (
          nx4878), .S0 (nx8172)) ;
    inv01 ix4875 (.Y (nx4876), .A (L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_2)) ;
    inv01 ix4877 (.Y (nx4878), .A (WindowDin_2__4__0)) ;
    mux21 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix133 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_2), .A0 (nx4880), .A1 (
          nx4882), .S0 (nx8172)) ;
    inv01 ix4879 (.Y (nx4880), .A (L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_3)) ;
    inv01 ix4881 (.Y (nx4882), .A (WindowDin_2__4__1)) ;
    mux21 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix141 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_3), .A0 (nx4884), .A1 (
          nx4886), .S0 (nx8172)) ;
    inv01 ix4883 (.Y (nx4884), .A (L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_4)) ;
    inv01 ix4885 (.Y (nx4886), .A (WindowDin_2__4__2)) ;
    mux21 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix149 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_4), .A0 (nx4888), .A1 (
          nx4890), .S0 (nx8172)) ;
    inv01 ix4887 (.Y (nx4888), .A (L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_5)) ;
    inv01 ix4889 (.Y (nx4890), .A (WindowDin_2__4__3)) ;
    mux21 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix157 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_5), .A0 (nx4892), .A1 (
          nx4894), .S0 (nx8172)) ;
    inv01 ix4891 (.Y (nx4892), .A (L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_6)) ;
    inv01 ix4893 (.Y (nx4894), .A (WindowDin_2__4__4)) ;
    mux21 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix165 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_6), .A0 (nx4896), .A1 (
          nx4898), .S0 (nx8172)) ;
    inv01 ix4895 (.Y (nx4896), .A (L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_7)) ;
    inv01 ix4897 (.Y (nx4898), .A (WindowDin_2__4__5)) ;
    mux21 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix173 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_7), .A0 (nx4900), .A1 (
          nx4902), .S0 (nx8174)) ;
    inv01 ix4899 (.Y (nx4900), .A (L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_8)) ;
    inv01 ix4901 (.Y (nx4902), .A (WindowDin_2__4__6)) ;
    mux21 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix181 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_8), .A0 (nx4904), .A1 (
          nx4906), .S0 (nx8174)) ;
    inv01 ix4903 (.Y (nx4904), .A (L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_9)) ;
    inv01 ix4905 (.Y (nx4906), .A (WindowDin_2__4__7)) ;
    nor02_2x L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix89 (.Y (
             L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_9), .A0 (nx8174), .A1 (
             nx4908)) ;
    inv01 ix4907 (.Y (nx4908), .A (L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_10)
          ) ;
    nor02_2x L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix93 (.Y (
             L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_10), .A0 (nx8174), .A1 (
             nx4910)) ;
    inv01 ix4909 (.Y (nx4910), .A (L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_11)
          ) ;
    nor02_2x L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix97 (.Y (
             L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_11), .A0 (nx8174), .A1 (
             nx4912)) ;
    inv01 ix4911 (.Y (nx4912), .A (L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_12)
          ) ;
    nor02_2x L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix101 (.Y (
             L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_12), .A0 (nx8174), .A1 (
             nx4914)) ;
    inv01 ix4913 (.Y (nx4914), .A (L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_13)
          ) ;
    nor02_2x L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix105 (.Y (
             L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_13), .A0 (nx8174), .A1 (
             nx4916)) ;
    inv01 ix4915 (.Y (nx4916), .A (L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_14)
          ) ;
    nor02_2x L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix109 (.Y (
             L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_14), .A0 (nx8176), .A1 (
             nx4918)) ;
    inv01 ix4917 (.Y (nx4918), .A (L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_15)
          ) ;
    nor02_2x L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix113 (.Y (
             L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_15), .A0 (nx8176), .A1 (
             nx4920)) ;
    inv01 ix4919 (.Y (nx4920), .A (L1_2_L2_4_G2_MINI_ALU_BoothPBeforeShift_16)
          ) ;
    nor02_2x L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix117 (.Y (
             L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_16), .A0 (nx8176), .A1 (
             nx4920)) ;
    mux21 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix189 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BoothOperand_0), .A0 (nx4922), .A1 (nx4924), .S0 (
          nx8164)) ;
    inv01 ix4921 (.Y (nx4922), .A (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_0)) ;
    inv01 ix4923 (.Y (nx4924), .A (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_0)) ;
    mux21 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix197 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BoothOperand_1), .A0 (nx4926), .A1 (nx4928), .S0 (
          nx8164)) ;
    inv01 ix4925 (.Y (nx4926), .A (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_1)) ;
    inv01 ix4927 (.Y (nx4928), .A (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_1)) ;
    mux21 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix205 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BoothOperand_2), .A0 (nx4930), .A1 (nx4932), .S0 (
          nx8164)) ;
    inv01 ix4929 (.Y (nx4930), .A (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_2)) ;
    inv01 ix4931 (.Y (nx4932), .A (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_2)) ;
    mux21 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix213 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BoothOperand_3), .A0 (nx4934), .A1 (nx4936), .S0 (
          nx8164)) ;
    inv01 ix4933 (.Y (nx4934), .A (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_3)) ;
    inv01 ix4935 (.Y (nx4936), .A (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_3)) ;
    mux21 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix221 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BoothOperand_4), .A0 (nx4938), .A1 (nx4940), .S0 (
          nx8164)) ;
    inv01 ix4937 (.Y (nx4938), .A (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_4)) ;
    inv01 ix4939 (.Y (nx4940), .A (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_4)) ;
    mux21 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix229 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BoothOperand_5), .A0 (nx4942), .A1 (nx4944), .S0 (
          nx8166)) ;
    inv01 ix4941 (.Y (nx4942), .A (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_5)) ;
    inv01 ix4943 (.Y (nx4944), .A (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_5)) ;
    mux21 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix237 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BoothOperand_6), .A0 (nx4946), .A1 (nx4948), .S0 (
          nx8166)) ;
    inv01 ix4945 (.Y (nx4946), .A (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_6)) ;
    inv01 ix4947 (.Y (nx4948), .A (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_6)) ;
    mux21 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix245 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BoothOperand_7), .A0 (nx4950), .A1 (nx4952), .S0 (
          nx8166)) ;
    inv01 ix4949 (.Y (nx4950), .A (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_7)) ;
    inv01 ix4951 (.Y (nx4952), .A (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_7)) ;
    mux21 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix253 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BoothOperand_8), .A0 (nx4954), .A1 (nx4956), .S0 (
          nx8166)) ;
    inv01 ix4953 (.Y (nx4954), .A (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_8)) ;
    inv01 ix4955 (.Y (nx4956), .A (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_8)) ;
    mux21 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix261 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BoothOperand_9), .A0 (nx4958), .A1 (nx4960), .S0 (
          nx8166)) ;
    inv01 ix4957 (.Y (nx4958), .A (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_9)) ;
    inv01 ix4959 (.Y (nx4960), .A (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_9)) ;
    mux21 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix269 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BoothOperand_10), .A0 (nx4962), .A1 (nx4964), .S0 (
          nx8166)) ;
    inv01 ix4961 (.Y (nx4962), .A (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_10)) ;
    inv01 ix4963 (.Y (nx4964), .A (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_10)) ;
    mux21 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix277 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BoothOperand_11), .A0 (nx4966), .A1 (nx4968), .S0 (
          nx8166)) ;
    inv01 ix4965 (.Y (nx4966), .A (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_11)) ;
    inv01 ix4967 (.Y (nx4968), .A (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_11)) ;
    mux21 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix285 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BoothOperand_12), .A0 (nx4970), .A1 (nx4972), .S0 (
          nx8168)) ;
    inv01 ix4969 (.Y (nx4970), .A (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_12)) ;
    inv01 ix4971 (.Y (nx4972), .A (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_12)) ;
    mux21 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix293 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BoothOperand_13), .A0 (nx4974), .A1 (nx4976), .S0 (
          nx8168)) ;
    inv01 ix4973 (.Y (nx4974), .A (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_13)) ;
    inv01 ix4975 (.Y (nx4976), .A (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_13)) ;
    mux21 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix301 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BoothOperand_14), .A0 (nx4978), .A1 (nx4980), .S0 (
          nx8168)) ;
    inv01 ix4977 (.Y (nx4978), .A (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_14)) ;
    inv01 ix4979 (.Y (nx4980), .A (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_14)) ;
    mux21 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix309 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BoothOperand_15), .A0 (nx4982), .A1 (nx4984), .S0 (
          nx8168)) ;
    inv01 ix4981 (.Y (nx4982), .A (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_15)) ;
    inv01 ix4983 (.Y (nx4984), .A (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_15)) ;
    mux21 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix317 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BoothOperand_16), .A0 (nx4986), .A1 (nx4988), .S0 (
          nx8168)) ;
    inv01 ix4985 (.Y (nx4986), .A (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_16)) ;
    inv01 ix4987 (.Y (nx4988), .A (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_16)) ;
    xnor2 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_ix321 (.Y (
          L1_2_L2_4_G2_MINI_ALU_AddPToBoothOperand), .A0 (nx8168), .A1 (nx4854)
          ) ;
    oai32 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix393 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .A0 (nx8680), .A1 (
          RST), .A2 (nx8178), .B0 (nx4924), .B1 (nx4992)) ;
    oai32 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix403 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .A0 (nx8680), .A1 (
          RST), .A2 (nx8178), .B0 (nx4928), .B1 (nx4992)) ;
    oai32 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix413 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .A0 (nx8680), .A1 (
          RST), .A2 (nx8178), .B0 (nx4932), .B1 (nx4992)) ;
    oai32 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix423 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .A0 (nx8680), .A1 (
          RST), .A2 (nx8178), .B0 (nx4936), .B1 (nx4992)) ;
    oai32 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix433 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .A0 (nx8680), .A1 (
          RST), .A2 (nx8178), .B0 (nx4940), .B1 (nx4992)) ;
    oai32 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix443 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .A0 (nx8680), .A1 (
          RST), .A2 (nx8178), .B0 (nx4944), .B1 (nx4992)) ;
    oai32 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix453 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .A0 (nx8680), .A1 (
          RST), .A2 (nx8180), .B0 (nx4948), .B1 (nx4992)) ;
    oai32 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix463 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .A0 (nx8682), .A1 (
          RST), .A2 (nx8180), .B0 (nx4952), .B1 (nx4994)) ;
    oai32 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix473 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .A0 (nx8682), .A1 (
          RST), .A2 (nx8180), .B0 (nx4956), .B1 (nx4994)) ;
    oai32 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix483 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .A0 (nx4996), .A1 (
          RST), .A2 (nx8180), .B0 (nx4960), .B1 (nx4994)) ;
    inv01 ix4995 (.Y (nx4996), .A (FilterDin_2__4__0)) ;
    oai32 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix493 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .A0 (nx4998), .A1 (
          RST), .A2 (nx8180), .B0 (nx4964), .B1 (nx4994)) ;
    inv01 ix4997 (.Y (nx4998), .A (FilterDin_2__4__1)) ;
    oai32 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix503 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .A0 (nx5000), .A1 (
          RST), .A2 (nx8180), .B0 (nx4968), .B1 (nx4994)) ;
    inv01 ix4999 (.Y (nx5000), .A (FilterDin_2__4__2)) ;
    oai32 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix513 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .A0 (nx5002), .A1 (
          RST), .A2 (nx8180), .B0 (nx4972), .B1 (nx4994)) ;
    inv01 ix5001 (.Y (nx5002), .A (FilterDin_2__4__3)) ;
    oai32 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix523 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .A0 (nx5004), .A1 (
          RST), .A2 (nx8182), .B0 (nx4976), .B1 (nx4994)) ;
    inv01 ix5003 (.Y (nx5004), .A (FilterDin_2__4__4)) ;
    oai32 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix533 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .A0 (nx5006), .A1 (
          RST), .A2 (nx8182), .B0 (nx4980), .B1 (nx5008)) ;
    inv01 ix5005 (.Y (nx5006), .A (FilterDin_2__4__5)) ;
    inv01 ix5007 (.Y (nx5008), .A (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566)) ;
    oai32 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix543 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .A0 (nx5010), .A1 (
          RST), .A2 (nx8182), .B0 (nx4984), .B1 (nx5008)) ;
    inv01 ix5009 (.Y (nx5010), .A (FilterDin_2__4__6)) ;
    oai32 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix553 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .A0 (nx5012), .A1 (
          RST), .A2 (nx8182), .B0 (nx4988), .B1 (nx5008)) ;
    inv01 ix5011 (.Y (nx5012), .A (FilterDin_2__4__7)) ;
    nand02_2x L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix633 (.Y (nx4992), .A0 (
              nx7600), .A1 (nx8182)) ;
    nand02_2x L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix635 (.Y (nx4994), .A0 (
              nx7600), .A1 (nx8182)) ;
    oai32 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix393 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .A0 (nx8682), .A1 (
          RST), .A2 (nx8184), .B0 (nx4922), .B1 (nx5014)) ;
    oai32 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix403 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .A0 (nx8682), .A1 (
          RST), .A2 (nx8184), .B0 (nx4926), .B1 (nx5014)) ;
    oai32 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix413 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .A0 (nx8682), .A1 (
          RST), .A2 (nx8184), .B0 (nx4930), .B1 (nx5014)) ;
    oai32 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix423 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .A0 (nx8682), .A1 (
          RST), .A2 (nx8184), .B0 (nx4934), .B1 (nx5014)) ;
    oai32 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix433 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .A0 (nx8682), .A1 (
          RST), .A2 (nx8184), .B0 (nx4938), .B1 (nx5014)) ;
    oai32 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix443 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .A0 (nx8684), .A1 (
          RST), .A2 (nx8184), .B0 (nx4942), .B1 (nx5014)) ;
    oai32 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix453 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .A0 (nx8684), .A1 (
          RST), .A2 (nx8186), .B0 (nx4946), .B1 (nx5014)) ;
    oai32 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix463 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .A0 (nx8684), .A1 (
          RST), .A2 (nx8186), .B0 (nx4950), .B1 (nx5016)) ;
    oai32 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix473 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .A0 (nx8684), .A1 (
          RST), .A2 (nx8186), .B0 (nx4954), .B1 (nx5016)) ;
    oai32 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix483 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .A0 (nx4996), .A1 (
          RST), .A2 (nx8186), .B0 (nx4958), .B1 (nx5016)) ;
    oai32 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix493 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .A0 (nx5018), .A1 (
          RST), .A2 (nx8186), .B0 (nx4962), .B1 (nx5016)) ;
    inv01 ix5017 (.Y (nx5018), .A (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_10)) ;
    oai32 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix503 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .A0 (nx5020), .A1 (
          RST), .A2 (nx8186), .B0 (nx4966), .B1 (nx5016)) ;
    inv01 ix5019 (.Y (nx5020), .A (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_11)) ;
    oai32 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix513 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .A0 (nx5022), .A1 (
          RST), .A2 (nx8186), .B0 (nx4970), .B1 (nx5016)) ;
    inv01 ix5021 (.Y (nx5022), .A (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_12)) ;
    oai32 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix523 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .A0 (nx5024), .A1 (
          RST), .A2 (nx8188), .B0 (nx4974), .B1 (nx5016)) ;
    inv01 ix5023 (.Y (nx5024), .A (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_13)) ;
    oai32 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix533 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .A0 (nx5026), .A1 (
          RST), .A2 (nx8188), .B0 (nx4978), .B1 (nx5028)) ;
    inv01 ix5025 (.Y (nx5026), .A (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_14)) ;
    inv01 ix5027 (.Y (nx5028), .A (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566)) ;
    oai32 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix543 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .A0 (nx5030), .A1 (
          RST), .A2 (nx8188), .B0 (nx4982), .B1 (nx5028)) ;
    inv01 ix5029 (.Y (nx5030), .A (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_15)) ;
    oai32 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix553 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .A0 (nx5032), .A1 (
          RST), .A2 (nx8188), .B0 (nx4986), .B1 (nx5028)) ;
    inv01 ix5031 (.Y (nx5032), .A (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_16)) ;
    nand02_2x L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix633 (.Y (nx5014), .A0 (
              nx7600), .A1 (nx8188)) ;
    nand02_2x L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix635 (.Y (nx5016), .A0 (
              nx7600), .A1 (nx8188)) ;
    oai32 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix393 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .A0 (nx5034), .A1 (
          RST), .A2 (nx8190), .B0 (L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_nx384), .B1 (
          nx5036)) ;
    inv01 ix5033 (.Y (nx5034), .A (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_0)) ;
    oai32 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix403 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .A0 (nx5038), .A1 (
          RST), .A2 (nx8190), .B0 (nx4854), .B1 (nx5036)) ;
    inv01 ix5037 (.Y (nx5038), .A (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_1)) ;
    oai32 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix413 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .A0 (nx5040), .A1 (
          RST), .A2 (nx8190), .B0 (L1_2_L2_4_G2_MINI_ALU_nx387), .B1 (nx5036)) ;
    inv01 ix5039 (.Y (nx5040), .A (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_2)) ;
    oai32 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix423 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .A0 (nx5042), .A1 (
          RST), .A2 (nx8190), .B0 (L1_2_L2_4_G2_MINI_ALU_nx399), .B1 (nx5036)) ;
    inv01 ix5041 (.Y (nx5042), .A (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_3)) ;
    oai32 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix433 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .A0 (nx5044), .A1 (
          RST), .A2 (nx8190), .B0 (L1_2_L2_4_G2_MINI_ALU_nx409), .B1 (nx5036)) ;
    inv01 ix5043 (.Y (nx5044), .A (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_4)) ;
    oai32 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix443 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .A0 (nx5046), .A1 (
          RST), .A2 (nx8190), .B0 (L1_2_L2_4_G2_MINI_ALU_nx419), .B1 (nx5036)) ;
    inv01 ix5045 (.Y (nx5046), .A (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_5)) ;
    oai32 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix453 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .A0 (nx5048), .A1 (
          RST), .A2 (nx8190), .B0 (L1_2_L2_4_G2_MINI_ALU_nx429), .B1 (nx5036)) ;
    inv01 ix5047 (.Y (nx5048), .A (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_6)) ;
    oai32 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix463 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .A0 (nx5050), .A1 (
          RST), .A2 (nx8192), .B0 (L1_2_L2_4_G2_MINI_ALU_nx439), .B1 (nx5052)) ;
    inv01 ix5049 (.Y (nx5050), .A (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_7)) ;
    oai32 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix473 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .A0 (nx5054), .A1 (
          RST), .A2 (nx8192), .B0 (L1_2_L2_4_G2_MINI_ALU_nx449), .B1 (nx5052)) ;
    inv01 ix5053 (.Y (nx5054), .A (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_8)) ;
    oai32 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix483 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .A0 (nx5056), .A1 (
          RST), .A2 (nx8192), .B0 (L1_2_L2_4_G2_MINI_ALU_nx469), .B1 (nx5052)) ;
    inv01 ix5055 (.Y (nx5056), .A (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_9)) ;
    oai32 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix493 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .A0 (nx5058), .A1 (
          RST), .A2 (nx8192), .B0 (L1_2_L2_4_G2_MINI_ALU_nx477), .B1 (nx5052)) ;
    inv01 ix5057 (.Y (nx5058), .A (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_10)) ;
    oai32 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix503 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .A0 (nx5060), .A1 (
          RST), .A2 (nx8192), .B0 (L1_2_L2_4_G2_MINI_ALU_nx485), .B1 (nx5052)) ;
    inv01 ix5059 (.Y (nx5060), .A (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_11)) ;
    oai32 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix513 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .A0 (nx5062), .A1 (
          RST), .A2 (nx8192), .B0 (L1_2_L2_4_G2_MINI_ALU_nx493), .B1 (nx5052)) ;
    inv01 ix5061 (.Y (nx5062), .A (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_12)) ;
    oai32 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix523 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .A0 (nx5064), .A1 (
          RST), .A2 (nx8192), .B0 (L1_2_L2_4_G2_MINI_ALU_nx501), .B1 (nx5052)) ;
    inv01 ix5063 (.Y (nx5064), .A (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_13)) ;
    oai32 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix533 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .A0 (nx5066), .A1 (
          RST), .A2 (nx8194), .B0 (L1_2_L2_4_G2_MINI_ALU_nx509), .B1 (nx5068)) ;
    inv01 ix5065 (.Y (nx5066), .A (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_14)) ;
    inv01 ix5067 (.Y (nx5068), .A (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566)) ;
    oai32 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix543 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .A0 (nx5070), .A1 (
          RST), .A2 (nx8194), .B0 (L1_2_L2_4_G2_MINI_ALU_nx517), .B1 (nx5068)) ;
    inv01 ix5069 (.Y (nx5070), .A (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_15)) ;
    oai32 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix553 (.Y (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .A0 (nx5072), .A1 (
          RST), .A2 (nx8194), .B0 (nx4870), .B1 (nx5068)) ;
    inv01 ix5071 (.Y (nx5072), .A (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_16)) ;
    nand02_2x L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix633 (.Y (nx5036), .A0 (
              nx7600), .A1 (nx8194)) ;
    nand02_2x L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix635 (.Y (nx5052), .A0 (
              nx7600), .A1 (nx8194)) ;
    mux21 L1_3_L2_0_G2_MINI_ALU_ix404 (.Y (L1_3_L2_0_G2_MINI_ALU_nx403), .A0 (
          nx5074), .A1 (L1_3_L2_0_G2_MINI_ALU_BoothP_2), .S0 (
          L1_3_L2_0_G2_MINI_ALU_nx395)) ;
    inv01 ix5073 (.Y (nx5074), .A (L1_3_L2_0_G2_MINI_ALU_nx391)) ;
    mux21 L1_3_L2_0_G2_MINI_ALU_ix414 (.Y (L1_3_L2_0_G2_MINI_ALU_nx413), .A0 (
          nx5076), .A1 (L1_3_L2_0_G2_MINI_ALU_BoothP_3), .S0 (
          L1_3_L2_0_G2_MINI_ALU_nx405)) ;
    inv01 ix5075 (.Y (nx5076), .A (L1_3_L2_0_G2_MINI_ALU_nx403)) ;
    mux21 L1_3_L2_0_G2_MINI_ALU_ix424 (.Y (L1_3_L2_0_G2_MINI_ALU_nx423), .A0 (
          nx5078), .A1 (L1_3_L2_0_G2_MINI_ALU_BoothP_4), .S0 (
          L1_3_L2_0_G2_MINI_ALU_nx415)) ;
    inv01 ix5077 (.Y (nx5078), .A (L1_3_L2_0_G2_MINI_ALU_nx413)) ;
    mux21 L1_3_L2_0_G2_MINI_ALU_ix434 (.Y (L1_3_L2_0_G2_MINI_ALU_nx433), .A0 (
          nx5080), .A1 (L1_3_L2_0_G2_MINI_ALU_BoothP_5), .S0 (
          L1_3_L2_0_G2_MINI_ALU_nx425)) ;
    inv01 ix5079 (.Y (nx5080), .A (L1_3_L2_0_G2_MINI_ALU_nx423)) ;
    mux21 L1_3_L2_0_G2_MINI_ALU_ix444 (.Y (L1_3_L2_0_G2_MINI_ALU_nx443), .A0 (
          nx5082), .A1 (L1_3_L2_0_G2_MINI_ALU_BoothP_6), .S0 (
          L1_3_L2_0_G2_MINI_ALU_nx435)) ;
    inv01 ix5081 (.Y (nx5082), .A (L1_3_L2_0_G2_MINI_ALU_nx433)) ;
    mux21 L1_3_L2_0_G2_MINI_ALU_ix454 (.Y (L1_3_L2_0_G2_MINI_ALU_nx453), .A0 (
          nx5084), .A1 (L1_3_L2_0_G2_MINI_ALU_BoothP_7), .S0 (
          L1_3_L2_0_G2_MINI_ALU_nx445)) ;
    inv01 ix5083 (.Y (nx5084), .A (L1_3_L2_0_G2_MINI_ALU_nx443)) ;
    mux21 L1_3_L2_0_G2_MINI_ALU_ix462 (.Y (L1_3_L2_0_G2_MINI_ALU_nx461), .A0 (
          nx5086), .A1 (L1_3_L2_0_G2_MINI_ALU_BoothP_8), .S0 (
          L1_3_L2_0_G2_MINI_ALU_nx455)) ;
    inv01 ix5085 (.Y (nx5086), .A (L1_3_L2_0_G2_MINI_ALU_nx453)) ;
    mux21 L1_3_L2_0_G2_MINI_ALU_ix468 (.Y (L1_3_L2_0_G2_MINI_ALU_nx467), .A0 (
          nx5088), .A1 (L1_3_L2_0_G2_MINI_ALU_BoothP_9), .S0 (
          L1_3_L2_0_G2_MINI_ALU_nx463)) ;
    inv01 ix5087 (.Y (nx5088), .A (L1_3_L2_0_G2_MINI_ALU_nx461)) ;
    mux21 L1_3_L2_0_G2_MINI_ALU_ix476 (.Y (L1_3_L2_0_G2_MINI_ALU_nx475), .A0 (
          nx5090), .A1 (L1_3_L2_0_G2_MINI_ALU_BoothP_10), .S0 (
          L1_3_L2_0_G2_MINI_ALU_nx471)) ;
    inv01 ix5089 (.Y (nx5090), .A (L1_3_L2_0_G2_MINI_ALU_nx467)) ;
    mux21 L1_3_L2_0_G2_MINI_ALU_ix484 (.Y (L1_3_L2_0_G2_MINI_ALU_nx483), .A0 (
          nx5092), .A1 (L1_3_L2_0_G2_MINI_ALU_BoothP_11), .S0 (
          L1_3_L2_0_G2_MINI_ALU_nx479)) ;
    inv01 ix5091 (.Y (nx5092), .A (L1_3_L2_0_G2_MINI_ALU_nx475)) ;
    mux21 L1_3_L2_0_G2_MINI_ALU_ix492 (.Y (L1_3_L2_0_G2_MINI_ALU_nx491), .A0 (
          nx5094), .A1 (L1_3_L2_0_G2_MINI_ALU_BoothP_12), .S0 (
          L1_3_L2_0_G2_MINI_ALU_nx487)) ;
    inv01 ix5093 (.Y (nx5094), .A (L1_3_L2_0_G2_MINI_ALU_nx483)) ;
    mux21 L1_3_L2_0_G2_MINI_ALU_ix500 (.Y (L1_3_L2_0_G2_MINI_ALU_nx499), .A0 (
          nx5096), .A1 (L1_3_L2_0_G2_MINI_ALU_BoothP_13), .S0 (
          L1_3_L2_0_G2_MINI_ALU_nx495)) ;
    inv01 ix5095 (.Y (nx5096), .A (L1_3_L2_0_G2_MINI_ALU_nx491)) ;
    mux21 L1_3_L2_0_G2_MINI_ALU_ix508 (.Y (L1_3_L2_0_G2_MINI_ALU_nx507), .A0 (
          nx5098), .A1 (L1_3_L2_0_G2_MINI_ALU_BoothP_14), .S0 (
          L1_3_L2_0_G2_MINI_ALU_nx503)) ;
    inv01 ix5097 (.Y (nx5098), .A (L1_3_L2_0_G2_MINI_ALU_nx499)) ;
    mux21 L1_3_L2_0_G2_MINI_ALU_ix516 (.Y (L1_3_L2_0_G2_MINI_ALU_nx515), .A0 (
          nx5100), .A1 (L1_3_L2_0_G2_MINI_ALU_BoothP_15), .S0 (
          L1_3_L2_0_G2_MINI_ALU_nx511)) ;
    inv01 ix5099 (.Y (nx5100), .A (L1_3_L2_0_G2_MINI_ALU_nx507)) ;
    mux21 L1_3_L2_0_G2_MINI_ALU_ix161 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_1), .A0 (nx5102), .A1 (
          L1_3_L2_0_G2_MINI_ALU_nx379), .S0 (nx8198)) ;
    inv01 ix5101 (.Y (nx5102), .A (L1_3_L2_0_G2_MINI_ALU_BoothP_1)) ;
    mux21 L1_3_L2_0_G2_MINI_ALU_ix181 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_2), .A0 (
          L1_3_L2_0_G2_MINI_ALU_nx387), .A1 (L1_3_L2_0_G2_MINI_ALU_nx389), .S0 (
          nx8198)) ;
    mux21 L1_3_L2_0_G2_MINI_ALU_ix201 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_3), .A0 (
          L1_3_L2_0_G2_MINI_ALU_nx399), .A1 (L1_3_L2_0_G2_MINI_ALU_nx401), .S0 (
          nx8198)) ;
    mux21 L1_3_L2_0_G2_MINI_ALU_ix221 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_4), .A0 (
          L1_3_L2_0_G2_MINI_ALU_nx409), .A1 (L1_3_L2_0_G2_MINI_ALU_nx411), .S0 (
          nx8198)) ;
    mux21 L1_3_L2_0_G2_MINI_ALU_ix241 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_5), .A0 (
          L1_3_L2_0_G2_MINI_ALU_nx419), .A1 (L1_3_L2_0_G2_MINI_ALU_nx421), .S0 (
          nx8198)) ;
    mux21 L1_3_L2_0_G2_MINI_ALU_ix261 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_6), .A0 (
          L1_3_L2_0_G2_MINI_ALU_nx429), .A1 (L1_3_L2_0_G2_MINI_ALU_nx431), .S0 (
          nx8198)) ;
    mux21 L1_3_L2_0_G2_MINI_ALU_ix281 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_7), .A0 (
          L1_3_L2_0_G2_MINI_ALU_nx439), .A1 (L1_3_L2_0_G2_MINI_ALU_nx441), .S0 (
          nx8198)) ;
    mux21 L1_3_L2_0_G2_MINI_ALU_ix301 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_8), .A0 (
          L1_3_L2_0_G2_MINI_ALU_nx449), .A1 (L1_3_L2_0_G2_MINI_ALU_nx451), .S0 (
          nx8200)) ;
    mux21 L1_3_L2_0_G2_MINI_ALU_ix321 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_9), .A0 (
          L1_3_L2_0_G2_MINI_ALU_nx469), .A1 (nx5104), .S0 (nx8200)) ;
    inv01 ix5103 (.Y (nx5104), .A (L1_3_L2_0_G2_MINI_ALU_nx316)) ;
    mux21 L1_3_L2_0_G2_MINI_ALU_ix341 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_10), .A0 (
          L1_3_L2_0_G2_MINI_ALU_nx477), .A1 (nx5106), .S0 (nx8200)) ;
    inv01 ix5105 (.Y (nx5106), .A (L1_3_L2_0_G2_MINI_ALU_nx336)) ;
    mux21 L1_3_L2_0_G2_MINI_ALU_ix361 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_11), .A0 (
          L1_3_L2_0_G2_MINI_ALU_nx485), .A1 (nx5108), .S0 (nx8200)) ;
    inv01 ix5107 (.Y (nx5108), .A (L1_3_L2_0_G2_MINI_ALU_nx356)) ;
    mux21 L1_3_L2_0_G2_MINI_ALU_ix381 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_12), .A0 (
          L1_3_L2_0_G2_MINI_ALU_nx493), .A1 (nx5110), .S0 (nx8200)) ;
    inv01 ix5109 (.Y (nx5110), .A (L1_3_L2_0_G2_MINI_ALU_nx376)) ;
    mux21 L1_3_L2_0_G2_MINI_ALU_ix401 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_13), .A0 (
          L1_3_L2_0_G2_MINI_ALU_nx501), .A1 (nx5112), .S0 (nx8200)) ;
    inv01 ix5111 (.Y (nx5112), .A (L1_3_L2_0_G2_MINI_ALU_nx396)) ;
    mux21 L1_3_L2_0_G2_MINI_ALU_ix421 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_14), .A0 (
          L1_3_L2_0_G2_MINI_ALU_nx509), .A1 (nx5114), .S0 (nx8200)) ;
    inv01 ix5113 (.Y (nx5114), .A (L1_3_L2_0_G2_MINI_ALU_nx416)) ;
    mux21 L1_3_L2_0_G2_MINI_ALU_ix441 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_15), .A0 (
          L1_3_L2_0_G2_MINI_ALU_nx517), .A1 (nx5116), .S0 (nx8202)) ;
    inv01 ix5115 (.Y (nx5116), .A (L1_3_L2_0_G2_MINI_ALU_nx436)) ;
    mux21 L1_3_L2_0_G2_MINI_ALU_ix461 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_16), .A0 (nx5118), .A1 (nx5120
          ), .S0 (nx8202)) ;
    inv01 ix5117 (.Y (nx5118), .A (L1_3_L2_0_G2_MINI_ALU_BoothP_16)) ;
    inv01 ix5119 (.Y (nx5120), .A (L1_3_L2_0_G2_MINI_ALU_nx456)) ;
    nor02_2x L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix319 (.Y (
             L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642), .A0 (Start), .A1 (
             CalculatingBooth_dup_1162)) ;
    nor02_2x L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix85 (.Y (
             L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_0), .A0 (nx8212), .A1 (
             nx5122)) ;
    inv01 ix5121 (.Y (nx5122), .A (L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_1)) ;
    mux21 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix125 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_1), .A0 (nx5124), .A1 (
          nx5126), .S0 (nx8212)) ;
    inv01 ix5123 (.Y (nx5124), .A (L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_2)) ;
    inv01 ix5125 (.Y (nx5126), .A (WindowDin_3__0__0)) ;
    mux21 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix133 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_2), .A0 (nx5128), .A1 (
          nx5130), .S0 (nx8212)) ;
    inv01 ix5127 (.Y (nx5128), .A (L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_3)) ;
    inv01 ix5129 (.Y (nx5130), .A (WindowDin_3__0__1)) ;
    mux21 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix141 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_3), .A0 (nx5132), .A1 (
          nx5134), .S0 (nx8212)) ;
    inv01 ix5131 (.Y (nx5132), .A (L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_4)) ;
    inv01 ix5133 (.Y (nx5134), .A (WindowDin_3__0__2)) ;
    mux21 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix149 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_4), .A0 (nx5136), .A1 (
          nx5138), .S0 (nx8212)) ;
    inv01 ix5135 (.Y (nx5136), .A (L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_5)) ;
    inv01 ix5137 (.Y (nx5138), .A (WindowDin_3__0__3)) ;
    mux21 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix157 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_5), .A0 (nx5140), .A1 (
          nx5142), .S0 (nx8212)) ;
    inv01 ix5139 (.Y (nx5140), .A (L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_6)) ;
    inv01 ix5141 (.Y (nx5142), .A (WindowDin_3__0__4)) ;
    mux21 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix165 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_6), .A0 (nx5144), .A1 (
          nx5146), .S0 (nx8212)) ;
    inv01 ix5143 (.Y (nx5144), .A (L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_7)) ;
    inv01 ix5145 (.Y (nx5146), .A (WindowDin_3__0__5)) ;
    mux21 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix173 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_7), .A0 (nx5148), .A1 (
          nx5150), .S0 (nx8214)) ;
    inv01 ix5147 (.Y (nx5148), .A (L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_8)) ;
    inv01 ix5149 (.Y (nx5150), .A (WindowDin_3__0__6)) ;
    mux21 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix181 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_8), .A0 (nx5152), .A1 (
          nx5154), .S0 (nx8214)) ;
    inv01 ix5151 (.Y (nx5152), .A (L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_9)) ;
    inv01 ix5153 (.Y (nx5154), .A (WindowDin_3__0__7)) ;
    nor02_2x L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix89 (.Y (
             L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_9), .A0 (nx8214), .A1 (
             nx5156)) ;
    inv01 ix5155 (.Y (nx5156), .A (L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_10)
          ) ;
    nor02_2x L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix93 (.Y (
             L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_10), .A0 (nx8214), .A1 (
             nx5158)) ;
    inv01 ix5157 (.Y (nx5158), .A (L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_11)
          ) ;
    nor02_2x L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix97 (.Y (
             L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_11), .A0 (nx8214), .A1 (
             nx5160)) ;
    inv01 ix5159 (.Y (nx5160), .A (L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_12)
          ) ;
    nor02_2x L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix101 (.Y (
             L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_12), .A0 (nx8214), .A1 (
             nx5162)) ;
    inv01 ix5161 (.Y (nx5162), .A (L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_13)
          ) ;
    nor02_2x L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix105 (.Y (
             L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_13), .A0 (nx8214), .A1 (
             nx5164)) ;
    inv01 ix5163 (.Y (nx5164), .A (L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_14)
          ) ;
    nor02_2x L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix109 (.Y (
             L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_14), .A0 (nx8216), .A1 (
             nx5166)) ;
    inv01 ix5165 (.Y (nx5166), .A (L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_15)
          ) ;
    nor02_2x L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix113 (.Y (
             L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_15), .A0 (nx8216), .A1 (
             nx5168)) ;
    inv01 ix5167 (.Y (nx5168), .A (L1_3_L2_0_G2_MINI_ALU_BoothPBeforeShift_16)
          ) ;
    nor02_2x L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix117 (.Y (
             L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_16), .A0 (nx8216), .A1 (
             nx5168)) ;
    mux21 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix189 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BoothOperand_0), .A0 (nx5170), .A1 (nx5172), .S0 (
          nx8204)) ;
    inv01 ix5169 (.Y (nx5170), .A (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_0)) ;
    inv01 ix5171 (.Y (nx5172), .A (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_0)) ;
    mux21 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix197 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BoothOperand_1), .A0 (nx5174), .A1 (nx5176), .S0 (
          nx8204)) ;
    inv01 ix5173 (.Y (nx5174), .A (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_1)) ;
    inv01 ix5175 (.Y (nx5176), .A (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_1)) ;
    mux21 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix205 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BoothOperand_2), .A0 (nx5178), .A1 (nx5180), .S0 (
          nx8204)) ;
    inv01 ix5177 (.Y (nx5178), .A (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_2)) ;
    inv01 ix5179 (.Y (nx5180), .A (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_2)) ;
    mux21 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix213 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BoothOperand_3), .A0 (nx5182), .A1 (nx5184), .S0 (
          nx8204)) ;
    inv01 ix5181 (.Y (nx5182), .A (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_3)) ;
    inv01 ix5183 (.Y (nx5184), .A (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_3)) ;
    mux21 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix221 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BoothOperand_4), .A0 (nx5186), .A1 (nx5188), .S0 (
          nx8204)) ;
    inv01 ix5185 (.Y (nx5186), .A (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_4)) ;
    inv01 ix5187 (.Y (nx5188), .A (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_4)) ;
    mux21 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix229 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BoothOperand_5), .A0 (nx5190), .A1 (nx5192), .S0 (
          nx8206)) ;
    inv01 ix5189 (.Y (nx5190), .A (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_5)) ;
    inv01 ix5191 (.Y (nx5192), .A (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_5)) ;
    mux21 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix237 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BoothOperand_6), .A0 (nx5194), .A1 (nx5196), .S0 (
          nx8206)) ;
    inv01 ix5193 (.Y (nx5194), .A (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_6)) ;
    inv01 ix5195 (.Y (nx5196), .A (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_6)) ;
    mux21 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix245 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BoothOperand_7), .A0 (nx5198), .A1 (nx5200), .S0 (
          nx8206)) ;
    inv01 ix5197 (.Y (nx5198), .A (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_7)) ;
    inv01 ix5199 (.Y (nx5200), .A (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_7)) ;
    mux21 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix253 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BoothOperand_8), .A0 (nx5202), .A1 (nx5204), .S0 (
          nx8206)) ;
    inv01 ix5201 (.Y (nx5202), .A (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_8)) ;
    inv01 ix5203 (.Y (nx5204), .A (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_8)) ;
    mux21 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix261 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BoothOperand_9), .A0 (nx5206), .A1 (nx5208), .S0 (
          nx8206)) ;
    inv01 ix5205 (.Y (nx5206), .A (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_9)) ;
    inv01 ix5207 (.Y (nx5208), .A (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_9)) ;
    mux21 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix269 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BoothOperand_10), .A0 (nx5210), .A1 (nx5212), .S0 (
          nx8206)) ;
    inv01 ix5209 (.Y (nx5210), .A (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_10)) ;
    inv01 ix5211 (.Y (nx5212), .A (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_10)) ;
    mux21 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix277 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BoothOperand_11), .A0 (nx5214), .A1 (nx5216), .S0 (
          nx8206)) ;
    inv01 ix5213 (.Y (nx5214), .A (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_11)) ;
    inv01 ix5215 (.Y (nx5216), .A (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_11)) ;
    mux21 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix285 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BoothOperand_12), .A0 (nx5218), .A1 (nx5220), .S0 (
          nx8208)) ;
    inv01 ix5217 (.Y (nx5218), .A (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_12)) ;
    inv01 ix5219 (.Y (nx5220), .A (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_12)) ;
    mux21 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix293 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BoothOperand_13), .A0 (nx5222), .A1 (nx5224), .S0 (
          nx8208)) ;
    inv01 ix5221 (.Y (nx5222), .A (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_13)) ;
    inv01 ix5223 (.Y (nx5224), .A (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_13)) ;
    mux21 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix301 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BoothOperand_14), .A0 (nx5226), .A1 (nx5228), .S0 (
          nx8208)) ;
    inv01 ix5225 (.Y (nx5226), .A (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_14)) ;
    inv01 ix5227 (.Y (nx5228), .A (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_14)) ;
    mux21 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix309 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BoothOperand_15), .A0 (nx5230), .A1 (nx5232), .S0 (
          nx8208)) ;
    inv01 ix5229 (.Y (nx5230), .A (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_15)) ;
    inv01 ix5231 (.Y (nx5232), .A (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_15)) ;
    mux21 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix317 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BoothOperand_16), .A0 (nx5234), .A1 (nx5236), .S0 (
          nx8208)) ;
    inv01 ix5233 (.Y (nx5234), .A (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_16)) ;
    inv01 ix5235 (.Y (nx5236), .A (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_16)) ;
    xnor2 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_ix321 (.Y (
          L1_3_L2_0_G2_MINI_ALU_AddPToBoothOperand), .A0 (nx8208), .A1 (nx5102)
          ) ;
    oai32 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix393 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .A0 (nx8686), .A1 (
          RST), .A2 (nx8218), .B0 (nx5172), .B1 (nx5240)) ;
    oai32 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix403 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .A0 (nx8686), .A1 (
          RST), .A2 (nx8218), .B0 (nx5176), .B1 (nx5240)) ;
    oai32 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix413 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .A0 (nx8686), .A1 (
          RST), .A2 (nx8218), .B0 (nx5180), .B1 (nx5240)) ;
    oai32 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix423 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .A0 (nx8686), .A1 (
          RST), .A2 (nx8218), .B0 (nx5184), .B1 (nx5240)) ;
    oai32 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix433 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .A0 (nx8686), .A1 (
          RST), .A2 (nx8218), .B0 (nx5188), .B1 (nx5240)) ;
    oai32 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix443 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .A0 (nx8686), .A1 (
          RST), .A2 (nx8218), .B0 (nx5192), .B1 (nx5240)) ;
    oai32 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix453 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .A0 (nx8686), .A1 (
          RST), .A2 (nx8220), .B0 (nx5196), .B1 (nx5240)) ;
    oai32 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix463 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .A0 (nx8688), .A1 (
          RST), .A2 (nx8220), .B0 (nx5200), .B1 (nx5242)) ;
    oai32 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix473 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .A0 (nx8688), .A1 (
          RST), .A2 (nx8220), .B0 (nx5204), .B1 (nx5242)) ;
    oai32 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix483 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .A0 (nx5244), .A1 (
          RST), .A2 (nx8220), .B0 (nx5208), .B1 (nx5242)) ;
    inv01 ix5243 (.Y (nx5244), .A (FilterDin_3__0__0)) ;
    oai32 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix493 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .A0 (nx5246), .A1 (
          RST), .A2 (nx8220), .B0 (nx5212), .B1 (nx5242)) ;
    inv01 ix5245 (.Y (nx5246), .A (FilterDin_3__0__1)) ;
    oai32 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix503 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .A0 (nx5248), .A1 (
          RST), .A2 (nx8220), .B0 (nx5216), .B1 (nx5242)) ;
    inv01 ix5247 (.Y (nx5248), .A (FilterDin_3__0__2)) ;
    oai32 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix513 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .A0 (nx5250), .A1 (
          RST), .A2 (nx8220), .B0 (nx5220), .B1 (nx5242)) ;
    inv01 ix5249 (.Y (nx5250), .A (FilterDin_3__0__3)) ;
    oai32 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix523 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .A0 (nx5252), .A1 (
          RST), .A2 (nx8222), .B0 (nx5224), .B1 (nx5242)) ;
    inv01 ix5251 (.Y (nx5252), .A (FilterDin_3__0__4)) ;
    oai32 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix533 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .A0 (nx5254), .A1 (
          RST), .A2 (nx8222), .B0 (nx5228), .B1 (nx5256)) ;
    inv01 ix5253 (.Y (nx5254), .A (FilterDin_3__0__5)) ;
    inv01 ix5255 (.Y (nx5256), .A (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566)) ;
    oai32 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix543 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .A0 (nx5258), .A1 (
          RST), .A2 (nx8222), .B0 (nx5232), .B1 (nx5256)) ;
    inv01 ix5257 (.Y (nx5258), .A (FilterDin_3__0__6)) ;
    oai32 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix553 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .A0 (nx5260), .A1 (
          RST), .A2 (nx8222), .B0 (nx5236), .B1 (nx5256)) ;
    inv01 ix5259 (.Y (nx5260), .A (FilterDin_3__0__7)) ;
    nand02_2x L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix633 (.Y (nx5240), .A0 (
              nx7600), .A1 (nx8222)) ;
    nand02_2x L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix635 (.Y (nx5242), .A0 (
              nx7602), .A1 (nx8222)) ;
    oai32 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix393 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .A0 (nx8688), .A1 (
          RST), .A2 (nx8224), .B0 (nx5170), .B1 (nx5262)) ;
    oai32 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix403 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .A0 (nx8688), .A1 (
          RST), .A2 (nx8224), .B0 (nx5174), .B1 (nx5262)) ;
    oai32 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix413 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .A0 (nx8688), .A1 (
          RST), .A2 (nx8224), .B0 (nx5178), .B1 (nx5262)) ;
    oai32 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix423 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .A0 (nx8688), .A1 (
          RST), .A2 (nx8224), .B0 (nx5182), .B1 (nx5262)) ;
    oai32 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix433 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .A0 (nx8688), .A1 (
          RST), .A2 (nx8224), .B0 (nx5186), .B1 (nx5262)) ;
    oai32 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix443 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .A0 (nx8690), .A1 (
          RST), .A2 (nx8224), .B0 (nx5190), .B1 (nx5262)) ;
    oai32 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix453 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .A0 (nx8690), .A1 (
          RST), .A2 (nx8226), .B0 (nx5194), .B1 (nx5262)) ;
    oai32 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix463 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .A0 (nx8690), .A1 (
          RST), .A2 (nx8226), .B0 (nx5198), .B1 (nx5264)) ;
    oai32 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix473 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .A0 (nx8690), .A1 (
          RST), .A2 (nx8226), .B0 (nx5202), .B1 (nx5264)) ;
    oai32 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix483 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .A0 (nx5244), .A1 (
          RST), .A2 (nx8226), .B0 (nx5206), .B1 (nx5264)) ;
    oai32 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix493 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .A0 (nx5266), .A1 (
          RST), .A2 (nx8226), .B0 (nx5210), .B1 (nx5264)) ;
    inv01 ix5265 (.Y (nx5266), .A (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_10)) ;
    oai32 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix503 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .A0 (nx5268), .A1 (
          RST), .A2 (nx8226), .B0 (nx5214), .B1 (nx5264)) ;
    inv01 ix5267 (.Y (nx5268), .A (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_11)) ;
    oai32 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix513 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .A0 (nx5270), .A1 (
          RST), .A2 (nx8226), .B0 (nx5218), .B1 (nx5264)) ;
    inv01 ix5269 (.Y (nx5270), .A (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_12)) ;
    oai32 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix523 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .A0 (nx5272), .A1 (
          RST), .A2 (nx8228), .B0 (nx5222), .B1 (nx5264)) ;
    inv01 ix5271 (.Y (nx5272), .A (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_13)) ;
    oai32 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix533 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .A0 (nx5274), .A1 (
          RST), .A2 (nx8228), .B0 (nx5226), .B1 (nx5276)) ;
    inv01 ix5273 (.Y (nx5274), .A (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_14)) ;
    inv01 ix5275 (.Y (nx5276), .A (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566)) ;
    oai32 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix543 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .A0 (nx5278), .A1 (
          RST), .A2 (nx8228), .B0 (nx5230), .B1 (nx5276)) ;
    inv01 ix5277 (.Y (nx5278), .A (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_15)) ;
    oai32 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix553 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .A0 (nx5280), .A1 (
          RST), .A2 (nx8228), .B0 (nx5234), .B1 (nx5276)) ;
    inv01 ix5279 (.Y (nx5280), .A (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_16)) ;
    nand02_2x L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix633 (.Y (nx5262), .A0 (
              nx7602), .A1 (nx8228)) ;
    nand02_2x L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix635 (.Y (nx5264), .A0 (
              nx7602), .A1 (nx8228)) ;
    oai32 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix393 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .A0 (nx5282), .A1 (
          RST), .A2 (nx8230), .B0 (L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_nx384), .B1 (
          nx5284)) ;
    inv01 ix5281 (.Y (nx5282), .A (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_0)) ;
    oai32 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix403 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .A0 (nx5286), .A1 (
          RST), .A2 (nx8230), .B0 (nx5102), .B1 (nx5284)) ;
    inv01 ix5285 (.Y (nx5286), .A (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_1)) ;
    oai32 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix413 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .A0 (nx5288), .A1 (
          RST), .A2 (nx8230), .B0 (L1_3_L2_0_G2_MINI_ALU_nx387), .B1 (nx5284)) ;
    inv01 ix5287 (.Y (nx5288), .A (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_2)) ;
    oai32 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix423 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .A0 (nx5290), .A1 (
          RST), .A2 (nx8230), .B0 (L1_3_L2_0_G2_MINI_ALU_nx399), .B1 (nx5284)) ;
    inv01 ix5289 (.Y (nx5290), .A (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_3)) ;
    oai32 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix433 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .A0 (nx5292), .A1 (
          RST), .A2 (nx8230), .B0 (L1_3_L2_0_G2_MINI_ALU_nx409), .B1 (nx5284)) ;
    inv01 ix5291 (.Y (nx5292), .A (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_4)) ;
    oai32 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix443 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .A0 (nx5294), .A1 (
          RST), .A2 (nx8230), .B0 (L1_3_L2_0_G2_MINI_ALU_nx419), .B1 (nx5284)) ;
    inv01 ix5293 (.Y (nx5294), .A (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_5)) ;
    oai32 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix453 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .A0 (nx5296), .A1 (
          RST), .A2 (nx8230), .B0 (L1_3_L2_0_G2_MINI_ALU_nx429), .B1 (nx5284)) ;
    inv01 ix5295 (.Y (nx5296), .A (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_6)) ;
    oai32 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix463 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .A0 (nx5298), .A1 (
          RST), .A2 (nx8232), .B0 (L1_3_L2_0_G2_MINI_ALU_nx439), .B1 (nx5300)) ;
    inv01 ix5297 (.Y (nx5298), .A (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_7)) ;
    oai32 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix473 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .A0 (nx5302), .A1 (
          RST), .A2 (nx8232), .B0 (L1_3_L2_0_G2_MINI_ALU_nx449), .B1 (nx5300)) ;
    inv01 ix5301 (.Y (nx5302), .A (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_8)) ;
    oai32 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix483 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .A0 (nx5304), .A1 (
          RST), .A2 (nx8232), .B0 (L1_3_L2_0_G2_MINI_ALU_nx469), .B1 (nx5300)) ;
    inv01 ix5303 (.Y (nx5304), .A (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_9)) ;
    oai32 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix493 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .A0 (nx5306), .A1 (
          RST), .A2 (nx8232), .B0 (L1_3_L2_0_G2_MINI_ALU_nx477), .B1 (nx5300)) ;
    inv01 ix5305 (.Y (nx5306), .A (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_10)) ;
    oai32 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix503 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .A0 (nx5308), .A1 (
          RST), .A2 (nx8232), .B0 (L1_3_L2_0_G2_MINI_ALU_nx485), .B1 (nx5300)) ;
    inv01 ix5307 (.Y (nx5308), .A (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_11)) ;
    oai32 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix513 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .A0 (nx5310), .A1 (
          RST), .A2 (nx8232), .B0 (L1_3_L2_0_G2_MINI_ALU_nx493), .B1 (nx5300)) ;
    inv01 ix5309 (.Y (nx5310), .A (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_12)) ;
    oai32 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix523 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .A0 (nx5312), .A1 (
          RST), .A2 (nx8232), .B0 (L1_3_L2_0_G2_MINI_ALU_nx501), .B1 (nx5300)) ;
    inv01 ix5311 (.Y (nx5312), .A (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_13)) ;
    oai32 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix533 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .A0 (nx5314), .A1 (
          RST), .A2 (nx8234), .B0 (L1_3_L2_0_G2_MINI_ALU_nx509), .B1 (nx5316)) ;
    inv01 ix5313 (.Y (nx5314), .A (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_14)) ;
    inv01 ix5315 (.Y (nx5316), .A (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566)) ;
    oai32 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix543 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .A0 (nx5318), .A1 (
          RST), .A2 (nx8234), .B0 (L1_3_L2_0_G2_MINI_ALU_nx517), .B1 (nx5316)) ;
    inv01 ix5317 (.Y (nx5318), .A (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_15)) ;
    oai32 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix553 (.Y (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .A0 (nx5320), .A1 (
          RST), .A2 (nx8234), .B0 (nx5118), .B1 (nx5316)) ;
    inv01 ix5319 (.Y (nx5320), .A (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_16)) ;
    nand02_2x L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix633 (.Y (nx5284), .A0 (
              nx7602), .A1 (nx8234)) ;
    nand02_2x L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix635 (.Y (nx5300), .A0 (
              nx7602), .A1 (nx8234)) ;
    mux21 L1_3_L2_1_G2_MINI_ALU_ix404 (.Y (L1_3_L2_1_G2_MINI_ALU_nx403), .A0 (
          nx5322), .A1 (L1_3_L2_1_G2_MINI_ALU_BoothP_2), .S0 (
          L1_3_L2_1_G2_MINI_ALU_nx395)) ;
    inv01 ix5321 (.Y (nx5322), .A (L1_3_L2_1_G2_MINI_ALU_nx391)) ;
    mux21 L1_3_L2_1_G2_MINI_ALU_ix414 (.Y (L1_3_L2_1_G2_MINI_ALU_nx413), .A0 (
          nx5324), .A1 (L1_3_L2_1_G2_MINI_ALU_BoothP_3), .S0 (
          L1_3_L2_1_G2_MINI_ALU_nx405)) ;
    inv01 ix5323 (.Y (nx5324), .A (L1_3_L2_1_G2_MINI_ALU_nx403)) ;
    mux21 L1_3_L2_1_G2_MINI_ALU_ix424 (.Y (L1_3_L2_1_G2_MINI_ALU_nx423), .A0 (
          nx5326), .A1 (L1_3_L2_1_G2_MINI_ALU_BoothP_4), .S0 (
          L1_3_L2_1_G2_MINI_ALU_nx415)) ;
    inv01 ix5325 (.Y (nx5326), .A (L1_3_L2_1_G2_MINI_ALU_nx413)) ;
    mux21 L1_3_L2_1_G2_MINI_ALU_ix434 (.Y (L1_3_L2_1_G2_MINI_ALU_nx433), .A0 (
          nx5328), .A1 (L1_3_L2_1_G2_MINI_ALU_BoothP_5), .S0 (
          L1_3_L2_1_G2_MINI_ALU_nx425)) ;
    inv01 ix5327 (.Y (nx5328), .A (L1_3_L2_1_G2_MINI_ALU_nx423)) ;
    mux21 L1_3_L2_1_G2_MINI_ALU_ix444 (.Y (L1_3_L2_1_G2_MINI_ALU_nx443), .A0 (
          nx5330), .A1 (L1_3_L2_1_G2_MINI_ALU_BoothP_6), .S0 (
          L1_3_L2_1_G2_MINI_ALU_nx435)) ;
    inv01 ix5329 (.Y (nx5330), .A (L1_3_L2_1_G2_MINI_ALU_nx433)) ;
    mux21 L1_3_L2_1_G2_MINI_ALU_ix454 (.Y (L1_3_L2_1_G2_MINI_ALU_nx453), .A0 (
          nx5332), .A1 (L1_3_L2_1_G2_MINI_ALU_BoothP_7), .S0 (
          L1_3_L2_1_G2_MINI_ALU_nx445)) ;
    inv01 ix5331 (.Y (nx5332), .A (L1_3_L2_1_G2_MINI_ALU_nx443)) ;
    mux21 L1_3_L2_1_G2_MINI_ALU_ix462 (.Y (L1_3_L2_1_G2_MINI_ALU_nx461), .A0 (
          nx5334), .A1 (L1_3_L2_1_G2_MINI_ALU_BoothP_8), .S0 (
          L1_3_L2_1_G2_MINI_ALU_nx455)) ;
    inv01 ix5333 (.Y (nx5334), .A (L1_3_L2_1_G2_MINI_ALU_nx453)) ;
    mux21 L1_3_L2_1_G2_MINI_ALU_ix468 (.Y (L1_3_L2_1_G2_MINI_ALU_nx467), .A0 (
          nx5336), .A1 (L1_3_L2_1_G2_MINI_ALU_BoothP_9), .S0 (
          L1_3_L2_1_G2_MINI_ALU_nx463)) ;
    inv01 ix5335 (.Y (nx5336), .A (L1_3_L2_1_G2_MINI_ALU_nx461)) ;
    mux21 L1_3_L2_1_G2_MINI_ALU_ix476 (.Y (L1_3_L2_1_G2_MINI_ALU_nx475), .A0 (
          nx5338), .A1 (L1_3_L2_1_G2_MINI_ALU_BoothP_10), .S0 (
          L1_3_L2_1_G2_MINI_ALU_nx471)) ;
    inv01 ix5337 (.Y (nx5338), .A (L1_3_L2_1_G2_MINI_ALU_nx467)) ;
    mux21 L1_3_L2_1_G2_MINI_ALU_ix484 (.Y (L1_3_L2_1_G2_MINI_ALU_nx483), .A0 (
          nx5340), .A1 (L1_3_L2_1_G2_MINI_ALU_BoothP_11), .S0 (
          L1_3_L2_1_G2_MINI_ALU_nx479)) ;
    inv01 ix5339 (.Y (nx5340), .A (L1_3_L2_1_G2_MINI_ALU_nx475)) ;
    mux21 L1_3_L2_1_G2_MINI_ALU_ix492 (.Y (L1_3_L2_1_G2_MINI_ALU_nx491), .A0 (
          nx5342), .A1 (L1_3_L2_1_G2_MINI_ALU_BoothP_12), .S0 (
          L1_3_L2_1_G2_MINI_ALU_nx487)) ;
    inv01 ix5341 (.Y (nx5342), .A (L1_3_L2_1_G2_MINI_ALU_nx483)) ;
    mux21 L1_3_L2_1_G2_MINI_ALU_ix500 (.Y (L1_3_L2_1_G2_MINI_ALU_nx499), .A0 (
          nx5344), .A1 (L1_3_L2_1_G2_MINI_ALU_BoothP_13), .S0 (
          L1_3_L2_1_G2_MINI_ALU_nx495)) ;
    inv01 ix5343 (.Y (nx5344), .A (L1_3_L2_1_G2_MINI_ALU_nx491)) ;
    mux21 L1_3_L2_1_G2_MINI_ALU_ix508 (.Y (L1_3_L2_1_G2_MINI_ALU_nx507), .A0 (
          nx5346), .A1 (L1_3_L2_1_G2_MINI_ALU_BoothP_14), .S0 (
          L1_3_L2_1_G2_MINI_ALU_nx503)) ;
    inv01 ix5345 (.Y (nx5346), .A (L1_3_L2_1_G2_MINI_ALU_nx499)) ;
    mux21 L1_3_L2_1_G2_MINI_ALU_ix516 (.Y (L1_3_L2_1_G2_MINI_ALU_nx515), .A0 (
          nx5348), .A1 (L1_3_L2_1_G2_MINI_ALU_BoothP_15), .S0 (
          L1_3_L2_1_G2_MINI_ALU_nx511)) ;
    inv01 ix5347 (.Y (nx5348), .A (L1_3_L2_1_G2_MINI_ALU_nx507)) ;
    mux21 L1_3_L2_1_G2_MINI_ALU_ix161 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_1), .A0 (nx5350), .A1 (
          L1_3_L2_1_G2_MINI_ALU_nx379), .S0 (nx8238)) ;
    inv01 ix5349 (.Y (nx5350), .A (L1_3_L2_1_G2_MINI_ALU_BoothP_1)) ;
    mux21 L1_3_L2_1_G2_MINI_ALU_ix181 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_2), .A0 (
          L1_3_L2_1_G2_MINI_ALU_nx387), .A1 (L1_3_L2_1_G2_MINI_ALU_nx389), .S0 (
          nx8238)) ;
    mux21 L1_3_L2_1_G2_MINI_ALU_ix201 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_3), .A0 (
          L1_3_L2_1_G2_MINI_ALU_nx399), .A1 (L1_3_L2_1_G2_MINI_ALU_nx401), .S0 (
          nx8238)) ;
    mux21 L1_3_L2_1_G2_MINI_ALU_ix221 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_4), .A0 (
          L1_3_L2_1_G2_MINI_ALU_nx409), .A1 (L1_3_L2_1_G2_MINI_ALU_nx411), .S0 (
          nx8238)) ;
    mux21 L1_3_L2_1_G2_MINI_ALU_ix241 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_5), .A0 (
          L1_3_L2_1_G2_MINI_ALU_nx419), .A1 (L1_3_L2_1_G2_MINI_ALU_nx421), .S0 (
          nx8238)) ;
    mux21 L1_3_L2_1_G2_MINI_ALU_ix261 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_6), .A0 (
          L1_3_L2_1_G2_MINI_ALU_nx429), .A1 (L1_3_L2_1_G2_MINI_ALU_nx431), .S0 (
          nx8238)) ;
    mux21 L1_3_L2_1_G2_MINI_ALU_ix281 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_7), .A0 (
          L1_3_L2_1_G2_MINI_ALU_nx439), .A1 (L1_3_L2_1_G2_MINI_ALU_nx441), .S0 (
          nx8238)) ;
    mux21 L1_3_L2_1_G2_MINI_ALU_ix301 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_8), .A0 (
          L1_3_L2_1_G2_MINI_ALU_nx449), .A1 (L1_3_L2_1_G2_MINI_ALU_nx451), .S0 (
          nx8240)) ;
    mux21 L1_3_L2_1_G2_MINI_ALU_ix321 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_9), .A0 (
          L1_3_L2_1_G2_MINI_ALU_nx469), .A1 (nx5352), .S0 (nx8240)) ;
    inv01 ix5351 (.Y (nx5352), .A (L1_3_L2_1_G2_MINI_ALU_nx316)) ;
    mux21 L1_3_L2_1_G2_MINI_ALU_ix341 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_10), .A0 (
          L1_3_L2_1_G2_MINI_ALU_nx477), .A1 (nx5354), .S0 (nx8240)) ;
    inv01 ix5353 (.Y (nx5354), .A (L1_3_L2_1_G2_MINI_ALU_nx336)) ;
    mux21 L1_3_L2_1_G2_MINI_ALU_ix361 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_11), .A0 (
          L1_3_L2_1_G2_MINI_ALU_nx485), .A1 (nx5356), .S0 (nx8240)) ;
    inv01 ix5355 (.Y (nx5356), .A (L1_3_L2_1_G2_MINI_ALU_nx356)) ;
    mux21 L1_3_L2_1_G2_MINI_ALU_ix381 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_12), .A0 (
          L1_3_L2_1_G2_MINI_ALU_nx493), .A1 (nx5358), .S0 (nx8240)) ;
    inv01 ix5357 (.Y (nx5358), .A (L1_3_L2_1_G2_MINI_ALU_nx376)) ;
    mux21 L1_3_L2_1_G2_MINI_ALU_ix401 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_13), .A0 (
          L1_3_L2_1_G2_MINI_ALU_nx501), .A1 (nx5360), .S0 (nx8240)) ;
    inv01 ix5359 (.Y (nx5360), .A (L1_3_L2_1_G2_MINI_ALU_nx396)) ;
    mux21 L1_3_L2_1_G2_MINI_ALU_ix421 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_14), .A0 (
          L1_3_L2_1_G2_MINI_ALU_nx509), .A1 (nx5362), .S0 (nx8240)) ;
    inv01 ix5361 (.Y (nx5362), .A (L1_3_L2_1_G2_MINI_ALU_nx416)) ;
    mux21 L1_3_L2_1_G2_MINI_ALU_ix441 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_15), .A0 (
          L1_3_L2_1_G2_MINI_ALU_nx517), .A1 (nx5364), .S0 (nx8242)) ;
    inv01 ix5363 (.Y (nx5364), .A (L1_3_L2_1_G2_MINI_ALU_nx436)) ;
    mux21 L1_3_L2_1_G2_MINI_ALU_ix461 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_16), .A0 (nx5366), .A1 (nx5368
          ), .S0 (nx8242)) ;
    inv01 ix5365 (.Y (nx5366), .A (L1_3_L2_1_G2_MINI_ALU_BoothP_16)) ;
    inv01 ix5367 (.Y (nx5368), .A (L1_3_L2_1_G2_MINI_ALU_nx456)) ;
    nor02_2x L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix319 (.Y (
             L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642), .A0 (Start), .A1 (
             CalculatingBooth_dup_1162)) ;
    nor02_2x L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix85 (.Y (
             L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_0), .A0 (nx8252), .A1 (
             nx5370)) ;
    inv01 ix5369 (.Y (nx5370), .A (L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_1)) ;
    mux21 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix125 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_1), .A0 (nx5372), .A1 (
          nx5374), .S0 (nx8252)) ;
    inv01 ix5371 (.Y (nx5372), .A (L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_2)) ;
    inv01 ix5373 (.Y (nx5374), .A (WindowDin_3__1__0)) ;
    mux21 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix133 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_2), .A0 (nx5376), .A1 (
          nx5378), .S0 (nx8252)) ;
    inv01 ix5375 (.Y (nx5376), .A (L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_3)) ;
    inv01 ix5377 (.Y (nx5378), .A (WindowDin_3__1__1)) ;
    mux21 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix141 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_3), .A0 (nx5380), .A1 (
          nx5382), .S0 (nx8252)) ;
    inv01 ix5379 (.Y (nx5380), .A (L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_4)) ;
    inv01 ix5381 (.Y (nx5382), .A (WindowDin_3__1__2)) ;
    mux21 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix149 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_4), .A0 (nx5384), .A1 (
          nx5386), .S0 (nx8252)) ;
    inv01 ix5383 (.Y (nx5384), .A (L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_5)) ;
    inv01 ix5385 (.Y (nx5386), .A (WindowDin_3__1__3)) ;
    mux21 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix157 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_5), .A0 (nx5388), .A1 (
          nx5390), .S0 (nx8252)) ;
    inv01 ix5387 (.Y (nx5388), .A (L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_6)) ;
    inv01 ix5389 (.Y (nx5390), .A (WindowDin_3__1__4)) ;
    mux21 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix165 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_6), .A0 (nx5392), .A1 (
          nx5394), .S0 (nx8252)) ;
    inv01 ix5391 (.Y (nx5392), .A (L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_7)) ;
    inv01 ix5393 (.Y (nx5394), .A (WindowDin_3__1__5)) ;
    mux21 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix173 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_7), .A0 (nx5396), .A1 (
          nx5398), .S0 (nx8254)) ;
    inv01 ix5395 (.Y (nx5396), .A (L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_8)) ;
    inv01 ix5397 (.Y (nx5398), .A (WindowDin_3__1__6)) ;
    mux21 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix181 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_8), .A0 (nx5400), .A1 (
          nx5402), .S0 (nx8254)) ;
    inv01 ix5399 (.Y (nx5400), .A (L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_9)) ;
    inv01 ix5401 (.Y (nx5402), .A (WindowDin_3__1__7)) ;
    nor02_2x L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix89 (.Y (
             L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_9), .A0 (nx8254), .A1 (
             nx5404)) ;
    inv01 ix5403 (.Y (nx5404), .A (L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_10)
          ) ;
    nor02_2x L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix93 (.Y (
             L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_10), .A0 (nx8254), .A1 (
             nx5406)) ;
    inv01 ix5405 (.Y (nx5406), .A (L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_11)
          ) ;
    nor02_2x L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix97 (.Y (
             L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_11), .A0 (nx8254), .A1 (
             nx5408)) ;
    inv01 ix5407 (.Y (nx5408), .A (L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_12)
          ) ;
    nor02_2x L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix101 (.Y (
             L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_12), .A0 (nx8254), .A1 (
             nx5410)) ;
    inv01 ix5409 (.Y (nx5410), .A (L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_13)
          ) ;
    nor02_2x L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix105 (.Y (
             L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_13), .A0 (nx8254), .A1 (
             nx5412)) ;
    inv01 ix5411 (.Y (nx5412), .A (L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_14)
          ) ;
    nor02_2x L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix109 (.Y (
             L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_14), .A0 (nx8256), .A1 (
             nx5414)) ;
    inv01 ix5413 (.Y (nx5414), .A (L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_15)
          ) ;
    nor02_2x L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix113 (.Y (
             L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_15), .A0 (nx8256), .A1 (
             nx5416)) ;
    inv01 ix5415 (.Y (nx5416), .A (L1_3_L2_1_G2_MINI_ALU_BoothPBeforeShift_16)
          ) ;
    nor02_2x L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix117 (.Y (
             L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_16), .A0 (nx8256), .A1 (
             nx5416)) ;
    mux21 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix189 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BoothOperand_0), .A0 (nx5418), .A1 (nx5420), .S0 (
          nx8244)) ;
    inv01 ix5417 (.Y (nx5418), .A (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_0)) ;
    inv01 ix5419 (.Y (nx5420), .A (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_0)) ;
    mux21 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix197 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BoothOperand_1), .A0 (nx5422), .A1 (nx5424), .S0 (
          nx8244)) ;
    inv01 ix5421 (.Y (nx5422), .A (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_1)) ;
    inv01 ix5423 (.Y (nx5424), .A (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_1)) ;
    mux21 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix205 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BoothOperand_2), .A0 (nx5426), .A1 (nx5428), .S0 (
          nx8244)) ;
    inv01 ix5425 (.Y (nx5426), .A (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_2)) ;
    inv01 ix5427 (.Y (nx5428), .A (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_2)) ;
    mux21 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix213 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BoothOperand_3), .A0 (nx5430), .A1 (nx5432), .S0 (
          nx8244)) ;
    inv01 ix5429 (.Y (nx5430), .A (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_3)) ;
    inv01 ix5431 (.Y (nx5432), .A (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_3)) ;
    mux21 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix221 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BoothOperand_4), .A0 (nx5434), .A1 (nx5436), .S0 (
          nx8244)) ;
    inv01 ix5433 (.Y (nx5434), .A (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_4)) ;
    inv01 ix5435 (.Y (nx5436), .A (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_4)) ;
    mux21 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix229 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BoothOperand_5), .A0 (nx5438), .A1 (nx5440), .S0 (
          nx8246)) ;
    inv01 ix5437 (.Y (nx5438), .A (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_5)) ;
    inv01 ix5439 (.Y (nx5440), .A (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_5)) ;
    mux21 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix237 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BoothOperand_6), .A0 (nx5442), .A1 (nx5444), .S0 (
          nx8246)) ;
    inv01 ix5441 (.Y (nx5442), .A (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_6)) ;
    inv01 ix5443 (.Y (nx5444), .A (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_6)) ;
    mux21 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix245 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BoothOperand_7), .A0 (nx5446), .A1 (nx5448), .S0 (
          nx8246)) ;
    inv01 ix5445 (.Y (nx5446), .A (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_7)) ;
    inv01 ix5447 (.Y (nx5448), .A (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_7)) ;
    mux21 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix253 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BoothOperand_8), .A0 (nx5450), .A1 (nx5452), .S0 (
          nx8246)) ;
    inv01 ix5449 (.Y (nx5450), .A (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_8)) ;
    inv01 ix5451 (.Y (nx5452), .A (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_8)) ;
    mux21 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix261 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BoothOperand_9), .A0 (nx5454), .A1 (nx5456), .S0 (
          nx8246)) ;
    inv01 ix5453 (.Y (nx5454), .A (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_9)) ;
    inv01 ix5455 (.Y (nx5456), .A (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_9)) ;
    mux21 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix269 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BoothOperand_10), .A0 (nx5458), .A1 (nx5460), .S0 (
          nx8246)) ;
    inv01 ix5457 (.Y (nx5458), .A (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_10)) ;
    inv01 ix5459 (.Y (nx5460), .A (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_10)) ;
    mux21 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix277 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BoothOperand_11), .A0 (nx5462), .A1 (nx5464), .S0 (
          nx8246)) ;
    inv01 ix5461 (.Y (nx5462), .A (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_11)) ;
    inv01 ix5463 (.Y (nx5464), .A (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_11)) ;
    mux21 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix285 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BoothOperand_12), .A0 (nx5466), .A1 (nx5468), .S0 (
          nx8248)) ;
    inv01 ix5465 (.Y (nx5466), .A (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_12)) ;
    inv01 ix5467 (.Y (nx5468), .A (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_12)) ;
    mux21 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix293 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BoothOperand_13), .A0 (nx5470), .A1 (nx5472), .S0 (
          nx8248)) ;
    inv01 ix5469 (.Y (nx5470), .A (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_13)) ;
    inv01 ix5471 (.Y (nx5472), .A (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_13)) ;
    mux21 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix301 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BoothOperand_14), .A0 (nx5474), .A1 (nx5476), .S0 (
          nx8248)) ;
    inv01 ix5473 (.Y (nx5474), .A (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_14)) ;
    inv01 ix5475 (.Y (nx5476), .A (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_14)) ;
    mux21 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix309 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BoothOperand_15), .A0 (nx5478), .A1 (nx5480), .S0 (
          nx8248)) ;
    inv01 ix5477 (.Y (nx5478), .A (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_15)) ;
    inv01 ix5479 (.Y (nx5480), .A (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_15)) ;
    mux21 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix317 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BoothOperand_16), .A0 (nx5482), .A1 (nx5484), .S0 (
          nx8248)) ;
    inv01 ix5481 (.Y (nx5482), .A (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_16)) ;
    inv01 ix5483 (.Y (nx5484), .A (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_16)) ;
    xnor2 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_ix321 (.Y (
          L1_3_L2_1_G2_MINI_ALU_AddPToBoothOperand), .A0 (nx8248), .A1 (nx5350)
          ) ;
    oai32 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix393 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .A0 (nx8692), .A1 (
          RST), .A2 (nx8258), .B0 (nx5420), .B1 (nx5488)) ;
    oai32 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix403 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .A0 (nx8692), .A1 (
          RST), .A2 (nx8258), .B0 (nx5424), .B1 (nx5488)) ;
    oai32 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix413 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .A0 (nx8692), .A1 (
          RST), .A2 (nx8258), .B0 (nx5428), .B1 (nx5488)) ;
    oai32 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix423 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .A0 (nx8692), .A1 (
          RST), .A2 (nx8258), .B0 (nx5432), .B1 (nx5488)) ;
    oai32 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix433 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .A0 (nx8692), .A1 (
          RST), .A2 (nx8258), .B0 (nx5436), .B1 (nx5488)) ;
    oai32 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix443 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .A0 (nx8692), .A1 (
          RST), .A2 (nx8258), .B0 (nx5440), .B1 (nx5488)) ;
    oai32 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix453 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .A0 (nx8692), .A1 (
          RST), .A2 (nx8260), .B0 (nx5444), .B1 (nx5488)) ;
    oai32 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix463 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .A0 (nx8694), .A1 (
          RST), .A2 (nx8260), .B0 (nx5448), .B1 (nx5490)) ;
    oai32 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix473 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .A0 (nx8694), .A1 (
          RST), .A2 (nx8260), .B0 (nx5452), .B1 (nx5490)) ;
    oai32 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix483 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .A0 (nx5492), .A1 (
          RST), .A2 (nx8260), .B0 (nx5456), .B1 (nx5490)) ;
    inv01 ix5491 (.Y (nx5492), .A (FilterDin_3__1__0)) ;
    oai32 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix493 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .A0 (nx5494), .A1 (
          RST), .A2 (nx8260), .B0 (nx5460), .B1 (nx5490)) ;
    inv01 ix5493 (.Y (nx5494), .A (FilterDin_3__1__1)) ;
    oai32 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix503 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .A0 (nx5496), .A1 (
          RST), .A2 (nx8260), .B0 (nx5464), .B1 (nx5490)) ;
    inv01 ix5495 (.Y (nx5496), .A (FilterDin_3__1__2)) ;
    oai32 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix513 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .A0 (nx5498), .A1 (
          RST), .A2 (nx8260), .B0 (nx5468), .B1 (nx5490)) ;
    inv01 ix5497 (.Y (nx5498), .A (FilterDin_3__1__3)) ;
    oai32 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix523 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .A0 (nx5500), .A1 (
          RST), .A2 (nx8262), .B0 (nx5472), .B1 (nx5490)) ;
    inv01 ix5499 (.Y (nx5500), .A (FilterDin_3__1__4)) ;
    oai32 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix533 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .A0 (nx5502), .A1 (
          RST), .A2 (nx8262), .B0 (nx5476), .B1 (nx5504)) ;
    inv01 ix5501 (.Y (nx5502), .A (FilterDin_3__1__5)) ;
    inv01 ix5503 (.Y (nx5504), .A (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566)) ;
    oai32 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix543 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .A0 (nx5506), .A1 (
          RST), .A2 (nx8262), .B0 (nx5480), .B1 (nx5504)) ;
    inv01 ix5505 (.Y (nx5506), .A (FilterDin_3__1__6)) ;
    oai32 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix553 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .A0 (nx5508), .A1 (
          RST), .A2 (nx8262), .B0 (nx5484), .B1 (nx5504)) ;
    inv01 ix5507 (.Y (nx5508), .A (FilterDin_3__1__7)) ;
    nand02_2x L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix633 (.Y (nx5488), .A0 (
              nx7602), .A1 (nx8262)) ;
    nand02_2x L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix635 (.Y (nx5490), .A0 (
              nx7602), .A1 (nx8262)) ;
    oai32 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix393 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .A0 (nx8694), .A1 (
          RST), .A2 (nx8264), .B0 (nx5418), .B1 (nx5510)) ;
    oai32 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix403 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .A0 (nx8694), .A1 (
          RST), .A2 (nx8264), .B0 (nx5422), .B1 (nx5510)) ;
    oai32 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix413 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .A0 (nx8694), .A1 (
          RST), .A2 (nx8264), .B0 (nx5426), .B1 (nx5510)) ;
    oai32 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix423 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .A0 (nx8694), .A1 (
          RST), .A2 (nx8264), .B0 (nx5430), .B1 (nx5510)) ;
    oai32 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix433 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .A0 (nx8694), .A1 (
          RST), .A2 (nx8264), .B0 (nx5434), .B1 (nx5510)) ;
    oai32 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix443 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .A0 (nx8696), .A1 (
          RST), .A2 (nx8264), .B0 (nx5438), .B1 (nx5510)) ;
    oai32 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix453 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .A0 (nx8696), .A1 (
          RST), .A2 (nx8266), .B0 (nx5442), .B1 (nx5510)) ;
    oai32 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix463 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .A0 (nx8696), .A1 (
          RST), .A2 (nx8266), .B0 (nx5446), .B1 (nx5512)) ;
    oai32 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix473 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .A0 (nx8696), .A1 (
          RST), .A2 (nx8266), .B0 (nx5450), .B1 (nx5512)) ;
    oai32 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix483 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .A0 (nx5492), .A1 (
          RST), .A2 (nx8266), .B0 (nx5454), .B1 (nx5512)) ;
    oai32 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix493 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .A0 (nx5514), .A1 (
          RST), .A2 (nx8266), .B0 (nx5458), .B1 (nx5512)) ;
    inv01 ix5513 (.Y (nx5514), .A (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_10)) ;
    oai32 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix503 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .A0 (nx5516), .A1 (
          RST), .A2 (nx8266), .B0 (nx5462), .B1 (nx5512)) ;
    inv01 ix5515 (.Y (nx5516), .A (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_11)) ;
    oai32 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix513 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .A0 (nx5518), .A1 (
          RST), .A2 (nx8266), .B0 (nx5466), .B1 (nx5512)) ;
    inv01 ix5517 (.Y (nx5518), .A (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_12)) ;
    oai32 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix523 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .A0 (nx5520), .A1 (
          RST), .A2 (nx8268), .B0 (nx5470), .B1 (nx5512)) ;
    inv01 ix5519 (.Y (nx5520), .A (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_13)) ;
    oai32 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix533 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .A0 (nx5522), .A1 (
          RST), .A2 (nx8268), .B0 (nx5474), .B1 (nx5524)) ;
    inv01 ix5521 (.Y (nx5522), .A (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_14)) ;
    inv01 ix5523 (.Y (nx5524), .A (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566)) ;
    oai32 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix543 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .A0 (nx5526), .A1 (
          RST), .A2 (nx8268), .B0 (nx5478), .B1 (nx5524)) ;
    inv01 ix5525 (.Y (nx5526), .A (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_15)) ;
    oai32 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix553 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .A0 (nx5528), .A1 (
          RST), .A2 (nx8268), .B0 (nx5482), .B1 (nx5524)) ;
    inv01 ix5527 (.Y (nx5528), .A (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_16)) ;
    nand02_2x L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix633 (.Y (nx5510), .A0 (
              nx7604), .A1 (nx8268)) ;
    nand02_2x L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix635 (.Y (nx5512), .A0 (
              nx7604), .A1 (nx8268)) ;
    oai32 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix393 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .A0 (nx5530), .A1 (
          RST), .A2 (nx8270), .B0 (L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_nx384), .B1 (
          nx5532)) ;
    inv01 ix5529 (.Y (nx5530), .A (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_0)) ;
    oai32 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix403 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .A0 (nx5534), .A1 (
          RST), .A2 (nx8270), .B0 (nx5350), .B1 (nx5532)) ;
    inv01 ix5533 (.Y (nx5534), .A (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_1)) ;
    oai32 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix413 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .A0 (nx5536), .A1 (
          RST), .A2 (nx8270), .B0 (L1_3_L2_1_G2_MINI_ALU_nx387), .B1 (nx5532)) ;
    inv01 ix5535 (.Y (nx5536), .A (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_2)) ;
    oai32 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix423 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .A0 (nx5538), .A1 (
          RST), .A2 (nx8270), .B0 (L1_3_L2_1_G2_MINI_ALU_nx399), .B1 (nx5532)) ;
    inv01 ix5537 (.Y (nx5538), .A (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_3)) ;
    oai32 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix433 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .A0 (nx5540), .A1 (
          RST), .A2 (nx8270), .B0 (L1_3_L2_1_G2_MINI_ALU_nx409), .B1 (nx5532)) ;
    inv01 ix5539 (.Y (nx5540), .A (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_4)) ;
    oai32 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix443 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .A0 (nx5542), .A1 (
          RST), .A2 (nx8270), .B0 (L1_3_L2_1_G2_MINI_ALU_nx419), .B1 (nx5532)) ;
    inv01 ix5541 (.Y (nx5542), .A (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_5)) ;
    oai32 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix453 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .A0 (nx5544), .A1 (
          RST), .A2 (nx8270), .B0 (L1_3_L2_1_G2_MINI_ALU_nx429), .B1 (nx5532)) ;
    inv01 ix5543 (.Y (nx5544), .A (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_6)) ;
    oai32 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix463 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .A0 (nx5546), .A1 (
          RST), .A2 (nx8272), .B0 (L1_3_L2_1_G2_MINI_ALU_nx439), .B1 (nx5548)) ;
    inv01 ix5545 (.Y (nx5546), .A (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_7)) ;
    oai32 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix473 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .A0 (nx5550), .A1 (
          RST), .A2 (nx8272), .B0 (L1_3_L2_1_G2_MINI_ALU_nx449), .B1 (nx5548)) ;
    inv01 ix5549 (.Y (nx5550), .A (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_8)) ;
    oai32 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix483 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .A0 (nx5552), .A1 (
          RST), .A2 (nx8272), .B0 (L1_3_L2_1_G2_MINI_ALU_nx469), .B1 (nx5548)) ;
    inv01 ix5551 (.Y (nx5552), .A (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_9)) ;
    oai32 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix493 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .A0 (nx5554), .A1 (
          RST), .A2 (nx8272), .B0 (L1_3_L2_1_G2_MINI_ALU_nx477), .B1 (nx5548)) ;
    inv01 ix5553 (.Y (nx5554), .A (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_10)) ;
    oai32 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix503 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .A0 (nx5556), .A1 (
          RST), .A2 (nx8272), .B0 (L1_3_L2_1_G2_MINI_ALU_nx485), .B1 (nx5548)) ;
    inv01 ix5555 (.Y (nx5556), .A (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_11)) ;
    oai32 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix513 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .A0 (nx5558), .A1 (
          RST), .A2 (nx8272), .B0 (L1_3_L2_1_G2_MINI_ALU_nx493), .B1 (nx5548)) ;
    inv01 ix5557 (.Y (nx5558), .A (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_12)) ;
    oai32 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix523 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .A0 (nx5560), .A1 (
          RST), .A2 (nx8272), .B0 (L1_3_L2_1_G2_MINI_ALU_nx501), .B1 (nx5548)) ;
    inv01 ix5559 (.Y (nx5560), .A (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_13)) ;
    oai32 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix533 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .A0 (nx5562), .A1 (
          RST), .A2 (nx8274), .B0 (L1_3_L2_1_G2_MINI_ALU_nx509), .B1 (nx5564)) ;
    inv01 ix5561 (.Y (nx5562), .A (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_14)) ;
    inv01 ix5563 (.Y (nx5564), .A (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566)) ;
    oai32 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix543 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .A0 (nx5566), .A1 (
          RST), .A2 (nx8274), .B0 (L1_3_L2_1_G2_MINI_ALU_nx517), .B1 (nx5564)) ;
    inv01 ix5565 (.Y (nx5566), .A (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_15)) ;
    oai32 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix553 (.Y (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .A0 (nx5568), .A1 (
          RST), .A2 (nx8274), .B0 (nx5366), .B1 (nx5564)) ;
    inv01 ix5567 (.Y (nx5568), .A (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_16)) ;
    nand02_2x L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix633 (.Y (nx5532), .A0 (
              nx7604), .A1 (nx8274)) ;
    nand02_2x L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix635 (.Y (nx5548), .A0 (
              nx7604), .A1 (nx8274)) ;
    mux21 L1_3_L2_2_G2_MINI_ALU_ix404 (.Y (L1_3_L2_2_G2_MINI_ALU_nx403), .A0 (
          nx5570), .A1 (L1_3_L2_2_G2_MINI_ALU_BoothP_2), .S0 (
          L1_3_L2_2_G2_MINI_ALU_nx395)) ;
    inv01 ix5569 (.Y (nx5570), .A (L1_3_L2_2_G2_MINI_ALU_nx391)) ;
    mux21 L1_3_L2_2_G2_MINI_ALU_ix414 (.Y (L1_3_L2_2_G2_MINI_ALU_nx413), .A0 (
          nx5572), .A1 (L1_3_L2_2_G2_MINI_ALU_BoothP_3), .S0 (
          L1_3_L2_2_G2_MINI_ALU_nx405)) ;
    inv01 ix5571 (.Y (nx5572), .A (L1_3_L2_2_G2_MINI_ALU_nx403)) ;
    mux21 L1_3_L2_2_G2_MINI_ALU_ix424 (.Y (L1_3_L2_2_G2_MINI_ALU_nx423), .A0 (
          nx5574), .A1 (L1_3_L2_2_G2_MINI_ALU_BoothP_4), .S0 (
          L1_3_L2_2_G2_MINI_ALU_nx415)) ;
    inv01 ix5573 (.Y (nx5574), .A (L1_3_L2_2_G2_MINI_ALU_nx413)) ;
    mux21 L1_3_L2_2_G2_MINI_ALU_ix434 (.Y (L1_3_L2_2_G2_MINI_ALU_nx433), .A0 (
          nx5576), .A1 (L1_3_L2_2_G2_MINI_ALU_BoothP_5), .S0 (
          L1_3_L2_2_G2_MINI_ALU_nx425)) ;
    inv01 ix5575 (.Y (nx5576), .A (L1_3_L2_2_G2_MINI_ALU_nx423)) ;
    mux21 L1_3_L2_2_G2_MINI_ALU_ix444 (.Y (L1_3_L2_2_G2_MINI_ALU_nx443), .A0 (
          nx5578), .A1 (L1_3_L2_2_G2_MINI_ALU_BoothP_6), .S0 (
          L1_3_L2_2_G2_MINI_ALU_nx435)) ;
    inv01 ix5577 (.Y (nx5578), .A (L1_3_L2_2_G2_MINI_ALU_nx433)) ;
    mux21 L1_3_L2_2_G2_MINI_ALU_ix454 (.Y (L1_3_L2_2_G2_MINI_ALU_nx453), .A0 (
          nx5580), .A1 (L1_3_L2_2_G2_MINI_ALU_BoothP_7), .S0 (
          L1_3_L2_2_G2_MINI_ALU_nx445)) ;
    inv01 ix5579 (.Y (nx5580), .A (L1_3_L2_2_G2_MINI_ALU_nx443)) ;
    mux21 L1_3_L2_2_G2_MINI_ALU_ix462 (.Y (L1_3_L2_2_G2_MINI_ALU_nx461), .A0 (
          nx5582), .A1 (L1_3_L2_2_G2_MINI_ALU_BoothP_8), .S0 (
          L1_3_L2_2_G2_MINI_ALU_nx455)) ;
    inv01 ix5581 (.Y (nx5582), .A (L1_3_L2_2_G2_MINI_ALU_nx453)) ;
    mux21 L1_3_L2_2_G2_MINI_ALU_ix468 (.Y (L1_3_L2_2_G2_MINI_ALU_nx467), .A0 (
          nx5584), .A1 (L1_3_L2_2_G2_MINI_ALU_BoothP_9), .S0 (
          L1_3_L2_2_G2_MINI_ALU_nx463)) ;
    inv01 ix5583 (.Y (nx5584), .A (L1_3_L2_2_G2_MINI_ALU_nx461)) ;
    mux21 L1_3_L2_2_G2_MINI_ALU_ix476 (.Y (L1_3_L2_2_G2_MINI_ALU_nx475), .A0 (
          nx5586), .A1 (L1_3_L2_2_G2_MINI_ALU_BoothP_10), .S0 (
          L1_3_L2_2_G2_MINI_ALU_nx471)) ;
    inv01 ix5585 (.Y (nx5586), .A (L1_3_L2_2_G2_MINI_ALU_nx467)) ;
    mux21 L1_3_L2_2_G2_MINI_ALU_ix484 (.Y (L1_3_L2_2_G2_MINI_ALU_nx483), .A0 (
          nx5588), .A1 (L1_3_L2_2_G2_MINI_ALU_BoothP_11), .S0 (
          L1_3_L2_2_G2_MINI_ALU_nx479)) ;
    inv01 ix5587 (.Y (nx5588), .A (L1_3_L2_2_G2_MINI_ALU_nx475)) ;
    mux21 L1_3_L2_2_G2_MINI_ALU_ix492 (.Y (L1_3_L2_2_G2_MINI_ALU_nx491), .A0 (
          nx5590), .A1 (L1_3_L2_2_G2_MINI_ALU_BoothP_12), .S0 (
          L1_3_L2_2_G2_MINI_ALU_nx487)) ;
    inv01 ix5589 (.Y (nx5590), .A (L1_3_L2_2_G2_MINI_ALU_nx483)) ;
    mux21 L1_3_L2_2_G2_MINI_ALU_ix500 (.Y (L1_3_L2_2_G2_MINI_ALU_nx499), .A0 (
          nx5592), .A1 (L1_3_L2_2_G2_MINI_ALU_BoothP_13), .S0 (
          L1_3_L2_2_G2_MINI_ALU_nx495)) ;
    inv01 ix5591 (.Y (nx5592), .A (L1_3_L2_2_G2_MINI_ALU_nx491)) ;
    mux21 L1_3_L2_2_G2_MINI_ALU_ix508 (.Y (L1_3_L2_2_G2_MINI_ALU_nx507), .A0 (
          nx5594), .A1 (L1_3_L2_2_G2_MINI_ALU_BoothP_14), .S0 (
          L1_3_L2_2_G2_MINI_ALU_nx503)) ;
    inv01 ix5593 (.Y (nx5594), .A (L1_3_L2_2_G2_MINI_ALU_nx499)) ;
    mux21 L1_3_L2_2_G2_MINI_ALU_ix516 (.Y (L1_3_L2_2_G2_MINI_ALU_nx515), .A0 (
          nx5596), .A1 (L1_3_L2_2_G2_MINI_ALU_BoothP_15), .S0 (
          L1_3_L2_2_G2_MINI_ALU_nx511)) ;
    inv01 ix5595 (.Y (nx5596), .A (L1_3_L2_2_G2_MINI_ALU_nx507)) ;
    mux21 L1_3_L2_2_G2_MINI_ALU_ix161 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_1), .A0 (nx5598), .A1 (
          L1_3_L2_2_G2_MINI_ALU_nx379), .S0 (nx8278)) ;
    inv01 ix5597 (.Y (nx5598), .A (L1_3_L2_2_G2_MINI_ALU_BoothP_1)) ;
    mux21 L1_3_L2_2_G2_MINI_ALU_ix181 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_2), .A0 (
          L1_3_L2_2_G2_MINI_ALU_nx387), .A1 (L1_3_L2_2_G2_MINI_ALU_nx389), .S0 (
          nx8278)) ;
    mux21 L1_3_L2_2_G2_MINI_ALU_ix201 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_3), .A0 (
          L1_3_L2_2_G2_MINI_ALU_nx399), .A1 (L1_3_L2_2_G2_MINI_ALU_nx401), .S0 (
          nx8278)) ;
    mux21 L1_3_L2_2_G2_MINI_ALU_ix221 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_4), .A0 (
          L1_3_L2_2_G2_MINI_ALU_nx409), .A1 (L1_3_L2_2_G2_MINI_ALU_nx411), .S0 (
          nx8278)) ;
    mux21 L1_3_L2_2_G2_MINI_ALU_ix241 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_5), .A0 (
          L1_3_L2_2_G2_MINI_ALU_nx419), .A1 (L1_3_L2_2_G2_MINI_ALU_nx421), .S0 (
          nx8278)) ;
    mux21 L1_3_L2_2_G2_MINI_ALU_ix261 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_6), .A0 (
          L1_3_L2_2_G2_MINI_ALU_nx429), .A1 (L1_3_L2_2_G2_MINI_ALU_nx431), .S0 (
          nx8278)) ;
    mux21 L1_3_L2_2_G2_MINI_ALU_ix281 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_7), .A0 (
          L1_3_L2_2_G2_MINI_ALU_nx439), .A1 (L1_3_L2_2_G2_MINI_ALU_nx441), .S0 (
          nx8278)) ;
    mux21 L1_3_L2_2_G2_MINI_ALU_ix301 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_8), .A0 (
          L1_3_L2_2_G2_MINI_ALU_nx449), .A1 (L1_3_L2_2_G2_MINI_ALU_nx451), .S0 (
          nx8280)) ;
    mux21 L1_3_L2_2_G2_MINI_ALU_ix321 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_9), .A0 (
          L1_3_L2_2_G2_MINI_ALU_nx469), .A1 (nx5600), .S0 (nx8280)) ;
    inv01 ix5599 (.Y (nx5600), .A (L1_3_L2_2_G2_MINI_ALU_nx316)) ;
    mux21 L1_3_L2_2_G2_MINI_ALU_ix341 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_10), .A0 (
          L1_3_L2_2_G2_MINI_ALU_nx477), .A1 (nx5602), .S0 (nx8280)) ;
    inv01 ix5601 (.Y (nx5602), .A (L1_3_L2_2_G2_MINI_ALU_nx336)) ;
    mux21 L1_3_L2_2_G2_MINI_ALU_ix361 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_11), .A0 (
          L1_3_L2_2_G2_MINI_ALU_nx485), .A1 (nx5604), .S0 (nx8280)) ;
    inv01 ix5603 (.Y (nx5604), .A (L1_3_L2_2_G2_MINI_ALU_nx356)) ;
    mux21 L1_3_L2_2_G2_MINI_ALU_ix381 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_12), .A0 (
          L1_3_L2_2_G2_MINI_ALU_nx493), .A1 (nx5606), .S0 (nx8280)) ;
    inv01 ix5605 (.Y (nx5606), .A (L1_3_L2_2_G2_MINI_ALU_nx376)) ;
    mux21 L1_3_L2_2_G2_MINI_ALU_ix401 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_13), .A0 (
          L1_3_L2_2_G2_MINI_ALU_nx501), .A1 (nx5608), .S0 (nx8280)) ;
    inv01 ix5607 (.Y (nx5608), .A (L1_3_L2_2_G2_MINI_ALU_nx396)) ;
    mux21 L1_3_L2_2_G2_MINI_ALU_ix421 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_14), .A0 (
          L1_3_L2_2_G2_MINI_ALU_nx509), .A1 (nx5610), .S0 (nx8280)) ;
    inv01 ix5609 (.Y (nx5610), .A (L1_3_L2_2_G2_MINI_ALU_nx416)) ;
    mux21 L1_3_L2_2_G2_MINI_ALU_ix441 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_15), .A0 (
          L1_3_L2_2_G2_MINI_ALU_nx517), .A1 (nx5612), .S0 (nx8282)) ;
    inv01 ix5611 (.Y (nx5612), .A (L1_3_L2_2_G2_MINI_ALU_nx436)) ;
    mux21 L1_3_L2_2_G2_MINI_ALU_ix461 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_16), .A0 (nx5614), .A1 (nx5616
          ), .S0 (nx8282)) ;
    inv01 ix5613 (.Y (nx5614), .A (L1_3_L2_2_G2_MINI_ALU_BoothP_16)) ;
    inv01 ix5615 (.Y (nx5616), .A (L1_3_L2_2_G2_MINI_ALU_nx456)) ;
    nor02_2x L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix319 (.Y (
             L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642), .A0 (Start), .A1 (
             CalculatingBooth_dup_1162)) ;
    nor02_2x L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix85 (.Y (
             L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_0), .A0 (nx8292), .A1 (
             nx5618)) ;
    inv01 ix5617 (.Y (nx5618), .A (L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_1)) ;
    mux21 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix125 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_1), .A0 (nx5620), .A1 (
          nx5622), .S0 (nx8292)) ;
    inv01 ix5619 (.Y (nx5620), .A (L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_2)) ;
    inv01 ix5621 (.Y (nx5622), .A (WindowDin_3__2__0)) ;
    mux21 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix133 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_2), .A0 (nx5624), .A1 (
          nx5626), .S0 (nx8292)) ;
    inv01 ix5623 (.Y (nx5624), .A (L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_3)) ;
    inv01 ix5625 (.Y (nx5626), .A (WindowDin_3__2__1)) ;
    mux21 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix141 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_3), .A0 (nx5628), .A1 (
          nx5630), .S0 (nx8292)) ;
    inv01 ix5627 (.Y (nx5628), .A (L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_4)) ;
    inv01 ix5629 (.Y (nx5630), .A (WindowDin_3__2__2)) ;
    mux21 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix149 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_4), .A0 (nx5632), .A1 (
          nx5634), .S0 (nx8292)) ;
    inv01 ix5631 (.Y (nx5632), .A (L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_5)) ;
    inv01 ix5633 (.Y (nx5634), .A (WindowDin_3__2__3)) ;
    mux21 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix157 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_5), .A0 (nx5636), .A1 (
          nx5638), .S0 (nx8292)) ;
    inv01 ix5635 (.Y (nx5636), .A (L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_6)) ;
    inv01 ix5637 (.Y (nx5638), .A (WindowDin_3__2__4)) ;
    mux21 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix165 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_6), .A0 (nx5640), .A1 (
          nx5642), .S0 (nx8292)) ;
    inv01 ix5639 (.Y (nx5640), .A (L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_7)) ;
    inv01 ix5641 (.Y (nx5642), .A (WindowDin_3__2__5)) ;
    mux21 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix173 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_7), .A0 (nx5644), .A1 (
          nx5646), .S0 (nx8294)) ;
    inv01 ix5643 (.Y (nx5644), .A (L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_8)) ;
    inv01 ix5645 (.Y (nx5646), .A (WindowDin_3__2__6)) ;
    mux21 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix181 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_8), .A0 (nx5648), .A1 (
          nx5650), .S0 (nx8294)) ;
    inv01 ix5647 (.Y (nx5648), .A (L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_9)) ;
    inv01 ix5649 (.Y (nx5650), .A (WindowDin_3__2__7)) ;
    nor02_2x L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix89 (.Y (
             L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_9), .A0 (nx8294), .A1 (
             nx5652)) ;
    inv01 ix5651 (.Y (nx5652), .A (L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_10)
          ) ;
    nor02_2x L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix93 (.Y (
             L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_10), .A0 (nx8294), .A1 (
             nx5654)) ;
    inv01 ix5653 (.Y (nx5654), .A (L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_11)
          ) ;
    nor02_2x L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix97 (.Y (
             L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_11), .A0 (nx8294), .A1 (
             nx5656)) ;
    inv01 ix5655 (.Y (nx5656), .A (L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_12)
          ) ;
    nor02_2x L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix101 (.Y (
             L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_12), .A0 (nx8294), .A1 (
             nx5658)) ;
    inv01 ix5657 (.Y (nx5658), .A (L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_13)
          ) ;
    nor02_2x L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix105 (.Y (
             L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_13), .A0 (nx8294), .A1 (
             nx5660)) ;
    inv01 ix5659 (.Y (nx5660), .A (L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_14)
          ) ;
    nor02_2x L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix109 (.Y (
             L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_14), .A0 (nx8296), .A1 (
             nx5662)) ;
    inv01 ix5661 (.Y (nx5662), .A (L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_15)
          ) ;
    nor02_2x L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix113 (.Y (
             L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_15), .A0 (nx8296), .A1 (
             nx5664)) ;
    inv01 ix5663 (.Y (nx5664), .A (L1_3_L2_2_G2_MINI_ALU_BoothPBeforeShift_16)
          ) ;
    nor02_2x L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix117 (.Y (
             L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_16), .A0 (nx8296), .A1 (
             nx5664)) ;
    mux21 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix189 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BoothOperand_0), .A0 (nx5666), .A1 (nx5668), .S0 (
          nx8284)) ;
    inv01 ix5665 (.Y (nx5666), .A (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_0)) ;
    inv01 ix5667 (.Y (nx5668), .A (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_0)) ;
    mux21 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix197 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BoothOperand_1), .A0 (nx5670), .A1 (nx5672), .S0 (
          nx8284)) ;
    inv01 ix5669 (.Y (nx5670), .A (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_1)) ;
    inv01 ix5671 (.Y (nx5672), .A (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_1)) ;
    mux21 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix205 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BoothOperand_2), .A0 (nx5674), .A1 (nx5676), .S0 (
          nx8284)) ;
    inv01 ix5673 (.Y (nx5674), .A (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_2)) ;
    inv01 ix5675 (.Y (nx5676), .A (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_2)) ;
    mux21 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix213 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BoothOperand_3), .A0 (nx5678), .A1 (nx5680), .S0 (
          nx8284)) ;
    inv01 ix5677 (.Y (nx5678), .A (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_3)) ;
    inv01 ix5679 (.Y (nx5680), .A (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_3)) ;
    mux21 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix221 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BoothOperand_4), .A0 (nx5682), .A1 (nx5684), .S0 (
          nx8284)) ;
    inv01 ix5681 (.Y (nx5682), .A (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_4)) ;
    inv01 ix5683 (.Y (nx5684), .A (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_4)) ;
    mux21 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix229 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BoothOperand_5), .A0 (nx5686), .A1 (nx5688), .S0 (
          nx8286)) ;
    inv01 ix5685 (.Y (nx5686), .A (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_5)) ;
    inv01 ix5687 (.Y (nx5688), .A (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_5)) ;
    mux21 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix237 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BoothOperand_6), .A0 (nx5690), .A1 (nx5692), .S0 (
          nx8286)) ;
    inv01 ix5689 (.Y (nx5690), .A (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_6)) ;
    inv01 ix5691 (.Y (nx5692), .A (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_6)) ;
    mux21 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix245 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BoothOperand_7), .A0 (nx5694), .A1 (nx5696), .S0 (
          nx8286)) ;
    inv01 ix5693 (.Y (nx5694), .A (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_7)) ;
    inv01 ix5695 (.Y (nx5696), .A (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_7)) ;
    mux21 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix253 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BoothOperand_8), .A0 (nx5698), .A1 (nx5700), .S0 (
          nx8286)) ;
    inv01 ix5697 (.Y (nx5698), .A (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_8)) ;
    inv01 ix5699 (.Y (nx5700), .A (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_8)) ;
    mux21 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix261 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BoothOperand_9), .A0 (nx5702), .A1 (nx5704), .S0 (
          nx8286)) ;
    inv01 ix5701 (.Y (nx5702), .A (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_9)) ;
    inv01 ix5703 (.Y (nx5704), .A (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_9)) ;
    mux21 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix269 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BoothOperand_10), .A0 (nx5706), .A1 (nx5708), .S0 (
          nx8286)) ;
    inv01 ix5705 (.Y (nx5706), .A (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_10)) ;
    inv01 ix5707 (.Y (nx5708), .A (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_10)) ;
    mux21 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix277 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BoothOperand_11), .A0 (nx5710), .A1 (nx5712), .S0 (
          nx8286)) ;
    inv01 ix5709 (.Y (nx5710), .A (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_11)) ;
    inv01 ix5711 (.Y (nx5712), .A (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_11)) ;
    mux21 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix285 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BoothOperand_12), .A0 (nx5714), .A1 (nx5716), .S0 (
          nx8288)) ;
    inv01 ix5713 (.Y (nx5714), .A (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_12)) ;
    inv01 ix5715 (.Y (nx5716), .A (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_12)) ;
    mux21 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix293 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BoothOperand_13), .A0 (nx5718), .A1 (nx5720), .S0 (
          nx8288)) ;
    inv01 ix5717 (.Y (nx5718), .A (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_13)) ;
    inv01 ix5719 (.Y (nx5720), .A (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_13)) ;
    mux21 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix301 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BoothOperand_14), .A0 (nx5722), .A1 (nx5724), .S0 (
          nx8288)) ;
    inv01 ix5721 (.Y (nx5722), .A (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_14)) ;
    inv01 ix5723 (.Y (nx5724), .A (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_14)) ;
    mux21 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix309 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BoothOperand_15), .A0 (nx5726), .A1 (nx5728), .S0 (
          nx8288)) ;
    inv01 ix5725 (.Y (nx5726), .A (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_15)) ;
    inv01 ix5727 (.Y (nx5728), .A (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_15)) ;
    mux21 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix317 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BoothOperand_16), .A0 (nx5730), .A1 (nx5732), .S0 (
          nx8288)) ;
    inv01 ix5729 (.Y (nx5730), .A (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_16)) ;
    inv01 ix5731 (.Y (nx5732), .A (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_16)) ;
    xnor2 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_ix321 (.Y (
          L1_3_L2_2_G2_MINI_ALU_AddPToBoothOperand), .A0 (nx8288), .A1 (nx5598)
          ) ;
    oai32 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix393 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .A0 (nx8698), .A1 (
          RST), .A2 (nx8298), .B0 (nx5668), .B1 (nx5736)) ;
    oai32 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix403 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .A0 (nx8698), .A1 (
          RST), .A2 (nx8298), .B0 (nx5672), .B1 (nx5736)) ;
    oai32 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix413 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .A0 (nx8698), .A1 (
          RST), .A2 (nx8298), .B0 (nx5676), .B1 (nx5736)) ;
    oai32 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix423 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .A0 (nx8698), .A1 (
          RST), .A2 (nx8298), .B0 (nx5680), .B1 (nx5736)) ;
    oai32 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix433 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .A0 (nx8698), .A1 (
          RST), .A2 (nx8298), .B0 (nx5684), .B1 (nx5736)) ;
    oai32 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix443 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .A0 (nx8698), .A1 (
          RST), .A2 (nx8298), .B0 (nx5688), .B1 (nx5736)) ;
    oai32 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix453 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .A0 (nx8698), .A1 (
          RST), .A2 (nx8300), .B0 (nx5692), .B1 (nx5736)) ;
    oai32 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix463 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .A0 (nx8700), .A1 (
          RST), .A2 (nx8300), .B0 (nx5696), .B1 (nx5738)) ;
    oai32 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix473 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .A0 (nx8700), .A1 (
          RST), .A2 (nx8300), .B0 (nx5700), .B1 (nx5738)) ;
    oai32 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix483 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .A0 (nx5740), .A1 (
          RST), .A2 (nx8300), .B0 (nx5704), .B1 (nx5738)) ;
    inv01 ix5739 (.Y (nx5740), .A (FilterDin_3__2__0)) ;
    oai32 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix493 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .A0 (nx5742), .A1 (
          RST), .A2 (nx8300), .B0 (nx5708), .B1 (nx5738)) ;
    inv01 ix5741 (.Y (nx5742), .A (FilterDin_3__2__1)) ;
    oai32 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix503 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .A0 (nx5744), .A1 (
          RST), .A2 (nx8300), .B0 (nx5712), .B1 (nx5738)) ;
    inv01 ix5743 (.Y (nx5744), .A (FilterDin_3__2__2)) ;
    oai32 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix513 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .A0 (nx5746), .A1 (
          RST), .A2 (nx8300), .B0 (nx5716), .B1 (nx5738)) ;
    inv01 ix5745 (.Y (nx5746), .A (FilterDin_3__2__3)) ;
    oai32 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix523 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .A0 (nx5748), .A1 (
          RST), .A2 (nx8302), .B0 (nx5720), .B1 (nx5738)) ;
    inv01 ix5747 (.Y (nx5748), .A (FilterDin_3__2__4)) ;
    oai32 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix533 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .A0 (nx5750), .A1 (
          RST), .A2 (nx8302), .B0 (nx5724), .B1 (nx5752)) ;
    inv01 ix5749 (.Y (nx5750), .A (FilterDin_3__2__5)) ;
    inv01 ix5751 (.Y (nx5752), .A (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566)) ;
    oai32 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix543 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .A0 (nx5754), .A1 (
          RST), .A2 (nx8302), .B0 (nx5728), .B1 (nx5752)) ;
    inv01 ix5753 (.Y (nx5754), .A (FilterDin_3__2__6)) ;
    oai32 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix553 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .A0 (nx5756), .A1 (
          RST), .A2 (nx8302), .B0 (nx5732), .B1 (nx5752)) ;
    inv01 ix5755 (.Y (nx5756), .A (FilterDin_3__2__7)) ;
    nand02_2x L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix633 (.Y (nx5736), .A0 (
              nx7604), .A1 (nx8302)) ;
    nand02_2x L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix635 (.Y (nx5738), .A0 (
              nx7604), .A1 (nx8302)) ;
    oai32 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix393 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .A0 (nx8700), .A1 (
          RST), .A2 (nx8304), .B0 (nx5666), .B1 (nx5758)) ;
    oai32 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix403 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .A0 (nx8700), .A1 (
          RST), .A2 (nx8304), .B0 (nx5670), .B1 (nx5758)) ;
    oai32 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix413 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .A0 (nx8700), .A1 (
          RST), .A2 (nx8304), .B0 (nx5674), .B1 (nx5758)) ;
    oai32 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix423 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .A0 (nx8700), .A1 (
          RST), .A2 (nx8304), .B0 (nx5678), .B1 (nx5758)) ;
    oai32 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix433 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .A0 (nx8700), .A1 (
          RST), .A2 (nx8304), .B0 (nx5682), .B1 (nx5758)) ;
    oai32 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix443 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .A0 (nx8702), .A1 (
          RST), .A2 (nx8304), .B0 (nx5686), .B1 (nx5758)) ;
    oai32 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix453 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .A0 (nx8702), .A1 (
          RST), .A2 (nx8306), .B0 (nx5690), .B1 (nx5758)) ;
    oai32 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix463 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .A0 (nx8702), .A1 (
          RST), .A2 (nx8306), .B0 (nx5694), .B1 (nx5760)) ;
    oai32 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix473 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .A0 (nx8702), .A1 (
          RST), .A2 (nx8306), .B0 (nx5698), .B1 (nx5760)) ;
    oai32 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix483 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .A0 (nx5740), .A1 (
          RST), .A2 (nx8306), .B0 (nx5702), .B1 (nx5760)) ;
    oai32 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix493 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .A0 (nx5762), .A1 (
          RST), .A2 (nx8306), .B0 (nx5706), .B1 (nx5760)) ;
    inv01 ix5761 (.Y (nx5762), .A (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_10)) ;
    oai32 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix503 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .A0 (nx5764), .A1 (
          RST), .A2 (nx8306), .B0 (nx5710), .B1 (nx5760)) ;
    inv01 ix5763 (.Y (nx5764), .A (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_11)) ;
    oai32 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix513 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .A0 (nx5766), .A1 (
          RST), .A2 (nx8306), .B0 (nx5714), .B1 (nx5760)) ;
    inv01 ix5765 (.Y (nx5766), .A (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_12)) ;
    oai32 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix523 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .A0 (nx5768), .A1 (
          RST), .A2 (nx8308), .B0 (nx5718), .B1 (nx5760)) ;
    inv01 ix5767 (.Y (nx5768), .A (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_13)) ;
    oai32 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix533 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .A0 (nx5770), .A1 (
          RST), .A2 (nx8308), .B0 (nx5722), .B1 (nx5772)) ;
    inv01 ix5769 (.Y (nx5770), .A (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_14)) ;
    inv01 ix5771 (.Y (nx5772), .A (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566)) ;
    oai32 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix543 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .A0 (nx5774), .A1 (
          RST), .A2 (nx8308), .B0 (nx5726), .B1 (nx5772)) ;
    inv01 ix5773 (.Y (nx5774), .A (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_15)) ;
    oai32 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix553 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .A0 (nx5776), .A1 (
          RST), .A2 (nx8308), .B0 (nx5730), .B1 (nx5772)) ;
    inv01 ix5775 (.Y (nx5776), .A (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_16)) ;
    nand02_2x L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix633 (.Y (nx5758), .A0 (
              nx7604), .A1 (nx8308)) ;
    nand02_2x L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix635 (.Y (nx5760), .A0 (
              nx7606), .A1 (nx8308)) ;
    oai32 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix393 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .A0 (nx5778), .A1 (
          RST), .A2 (nx8310), .B0 (L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_nx384), .B1 (
          nx5780)) ;
    inv01 ix5777 (.Y (nx5778), .A (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_0)) ;
    oai32 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix403 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .A0 (nx5782), .A1 (
          RST), .A2 (nx8310), .B0 (nx5598), .B1 (nx5780)) ;
    inv01 ix5781 (.Y (nx5782), .A (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_1)) ;
    oai32 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix413 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .A0 (nx5784), .A1 (
          RST), .A2 (nx8310), .B0 (L1_3_L2_2_G2_MINI_ALU_nx387), .B1 (nx5780)) ;
    inv01 ix5783 (.Y (nx5784), .A (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_2)) ;
    oai32 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix423 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .A0 (nx5786), .A1 (
          RST), .A2 (nx8310), .B0 (L1_3_L2_2_G2_MINI_ALU_nx399), .B1 (nx5780)) ;
    inv01 ix5785 (.Y (nx5786), .A (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_3)) ;
    oai32 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix433 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .A0 (nx5788), .A1 (
          RST), .A2 (nx8310), .B0 (L1_3_L2_2_G2_MINI_ALU_nx409), .B1 (nx5780)) ;
    inv01 ix5787 (.Y (nx5788), .A (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_4)) ;
    oai32 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix443 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .A0 (nx5790), .A1 (
          RST), .A2 (nx8310), .B0 (L1_3_L2_2_G2_MINI_ALU_nx419), .B1 (nx5780)) ;
    inv01 ix5789 (.Y (nx5790), .A (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_5)) ;
    oai32 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix453 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .A0 (nx5792), .A1 (
          RST), .A2 (nx8310), .B0 (L1_3_L2_2_G2_MINI_ALU_nx429), .B1 (nx5780)) ;
    inv01 ix5791 (.Y (nx5792), .A (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_6)) ;
    oai32 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix463 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .A0 (nx5794), .A1 (
          RST), .A2 (nx8312), .B0 (L1_3_L2_2_G2_MINI_ALU_nx439), .B1 (nx5796)) ;
    inv01 ix5793 (.Y (nx5794), .A (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_7)) ;
    oai32 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix473 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .A0 (nx5798), .A1 (
          RST), .A2 (nx8312), .B0 (L1_3_L2_2_G2_MINI_ALU_nx449), .B1 (nx5796)) ;
    inv01 ix5797 (.Y (nx5798), .A (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_8)) ;
    oai32 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix483 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .A0 (nx5800), .A1 (
          RST), .A2 (nx8312), .B0 (L1_3_L2_2_G2_MINI_ALU_nx469), .B1 (nx5796)) ;
    inv01 ix5799 (.Y (nx5800), .A (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_9)) ;
    oai32 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix493 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .A0 (nx5802), .A1 (
          RST), .A2 (nx8312), .B0 (L1_3_L2_2_G2_MINI_ALU_nx477), .B1 (nx5796)) ;
    inv01 ix5801 (.Y (nx5802), .A (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_10)) ;
    oai32 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix503 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .A0 (nx5804), .A1 (
          RST), .A2 (nx8312), .B0 (L1_3_L2_2_G2_MINI_ALU_nx485), .B1 (nx5796)) ;
    inv01 ix5803 (.Y (nx5804), .A (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_11)) ;
    oai32 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix513 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .A0 (nx5806), .A1 (
          RST), .A2 (nx8312), .B0 (L1_3_L2_2_G2_MINI_ALU_nx493), .B1 (nx5796)) ;
    inv01 ix5805 (.Y (nx5806), .A (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_12)) ;
    oai32 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix523 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .A0 (nx5808), .A1 (
          RST), .A2 (nx8312), .B0 (L1_3_L2_2_G2_MINI_ALU_nx501), .B1 (nx5796)) ;
    inv01 ix5807 (.Y (nx5808), .A (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_13)) ;
    oai32 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix533 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .A0 (nx5810), .A1 (
          RST), .A2 (nx8314), .B0 (L1_3_L2_2_G2_MINI_ALU_nx509), .B1 (nx5812)) ;
    inv01 ix5809 (.Y (nx5810), .A (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_14)) ;
    inv01 ix5811 (.Y (nx5812), .A (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566)) ;
    oai32 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix543 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .A0 (nx5814), .A1 (
          RST), .A2 (nx8314), .B0 (L1_3_L2_2_G2_MINI_ALU_nx517), .B1 (nx5812)) ;
    inv01 ix5813 (.Y (nx5814), .A (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_15)) ;
    oai32 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix553 (.Y (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .A0 (nx5816), .A1 (
          RST), .A2 (nx8314), .B0 (nx5614), .B1 (nx5812)) ;
    inv01 ix5815 (.Y (nx5816), .A (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_16)) ;
    nand02_2x L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix633 (.Y (nx5780), .A0 (
              nx7606), .A1 (nx8314)) ;
    nand02_2x L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix635 (.Y (nx5796), .A0 (
              nx7606), .A1 (nx8314)) ;
    mux21 L1_3_L2_3_G2_MINI_ALU_ix404 (.Y (L1_3_L2_3_G2_MINI_ALU_nx403), .A0 (
          nx5818), .A1 (L1_3_L2_3_G2_MINI_ALU_BoothP_2), .S0 (
          L1_3_L2_3_G2_MINI_ALU_nx395)) ;
    inv01 ix5817 (.Y (nx5818), .A (L1_3_L2_3_G2_MINI_ALU_nx391)) ;
    mux21 L1_3_L2_3_G2_MINI_ALU_ix414 (.Y (L1_3_L2_3_G2_MINI_ALU_nx413), .A0 (
          nx5820), .A1 (L1_3_L2_3_G2_MINI_ALU_BoothP_3), .S0 (
          L1_3_L2_3_G2_MINI_ALU_nx405)) ;
    inv01 ix5819 (.Y (nx5820), .A (L1_3_L2_3_G2_MINI_ALU_nx403)) ;
    mux21 L1_3_L2_3_G2_MINI_ALU_ix424 (.Y (L1_3_L2_3_G2_MINI_ALU_nx423), .A0 (
          nx5822), .A1 (L1_3_L2_3_G2_MINI_ALU_BoothP_4), .S0 (
          L1_3_L2_3_G2_MINI_ALU_nx415)) ;
    inv01 ix5821 (.Y (nx5822), .A (L1_3_L2_3_G2_MINI_ALU_nx413)) ;
    mux21 L1_3_L2_3_G2_MINI_ALU_ix434 (.Y (L1_3_L2_3_G2_MINI_ALU_nx433), .A0 (
          nx5824), .A1 (L1_3_L2_3_G2_MINI_ALU_BoothP_5), .S0 (
          L1_3_L2_3_G2_MINI_ALU_nx425)) ;
    inv01 ix5823 (.Y (nx5824), .A (L1_3_L2_3_G2_MINI_ALU_nx423)) ;
    mux21 L1_3_L2_3_G2_MINI_ALU_ix444 (.Y (L1_3_L2_3_G2_MINI_ALU_nx443), .A0 (
          nx5826), .A1 (L1_3_L2_3_G2_MINI_ALU_BoothP_6), .S0 (
          L1_3_L2_3_G2_MINI_ALU_nx435)) ;
    inv01 ix5825 (.Y (nx5826), .A (L1_3_L2_3_G2_MINI_ALU_nx433)) ;
    mux21 L1_3_L2_3_G2_MINI_ALU_ix454 (.Y (L1_3_L2_3_G2_MINI_ALU_nx453), .A0 (
          nx5828), .A1 (L1_3_L2_3_G2_MINI_ALU_BoothP_7), .S0 (
          L1_3_L2_3_G2_MINI_ALU_nx445)) ;
    inv01 ix5827 (.Y (nx5828), .A (L1_3_L2_3_G2_MINI_ALU_nx443)) ;
    mux21 L1_3_L2_3_G2_MINI_ALU_ix462 (.Y (L1_3_L2_3_G2_MINI_ALU_nx461), .A0 (
          nx5830), .A1 (L1_3_L2_3_G2_MINI_ALU_BoothP_8), .S0 (
          L1_3_L2_3_G2_MINI_ALU_nx455)) ;
    inv01 ix5829 (.Y (nx5830), .A (L1_3_L2_3_G2_MINI_ALU_nx453)) ;
    mux21 L1_3_L2_3_G2_MINI_ALU_ix468 (.Y (L1_3_L2_3_G2_MINI_ALU_nx467), .A0 (
          nx5832), .A1 (L1_3_L2_3_G2_MINI_ALU_BoothP_9), .S0 (
          L1_3_L2_3_G2_MINI_ALU_nx463)) ;
    inv01 ix5831 (.Y (nx5832), .A (L1_3_L2_3_G2_MINI_ALU_nx461)) ;
    mux21 L1_3_L2_3_G2_MINI_ALU_ix476 (.Y (L1_3_L2_3_G2_MINI_ALU_nx475), .A0 (
          nx5834), .A1 (L1_3_L2_3_G2_MINI_ALU_BoothP_10), .S0 (
          L1_3_L2_3_G2_MINI_ALU_nx471)) ;
    inv01 ix5833 (.Y (nx5834), .A (L1_3_L2_3_G2_MINI_ALU_nx467)) ;
    mux21 L1_3_L2_3_G2_MINI_ALU_ix484 (.Y (L1_3_L2_3_G2_MINI_ALU_nx483), .A0 (
          nx5836), .A1 (L1_3_L2_3_G2_MINI_ALU_BoothP_11), .S0 (
          L1_3_L2_3_G2_MINI_ALU_nx479)) ;
    inv01 ix5835 (.Y (nx5836), .A (L1_3_L2_3_G2_MINI_ALU_nx475)) ;
    mux21 L1_3_L2_3_G2_MINI_ALU_ix492 (.Y (L1_3_L2_3_G2_MINI_ALU_nx491), .A0 (
          nx5838), .A1 (L1_3_L2_3_G2_MINI_ALU_BoothP_12), .S0 (
          L1_3_L2_3_G2_MINI_ALU_nx487)) ;
    inv01 ix5837 (.Y (nx5838), .A (L1_3_L2_3_G2_MINI_ALU_nx483)) ;
    mux21 L1_3_L2_3_G2_MINI_ALU_ix500 (.Y (L1_3_L2_3_G2_MINI_ALU_nx499), .A0 (
          nx5840), .A1 (L1_3_L2_3_G2_MINI_ALU_BoothP_13), .S0 (
          L1_3_L2_3_G2_MINI_ALU_nx495)) ;
    inv01 ix5839 (.Y (nx5840), .A (L1_3_L2_3_G2_MINI_ALU_nx491)) ;
    mux21 L1_3_L2_3_G2_MINI_ALU_ix508 (.Y (L1_3_L2_3_G2_MINI_ALU_nx507), .A0 (
          nx5842), .A1 (L1_3_L2_3_G2_MINI_ALU_BoothP_14), .S0 (
          L1_3_L2_3_G2_MINI_ALU_nx503)) ;
    inv01 ix5841 (.Y (nx5842), .A (L1_3_L2_3_G2_MINI_ALU_nx499)) ;
    mux21 L1_3_L2_3_G2_MINI_ALU_ix516 (.Y (L1_3_L2_3_G2_MINI_ALU_nx515), .A0 (
          nx5844), .A1 (L1_3_L2_3_G2_MINI_ALU_BoothP_15), .S0 (
          L1_3_L2_3_G2_MINI_ALU_nx511)) ;
    inv01 ix5843 (.Y (nx5844), .A (L1_3_L2_3_G2_MINI_ALU_nx507)) ;
    mux21 L1_3_L2_3_G2_MINI_ALU_ix161 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_1), .A0 (nx5846), .A1 (
          L1_3_L2_3_G2_MINI_ALU_nx379), .S0 (nx8318)) ;
    inv01 ix5845 (.Y (nx5846), .A (L1_3_L2_3_G2_MINI_ALU_BoothP_1)) ;
    mux21 L1_3_L2_3_G2_MINI_ALU_ix181 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_2), .A0 (
          L1_3_L2_3_G2_MINI_ALU_nx387), .A1 (L1_3_L2_3_G2_MINI_ALU_nx389), .S0 (
          nx8318)) ;
    mux21 L1_3_L2_3_G2_MINI_ALU_ix201 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_3), .A0 (
          L1_3_L2_3_G2_MINI_ALU_nx399), .A1 (L1_3_L2_3_G2_MINI_ALU_nx401), .S0 (
          nx8318)) ;
    mux21 L1_3_L2_3_G2_MINI_ALU_ix221 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_4), .A0 (
          L1_3_L2_3_G2_MINI_ALU_nx409), .A1 (L1_3_L2_3_G2_MINI_ALU_nx411), .S0 (
          nx8318)) ;
    mux21 L1_3_L2_3_G2_MINI_ALU_ix241 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_5), .A0 (
          L1_3_L2_3_G2_MINI_ALU_nx419), .A1 (L1_3_L2_3_G2_MINI_ALU_nx421), .S0 (
          nx8318)) ;
    mux21 L1_3_L2_3_G2_MINI_ALU_ix261 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_6), .A0 (
          L1_3_L2_3_G2_MINI_ALU_nx429), .A1 (L1_3_L2_3_G2_MINI_ALU_nx431), .S0 (
          nx8318)) ;
    mux21 L1_3_L2_3_G2_MINI_ALU_ix281 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_7), .A0 (
          L1_3_L2_3_G2_MINI_ALU_nx439), .A1 (L1_3_L2_3_G2_MINI_ALU_nx441), .S0 (
          nx8318)) ;
    mux21 L1_3_L2_3_G2_MINI_ALU_ix301 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_8), .A0 (
          L1_3_L2_3_G2_MINI_ALU_nx449), .A1 (L1_3_L2_3_G2_MINI_ALU_nx451), .S0 (
          nx8320)) ;
    mux21 L1_3_L2_3_G2_MINI_ALU_ix321 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_9), .A0 (
          L1_3_L2_3_G2_MINI_ALU_nx469), .A1 (nx5848), .S0 (nx8320)) ;
    inv01 ix5847 (.Y (nx5848), .A (L1_3_L2_3_G2_MINI_ALU_nx316)) ;
    mux21 L1_3_L2_3_G2_MINI_ALU_ix341 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_10), .A0 (
          L1_3_L2_3_G2_MINI_ALU_nx477), .A1 (nx5850), .S0 (nx8320)) ;
    inv01 ix5849 (.Y (nx5850), .A (L1_3_L2_3_G2_MINI_ALU_nx336)) ;
    mux21 L1_3_L2_3_G2_MINI_ALU_ix361 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_11), .A0 (
          L1_3_L2_3_G2_MINI_ALU_nx485), .A1 (nx5852), .S0 (nx8320)) ;
    inv01 ix5851 (.Y (nx5852), .A (L1_3_L2_3_G2_MINI_ALU_nx356)) ;
    mux21 L1_3_L2_3_G2_MINI_ALU_ix381 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_12), .A0 (
          L1_3_L2_3_G2_MINI_ALU_nx493), .A1 (nx5854), .S0 (nx8320)) ;
    inv01 ix5853 (.Y (nx5854), .A (L1_3_L2_3_G2_MINI_ALU_nx376)) ;
    mux21 L1_3_L2_3_G2_MINI_ALU_ix401 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_13), .A0 (
          L1_3_L2_3_G2_MINI_ALU_nx501), .A1 (nx5856), .S0 (nx8320)) ;
    inv01 ix5855 (.Y (nx5856), .A (L1_3_L2_3_G2_MINI_ALU_nx396)) ;
    mux21 L1_3_L2_3_G2_MINI_ALU_ix421 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_14), .A0 (
          L1_3_L2_3_G2_MINI_ALU_nx509), .A1 (nx5858), .S0 (nx8320)) ;
    inv01 ix5857 (.Y (nx5858), .A (L1_3_L2_3_G2_MINI_ALU_nx416)) ;
    mux21 L1_3_L2_3_G2_MINI_ALU_ix441 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_15), .A0 (
          L1_3_L2_3_G2_MINI_ALU_nx517), .A1 (nx5860), .S0 (nx8322)) ;
    inv01 ix5859 (.Y (nx5860), .A (L1_3_L2_3_G2_MINI_ALU_nx436)) ;
    mux21 L1_3_L2_3_G2_MINI_ALU_ix461 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_16), .A0 (nx5862), .A1 (nx5864
          ), .S0 (nx8322)) ;
    inv01 ix5861 (.Y (nx5862), .A (L1_3_L2_3_G2_MINI_ALU_BoothP_16)) ;
    inv01 ix5863 (.Y (nx5864), .A (L1_3_L2_3_G2_MINI_ALU_nx456)) ;
    nor02_2x L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix319 (.Y (
             L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642), .A0 (Start), .A1 (
             CalculatingBooth_dup_1162)) ;
    nor02_2x L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix85 (.Y (
             L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_0), .A0 (nx8332), .A1 (
             nx5866)) ;
    inv01 ix5865 (.Y (nx5866), .A (L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_1)) ;
    mux21 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix125 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_1), .A0 (nx5868), .A1 (
          nx5870), .S0 (nx8332)) ;
    inv01 ix5867 (.Y (nx5868), .A (L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_2)) ;
    inv01 ix5869 (.Y (nx5870), .A (WindowDin_3__3__0)) ;
    mux21 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix133 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_2), .A0 (nx5872), .A1 (
          nx5874), .S0 (nx8332)) ;
    inv01 ix5871 (.Y (nx5872), .A (L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_3)) ;
    inv01 ix5873 (.Y (nx5874), .A (WindowDin_3__3__1)) ;
    mux21 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix141 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_3), .A0 (nx5876), .A1 (
          nx5878), .S0 (nx8332)) ;
    inv01 ix5875 (.Y (nx5876), .A (L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_4)) ;
    inv01 ix5877 (.Y (nx5878), .A (WindowDin_3__3__2)) ;
    mux21 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix149 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_4), .A0 (nx5880), .A1 (
          nx5882), .S0 (nx8332)) ;
    inv01 ix5879 (.Y (nx5880), .A (L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_5)) ;
    inv01 ix5881 (.Y (nx5882), .A (WindowDin_3__3__3)) ;
    mux21 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix157 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_5), .A0 (nx5884), .A1 (
          nx5886), .S0 (nx8332)) ;
    inv01 ix5883 (.Y (nx5884), .A (L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_6)) ;
    inv01 ix5885 (.Y (nx5886), .A (WindowDin_3__3__4)) ;
    mux21 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix165 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_6), .A0 (nx5888), .A1 (
          nx5890), .S0 (nx8332)) ;
    inv01 ix5887 (.Y (nx5888), .A (L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_7)) ;
    inv01 ix5889 (.Y (nx5890), .A (WindowDin_3__3__5)) ;
    mux21 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix173 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_7), .A0 (nx5892), .A1 (
          nx5894), .S0 (nx8334)) ;
    inv01 ix5891 (.Y (nx5892), .A (L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_8)) ;
    inv01 ix5893 (.Y (nx5894), .A (WindowDin_3__3__6)) ;
    mux21 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix181 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_8), .A0 (nx5896), .A1 (
          nx5898), .S0 (nx8334)) ;
    inv01 ix5895 (.Y (nx5896), .A (L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_9)) ;
    inv01 ix5897 (.Y (nx5898), .A (WindowDin_3__3__7)) ;
    nor02_2x L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix89 (.Y (
             L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_9), .A0 (nx8334), .A1 (
             nx5900)) ;
    inv01 ix5899 (.Y (nx5900), .A (L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_10)
          ) ;
    nor02_2x L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix93 (.Y (
             L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_10), .A0 (nx8334), .A1 (
             nx5902)) ;
    inv01 ix5901 (.Y (nx5902), .A (L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_11)
          ) ;
    nor02_2x L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix97 (.Y (
             L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_11), .A0 (nx8334), .A1 (
             nx5904)) ;
    inv01 ix5903 (.Y (nx5904), .A (L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_12)
          ) ;
    nor02_2x L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix101 (.Y (
             L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_12), .A0 (nx8334), .A1 (
             nx5906)) ;
    inv01 ix5905 (.Y (nx5906), .A (L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_13)
          ) ;
    nor02_2x L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix105 (.Y (
             L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_13), .A0 (nx8334), .A1 (
             nx5908)) ;
    inv01 ix5907 (.Y (nx5908), .A (L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_14)
          ) ;
    nor02_2x L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix109 (.Y (
             L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_14), .A0 (nx8336), .A1 (
             nx5910)) ;
    inv01 ix5909 (.Y (nx5910), .A (L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_15)
          ) ;
    nor02_2x L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix113 (.Y (
             L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_15), .A0 (nx8336), .A1 (
             nx5912)) ;
    inv01 ix5911 (.Y (nx5912), .A (L1_3_L2_3_G2_MINI_ALU_BoothPBeforeShift_16)
          ) ;
    nor02_2x L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix117 (.Y (
             L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_16), .A0 (nx8336), .A1 (
             nx5912)) ;
    mux21 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix189 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BoothOperand_0), .A0 (nx5914), .A1 (nx5916), .S0 (
          nx8324)) ;
    inv01 ix5913 (.Y (nx5914), .A (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_0)) ;
    inv01 ix5915 (.Y (nx5916), .A (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_0)) ;
    mux21 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix197 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BoothOperand_1), .A0 (nx5918), .A1 (nx5920), .S0 (
          nx8324)) ;
    inv01 ix5917 (.Y (nx5918), .A (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_1)) ;
    inv01 ix5919 (.Y (nx5920), .A (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_1)) ;
    mux21 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix205 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BoothOperand_2), .A0 (nx5922), .A1 (nx5924), .S0 (
          nx8324)) ;
    inv01 ix5921 (.Y (nx5922), .A (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_2)) ;
    inv01 ix5923 (.Y (nx5924), .A (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_2)) ;
    mux21 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix213 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BoothOperand_3), .A0 (nx5926), .A1 (nx5928), .S0 (
          nx8324)) ;
    inv01 ix5925 (.Y (nx5926), .A (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_3)) ;
    inv01 ix5927 (.Y (nx5928), .A (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_3)) ;
    mux21 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix221 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BoothOperand_4), .A0 (nx5930), .A1 (nx5932), .S0 (
          nx8324)) ;
    inv01 ix5929 (.Y (nx5930), .A (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_4)) ;
    inv01 ix5931 (.Y (nx5932), .A (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_4)) ;
    mux21 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix229 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BoothOperand_5), .A0 (nx5934), .A1 (nx5936), .S0 (
          nx8326)) ;
    inv01 ix5933 (.Y (nx5934), .A (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_5)) ;
    inv01 ix5935 (.Y (nx5936), .A (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_5)) ;
    mux21 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix237 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BoothOperand_6), .A0 (nx5938), .A1 (nx5940), .S0 (
          nx8326)) ;
    inv01 ix5937 (.Y (nx5938), .A (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_6)) ;
    inv01 ix5939 (.Y (nx5940), .A (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_6)) ;
    mux21 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix245 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BoothOperand_7), .A0 (nx5942), .A1 (nx5944), .S0 (
          nx8326)) ;
    inv01 ix5941 (.Y (nx5942), .A (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_7)) ;
    inv01 ix5943 (.Y (nx5944), .A (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_7)) ;
    mux21 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix253 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BoothOperand_8), .A0 (nx5946), .A1 (nx5948), .S0 (
          nx8326)) ;
    inv01 ix5945 (.Y (nx5946), .A (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_8)) ;
    inv01 ix5947 (.Y (nx5948), .A (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_8)) ;
    mux21 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix261 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BoothOperand_9), .A0 (nx5950), .A1 (nx5952), .S0 (
          nx8326)) ;
    inv01 ix5949 (.Y (nx5950), .A (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_9)) ;
    inv01 ix5951 (.Y (nx5952), .A (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_9)) ;
    mux21 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix269 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BoothOperand_10), .A0 (nx5954), .A1 (nx5956), .S0 (
          nx8326)) ;
    inv01 ix5953 (.Y (nx5954), .A (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_10)) ;
    inv01 ix5955 (.Y (nx5956), .A (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_10)) ;
    mux21 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix277 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BoothOperand_11), .A0 (nx5958), .A1 (nx5960), .S0 (
          nx8326)) ;
    inv01 ix5957 (.Y (nx5958), .A (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_11)) ;
    inv01 ix5959 (.Y (nx5960), .A (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_11)) ;
    mux21 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix285 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BoothOperand_12), .A0 (nx5962), .A1 (nx5964), .S0 (
          nx8328)) ;
    inv01 ix5961 (.Y (nx5962), .A (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_12)) ;
    inv01 ix5963 (.Y (nx5964), .A (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_12)) ;
    mux21 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix293 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BoothOperand_13), .A0 (nx5966), .A1 (nx5968), .S0 (
          nx8328)) ;
    inv01 ix5965 (.Y (nx5966), .A (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_13)) ;
    inv01 ix5967 (.Y (nx5968), .A (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_13)) ;
    mux21 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix301 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BoothOperand_14), .A0 (nx5970), .A1 (nx5972), .S0 (
          nx8328)) ;
    inv01 ix5969 (.Y (nx5970), .A (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_14)) ;
    inv01 ix5971 (.Y (nx5972), .A (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_14)) ;
    mux21 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix309 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BoothOperand_15), .A0 (nx5974), .A1 (nx5976), .S0 (
          nx8328)) ;
    inv01 ix5973 (.Y (nx5974), .A (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_15)) ;
    inv01 ix5975 (.Y (nx5976), .A (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_15)) ;
    mux21 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix317 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BoothOperand_16), .A0 (nx5978), .A1 (nx5980), .S0 (
          nx8328)) ;
    inv01 ix5977 (.Y (nx5978), .A (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDout_16)) ;
    inv01 ix5979 (.Y (nx5980), .A (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterADout_16)) ;
    xnor2 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_ix321 (.Y (
          L1_3_L2_3_G2_MINI_ALU_AddPToBoothOperand), .A0 (nx8328), .A1 (nx5846)
          ) ;
    oai32 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix393 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .A0 (nx8704), .A1 (
          RST), .A2 (nx8338), .B0 (nx5916), .B1 (nx5984)) ;
    oai32 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix403 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .A0 (nx8704), .A1 (
          RST), .A2 (nx8338), .B0 (nx5920), .B1 (nx5984)) ;
    oai32 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix413 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .A0 (nx8704), .A1 (
          RST), .A2 (nx8338), .B0 (nx5924), .B1 (nx5984)) ;
    oai32 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix423 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .A0 (nx8704), .A1 (
          RST), .A2 (nx8338), .B0 (nx5928), .B1 (nx5984)) ;
    oai32 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix433 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .A0 (nx8704), .A1 (
          RST), .A2 (nx8338), .B0 (nx5932), .B1 (nx5984)) ;
    oai32 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix443 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .A0 (nx8704), .A1 (
          RST), .A2 (nx8338), .B0 (nx5936), .B1 (nx5984)) ;
    oai32 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix453 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .A0 (nx8704), .A1 (
          RST), .A2 (nx8340), .B0 (nx5940), .B1 (nx5984)) ;
    oai32 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix463 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .A0 (nx8706), .A1 (
          RST), .A2 (nx8340), .B0 (nx5944), .B1 (nx5986)) ;
    oai32 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix473 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .A0 (nx8706), .A1 (
          RST), .A2 (nx8340), .B0 (nx5948), .B1 (nx5986)) ;
    oai32 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix483 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .A0 (nx5988), .A1 (
          RST), .A2 (nx8340), .B0 (nx5952), .B1 (nx5986)) ;
    inv01 ix5987 (.Y (nx5988), .A (FilterDin_3__3__0)) ;
    oai32 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix493 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .A0 (nx5990), .A1 (
          RST), .A2 (nx8340), .B0 (nx5956), .B1 (nx5986)) ;
    inv01 ix5989 (.Y (nx5990), .A (FilterDin_3__3__1)) ;
    oai32 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix503 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .A0 (nx5992), .A1 (
          RST), .A2 (nx8340), .B0 (nx5960), .B1 (nx5986)) ;
    inv01 ix5991 (.Y (nx5992), .A (FilterDin_3__3__2)) ;
    oai32 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix513 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .A0 (nx5994), .A1 (
          RST), .A2 (nx8340), .B0 (nx5964), .B1 (nx5986)) ;
    inv01 ix5993 (.Y (nx5994), .A (FilterDin_3__3__3)) ;
    oai32 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix523 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .A0 (nx5996), .A1 (
          RST), .A2 (nx8342), .B0 (nx5968), .B1 (nx5986)) ;
    inv01 ix5995 (.Y (nx5996), .A (FilterDin_3__3__4)) ;
    oai32 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix533 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .A0 (nx5998), .A1 (
          RST), .A2 (nx8342), .B0 (nx5972), .B1 (nx6000)) ;
    inv01 ix5997 (.Y (nx5998), .A (FilterDin_3__3__5)) ;
    inv01 ix5999 (.Y (nx6000), .A (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566)) ;
    oai32 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix543 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .A0 (nx6002), .A1 (
          RST), .A2 (nx8342), .B0 (nx5976), .B1 (nx6000)) ;
    inv01 ix6001 (.Y (nx6002), .A (FilterDin_3__3__6)) ;
    oai32 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix553 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .A0 (nx6004), .A1 (
          RST), .A2 (nx8342), .B0 (nx5980), .B1 (nx6000)) ;
    inv01 ix6003 (.Y (nx6004), .A (FilterDin_3__3__7)) ;
    nand02_2x L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix633 (.Y (nx5984), .A0 (
              nx7606), .A1 (nx8342)) ;
    nand02_2x L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix635 (.Y (nx5986), .A0 (
              nx7606), .A1 (nx8342)) ;
    oai32 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix393 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .A0 (nx8706), .A1 (
          RST), .A2 (nx8344), .B0 (nx5914), .B1 (nx6006)) ;
    oai32 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix403 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .A0 (nx8706), .A1 (
          RST), .A2 (nx8344), .B0 (nx5918), .B1 (nx6006)) ;
    oai32 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix413 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .A0 (nx8706), .A1 (
          RST), .A2 (nx8344), .B0 (nx5922), .B1 (nx6006)) ;
    oai32 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix423 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .A0 (nx8706), .A1 (
          RST), .A2 (nx8344), .B0 (nx5926), .B1 (nx6006)) ;
    oai32 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix433 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .A0 (nx8706), .A1 (
          RST), .A2 (nx8344), .B0 (nx5930), .B1 (nx6006)) ;
    oai32 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix443 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .A0 (nx8708), .A1 (
          RST), .A2 (nx8344), .B0 (nx5934), .B1 (nx6006)) ;
    oai32 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix453 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .A0 (nx8708), .A1 (
          RST), .A2 (nx8346), .B0 (nx5938), .B1 (nx6006)) ;
    oai32 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix463 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .A0 (nx8708), .A1 (
          RST), .A2 (nx8346), .B0 (nx5942), .B1 (nx6008)) ;
    oai32 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix473 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .A0 (nx8708), .A1 (
          RST), .A2 (nx8346), .B0 (nx5946), .B1 (nx6008)) ;
    oai32 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix483 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .A0 (nx5988), .A1 (
          RST), .A2 (nx8346), .B0 (nx5950), .B1 (nx6008)) ;
    oai32 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix493 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .A0 (nx6010), .A1 (
          RST), .A2 (nx8346), .B0 (nx5954), .B1 (nx6008)) ;
    inv01 ix6009 (.Y (nx6010), .A (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_10)) ;
    oai32 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix503 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .A0 (nx6012), .A1 (
          RST), .A2 (nx8346), .B0 (nx5958), .B1 (nx6008)) ;
    inv01 ix6011 (.Y (nx6012), .A (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_11)) ;
    oai32 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix513 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .A0 (nx6014), .A1 (
          RST), .A2 (nx8346), .B0 (nx5962), .B1 (nx6008)) ;
    inv01 ix6013 (.Y (nx6014), .A (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_12)) ;
    oai32 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix523 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .A0 (nx6016), .A1 (
          RST), .A2 (nx8348), .B0 (nx5966), .B1 (nx6008)) ;
    inv01 ix6015 (.Y (nx6016), .A (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_13)) ;
    oai32 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix533 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .A0 (nx6018), .A1 (
          RST), .A2 (nx8348), .B0 (nx5970), .B1 (nx6020)) ;
    inv01 ix6017 (.Y (nx6018), .A (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_14)) ;
    inv01 ix6019 (.Y (nx6020), .A (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566)) ;
    oai32 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix543 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .A0 (nx6022), .A1 (
          RST), .A2 (nx8348), .B0 (nx5974), .B1 (nx6020)) ;
    inv01 ix6021 (.Y (nx6022), .A (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_15)) ;
    oai32 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix553 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .A0 (nx6024), .A1 (
          RST), .A2 (nx8348), .B0 (nx5978), .B1 (nx6020)) ;
    inv01 ix6023 (.Y (nx6024), .A (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterSDin_16)) ;
    nand02_2x L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix633 (.Y (nx6006), .A0 (
              nx7606), .A1 (nx8348)) ;
    nand02_2x L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix635 (.Y (nx6008), .A0 (
              nx7606), .A1 (nx8348)) ;
    oai32 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix393 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .A0 (nx6026), .A1 (
          RST), .A2 (nx8350), .B0 (L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx384), .B1 (
          nx6028)) ;
    inv01 ix6025 (.Y (nx6026), .A (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_0)) ;
    oai32 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix403 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .A0 (nx6030), .A1 (
          RST), .A2 (nx8350), .B0 (nx5846), .B1 (nx6028)) ;
    inv01 ix6029 (.Y (nx6030), .A (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_1)) ;
    oai32 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix413 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .A0 (nx6032), .A1 (
          RST), .A2 (nx8350), .B0 (L1_3_L2_3_G2_MINI_ALU_nx387), .B1 (nx6028)) ;
    inv01 ix6031 (.Y (nx6032), .A (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_2)) ;
    oai32 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix423 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .A0 (nx6034), .A1 (
          RST), .A2 (nx8350), .B0 (L1_3_L2_3_G2_MINI_ALU_nx399), .B1 (nx6028)) ;
    inv01 ix6033 (.Y (nx6034), .A (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_3)) ;
    oai32 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix433 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .A0 (nx6036), .A1 (
          RST), .A2 (nx8350), .B0 (L1_3_L2_3_G2_MINI_ALU_nx409), .B1 (nx6028)) ;
    inv01 ix6035 (.Y (nx6036), .A (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_4)) ;
    oai32 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix443 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .A0 (nx6038), .A1 (
          RST), .A2 (nx8350), .B0 (L1_3_L2_3_G2_MINI_ALU_nx419), .B1 (nx6028)) ;
    inv01 ix6037 (.Y (nx6038), .A (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_5)) ;
    oai32 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix453 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .A0 (nx6040), .A1 (
          RST), .A2 (nx8350), .B0 (L1_3_L2_3_G2_MINI_ALU_nx429), .B1 (nx6028)) ;
    inv01 ix6039 (.Y (nx6040), .A (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_6)) ;
    oai32 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix463 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .A0 (nx6042), .A1 (
          RST), .A2 (nx8352), .B0 (L1_3_L2_3_G2_MINI_ALU_nx439), .B1 (nx6044)) ;
    inv01 ix6041 (.Y (nx6042), .A (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_7)) ;
    oai32 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix473 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .A0 (nx6046), .A1 (
          RST), .A2 (nx8352), .B0 (L1_3_L2_3_G2_MINI_ALU_nx449), .B1 (nx6044)) ;
    inv01 ix6045 (.Y (nx6046), .A (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_8)) ;
    oai32 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix483 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .A0 (nx6048), .A1 (
          RST), .A2 (nx8352), .B0 (L1_3_L2_3_G2_MINI_ALU_nx469), .B1 (nx6044)) ;
    inv01 ix6047 (.Y (nx6048), .A (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_9)) ;
    oai32 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix493 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .A0 (nx6050), .A1 (
          RST), .A2 (nx8352), .B0 (L1_3_L2_3_G2_MINI_ALU_nx477), .B1 (nx6044)) ;
    inv01 ix6049 (.Y (nx6050), .A (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_10)) ;
    oai32 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix503 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .A0 (nx6052), .A1 (
          RST), .A2 (nx8352), .B0 (L1_3_L2_3_G2_MINI_ALU_nx485), .B1 (nx6044)) ;
    inv01 ix6051 (.Y (nx6052), .A (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_11)) ;
    oai32 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix513 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .A0 (nx6054), .A1 (
          RST), .A2 (nx8352), .B0 (L1_3_L2_3_G2_MINI_ALU_nx493), .B1 (nx6044)) ;
    inv01 ix6053 (.Y (nx6054), .A (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_12)) ;
    oai32 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix523 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .A0 (nx6056), .A1 (
          RST), .A2 (nx8352), .B0 (L1_3_L2_3_G2_MINI_ALU_nx501), .B1 (nx6044)) ;
    inv01 ix6055 (.Y (nx6056), .A (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_13)) ;
    oai32 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix533 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .A0 (nx6058), .A1 (
          RST), .A2 (nx8354), .B0 (L1_3_L2_3_G2_MINI_ALU_nx509), .B1 (nx6060)) ;
    inv01 ix6057 (.Y (nx6058), .A (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_14)) ;
    inv01 ix6059 (.Y (nx6060), .A (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566)) ;
    oai32 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix543 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .A0 (nx6062), .A1 (
          RST), .A2 (nx8354), .B0 (L1_3_L2_3_G2_MINI_ALU_nx517), .B1 (nx6060)) ;
    inv01 ix6061 (.Y (nx6062), .A (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_15)) ;
    oai32 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix553 (.Y (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .A0 (nx6064), .A1 (
          RST), .A2 (nx8354), .B0 (nx5862), .B1 (nx6060)) ;
    inv01 ix6063 (.Y (nx6064), .A (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_RegisterPDin_16)) ;
    nand02_2x L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix633 (.Y (nx6028), .A0 (
              nx7608), .A1 (nx8354)) ;
    nand02_2x L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix635 (.Y (nx6044), .A0 (
              nx7608), .A1 (nx8354)) ;
    mux21 L1_3_L2_4_G3_MINI_ALU_ix404 (.Y (L1_3_L2_4_G3_MINI_ALU_nx403), .A0 (
          nx6066), .A1 (L1_3_L2_4_G3_MINI_ALU_BoothP_2), .S0 (
          L1_3_L2_4_G3_MINI_ALU_nx395)) ;
    inv01 ix6065 (.Y (nx6066), .A (L1_3_L2_4_G3_MINI_ALU_nx391)) ;
    mux21 L1_3_L2_4_G3_MINI_ALU_ix414 (.Y (L1_3_L2_4_G3_MINI_ALU_nx413), .A0 (
          nx6068), .A1 (L1_3_L2_4_G3_MINI_ALU_BoothP_3), .S0 (
          L1_3_L2_4_G3_MINI_ALU_nx405)) ;
    inv01 ix6067 (.Y (nx6068), .A (L1_3_L2_4_G3_MINI_ALU_nx403)) ;
    mux21 L1_3_L2_4_G3_MINI_ALU_ix424 (.Y (L1_3_L2_4_G3_MINI_ALU_nx423), .A0 (
          nx6070), .A1 (L1_3_L2_4_G3_MINI_ALU_BoothP_4), .S0 (
          L1_3_L2_4_G3_MINI_ALU_nx415)) ;
    inv01 ix6069 (.Y (nx6070), .A (L1_3_L2_4_G3_MINI_ALU_nx413)) ;
    mux21 L1_3_L2_4_G3_MINI_ALU_ix434 (.Y (L1_3_L2_4_G3_MINI_ALU_nx433), .A0 (
          nx6072), .A1 (L1_3_L2_4_G3_MINI_ALU_BoothP_5), .S0 (
          L1_3_L2_4_G3_MINI_ALU_nx425)) ;
    inv01 ix6071 (.Y (nx6072), .A (L1_3_L2_4_G3_MINI_ALU_nx423)) ;
    mux21 L1_3_L2_4_G3_MINI_ALU_ix444 (.Y (L1_3_L2_4_G3_MINI_ALU_nx443), .A0 (
          nx6074), .A1 (L1_3_L2_4_G3_MINI_ALU_BoothP_6), .S0 (
          L1_3_L2_4_G3_MINI_ALU_nx435)) ;
    inv01 ix6073 (.Y (nx6074), .A (L1_3_L2_4_G3_MINI_ALU_nx433)) ;
    mux21 L1_3_L2_4_G3_MINI_ALU_ix454 (.Y (L1_3_L2_4_G3_MINI_ALU_nx453), .A0 (
          nx6076), .A1 (L1_3_L2_4_G3_MINI_ALU_BoothP_7), .S0 (
          L1_3_L2_4_G3_MINI_ALU_nx445)) ;
    inv01 ix6075 (.Y (nx6076), .A (L1_3_L2_4_G3_MINI_ALU_nx443)) ;
    mux21 L1_3_L2_4_G3_MINI_ALU_ix462 (.Y (L1_3_L2_4_G3_MINI_ALU_nx461), .A0 (
          nx6078), .A1 (L1_3_L2_4_G3_MINI_ALU_BoothP_8), .S0 (
          L1_3_L2_4_G3_MINI_ALU_nx455)) ;
    inv01 ix6077 (.Y (nx6078), .A (L1_3_L2_4_G3_MINI_ALU_nx453)) ;
    mux21 L1_3_L2_4_G3_MINI_ALU_ix468 (.Y (L1_3_L2_4_G3_MINI_ALU_nx467), .A0 (
          nx6080), .A1 (L1_3_L2_4_G3_MINI_ALU_BoothP_9), .S0 (
          L1_3_L2_4_G3_MINI_ALU_nx463)) ;
    inv01 ix6079 (.Y (nx6080), .A (L1_3_L2_4_G3_MINI_ALU_nx461)) ;
    mux21 L1_3_L2_4_G3_MINI_ALU_ix476 (.Y (L1_3_L2_4_G3_MINI_ALU_nx475), .A0 (
          nx6082), .A1 (L1_3_L2_4_G3_MINI_ALU_BoothP_10), .S0 (
          L1_3_L2_4_G3_MINI_ALU_nx471)) ;
    inv01 ix6081 (.Y (nx6082), .A (L1_3_L2_4_G3_MINI_ALU_nx467)) ;
    mux21 L1_3_L2_4_G3_MINI_ALU_ix484 (.Y (L1_3_L2_4_G3_MINI_ALU_nx483), .A0 (
          nx6084), .A1 (L1_3_L2_4_G3_MINI_ALU_BoothP_11), .S0 (
          L1_3_L2_4_G3_MINI_ALU_nx479)) ;
    inv01 ix6083 (.Y (nx6084), .A (L1_3_L2_4_G3_MINI_ALU_nx475)) ;
    mux21 L1_3_L2_4_G3_MINI_ALU_ix492 (.Y (L1_3_L2_4_G3_MINI_ALU_nx491), .A0 (
          nx6086), .A1 (L1_3_L2_4_G3_MINI_ALU_BoothP_12), .S0 (
          L1_3_L2_4_G3_MINI_ALU_nx487)) ;
    inv01 ix6085 (.Y (nx6086), .A (L1_3_L2_4_G3_MINI_ALU_nx483)) ;
    mux21 L1_3_L2_4_G3_MINI_ALU_ix500 (.Y (L1_3_L2_4_G3_MINI_ALU_nx499), .A0 (
          nx6088), .A1 (L1_3_L2_4_G3_MINI_ALU_BoothP_13), .S0 (
          L1_3_L2_4_G3_MINI_ALU_nx495)) ;
    inv01 ix6087 (.Y (nx6088), .A (L1_3_L2_4_G3_MINI_ALU_nx491)) ;
    mux21 L1_3_L2_4_G3_MINI_ALU_ix508 (.Y (L1_3_L2_4_G3_MINI_ALU_nx507), .A0 (
          nx6090), .A1 (L1_3_L2_4_G3_MINI_ALU_BoothP_14), .S0 (
          L1_3_L2_4_G3_MINI_ALU_nx503)) ;
    inv01 ix6089 (.Y (nx6090), .A (L1_3_L2_4_G3_MINI_ALU_nx499)) ;
    mux21 L1_3_L2_4_G3_MINI_ALU_ix516 (.Y (L1_3_L2_4_G3_MINI_ALU_nx515), .A0 (
          nx6092), .A1 (L1_3_L2_4_G3_MINI_ALU_BoothP_15), .S0 (
          L1_3_L2_4_G3_MINI_ALU_nx511)) ;
    inv01 ix6091 (.Y (nx6092), .A (L1_3_L2_4_G3_MINI_ALU_nx507)) ;
    mux21 L1_3_L2_4_G3_MINI_ALU_ix161 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_1), .A0 (nx6094), .A1 (
          L1_3_L2_4_G3_MINI_ALU_nx379), .S0 (nx8358)) ;
    inv01 ix6093 (.Y (nx6094), .A (L1_3_L2_4_G3_MINI_ALU_BoothP_1)) ;
    mux21 L1_3_L2_4_G3_MINI_ALU_ix181 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_2), .A0 (
          L1_3_L2_4_G3_MINI_ALU_nx387), .A1 (L1_3_L2_4_G3_MINI_ALU_nx389), .S0 (
          nx8358)) ;
    mux21 L1_3_L2_4_G3_MINI_ALU_ix201 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_3), .A0 (
          L1_3_L2_4_G3_MINI_ALU_nx399), .A1 (L1_3_L2_4_G3_MINI_ALU_nx401), .S0 (
          nx8358)) ;
    mux21 L1_3_L2_4_G3_MINI_ALU_ix221 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_4), .A0 (
          L1_3_L2_4_G3_MINI_ALU_nx409), .A1 (L1_3_L2_4_G3_MINI_ALU_nx411), .S0 (
          nx8358)) ;
    mux21 L1_3_L2_4_G3_MINI_ALU_ix241 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_5), .A0 (
          L1_3_L2_4_G3_MINI_ALU_nx419), .A1 (L1_3_L2_4_G3_MINI_ALU_nx421), .S0 (
          nx8358)) ;
    mux21 L1_3_L2_4_G3_MINI_ALU_ix261 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_6), .A0 (
          L1_3_L2_4_G3_MINI_ALU_nx429), .A1 (L1_3_L2_4_G3_MINI_ALU_nx431), .S0 (
          nx8358)) ;
    mux21 L1_3_L2_4_G3_MINI_ALU_ix281 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_7), .A0 (
          L1_3_L2_4_G3_MINI_ALU_nx439), .A1 (L1_3_L2_4_G3_MINI_ALU_nx441), .S0 (
          nx8358)) ;
    mux21 L1_3_L2_4_G3_MINI_ALU_ix301 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_8), .A0 (
          L1_3_L2_4_G3_MINI_ALU_nx449), .A1 (L1_3_L2_4_G3_MINI_ALU_nx451), .S0 (
          nx8360)) ;
    mux21 L1_3_L2_4_G3_MINI_ALU_ix321 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_9), .A0 (
          L1_3_L2_4_G3_MINI_ALU_nx469), .A1 (nx6096), .S0 (nx8360)) ;
    inv01 ix6095 (.Y (nx6096), .A (L1_3_L2_4_G3_MINI_ALU_nx316)) ;
    mux21 L1_3_L2_4_G3_MINI_ALU_ix341 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_10), .A0 (
          L1_3_L2_4_G3_MINI_ALU_nx477), .A1 (nx6098), .S0 (nx8360)) ;
    inv01 ix6097 (.Y (nx6098), .A (L1_3_L2_4_G3_MINI_ALU_nx336)) ;
    mux21 L1_3_L2_4_G3_MINI_ALU_ix361 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_11), .A0 (
          L1_3_L2_4_G3_MINI_ALU_nx485), .A1 (nx6100), .S0 (nx8360)) ;
    inv01 ix6099 (.Y (nx6100), .A (L1_3_L2_4_G3_MINI_ALU_nx356)) ;
    mux21 L1_3_L2_4_G3_MINI_ALU_ix381 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_12), .A0 (
          L1_3_L2_4_G3_MINI_ALU_nx493), .A1 (nx6102), .S0 (nx8360)) ;
    inv01 ix6101 (.Y (nx6102), .A (L1_3_L2_4_G3_MINI_ALU_nx376)) ;
    mux21 L1_3_L2_4_G3_MINI_ALU_ix401 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_13), .A0 (
          L1_3_L2_4_G3_MINI_ALU_nx501), .A1 (nx6104), .S0 (nx8360)) ;
    inv01 ix6103 (.Y (nx6104), .A (L1_3_L2_4_G3_MINI_ALU_nx396)) ;
    mux21 L1_3_L2_4_G3_MINI_ALU_ix421 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_14), .A0 (
          L1_3_L2_4_G3_MINI_ALU_nx509), .A1 (nx6106), .S0 (nx8360)) ;
    inv01 ix6105 (.Y (nx6106), .A (L1_3_L2_4_G3_MINI_ALU_nx416)) ;
    mux21 L1_3_L2_4_G3_MINI_ALU_ix441 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_15), .A0 (
          L1_3_L2_4_G3_MINI_ALU_nx517), .A1 (nx6108), .S0 (nx8362)) ;
    inv01 ix6107 (.Y (nx6108), .A (L1_3_L2_4_G3_MINI_ALU_nx436)) ;
    mux21 L1_3_L2_4_G3_MINI_ALU_ix461 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_16), .A0 (nx6110), .A1 (nx6112
          ), .S0 (nx8362)) ;
    inv01 ix6109 (.Y (nx6110), .A (L1_3_L2_4_G3_MINI_ALU_BoothP_16)) ;
    inv01 ix6111 (.Y (nx6112), .A (L1_3_L2_4_G3_MINI_ALU_nx456)) ;
    nor02_2x L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix319 (.Y (
             L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642), .A0 (Start), .A1 (
             CalculatingBooth_dup_1162)) ;
    nor02_2x L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix85 (.Y (
             L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_0), .A0 (nx8372), .A1 (
             nx6114)) ;
    inv01 ix6113 (.Y (nx6114), .A (L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_1)) ;
    mux21 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix125 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_1), .A0 (nx6116), .A1 (
          nx6118), .S0 (nx8372)) ;
    inv01 ix6115 (.Y (nx6116), .A (L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_2)) ;
    inv01 ix6117 (.Y (nx6118), .A (WindowDin_3__4__0)) ;
    mux21 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix133 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_2), .A0 (nx6120), .A1 (
          nx6122), .S0 (nx8372)) ;
    inv01 ix6119 (.Y (nx6120), .A (L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_3)) ;
    inv01 ix6121 (.Y (nx6122), .A (WindowDin_3__4__1)) ;
    mux21 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix141 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_3), .A0 (nx6124), .A1 (
          nx6126), .S0 (nx8372)) ;
    inv01 ix6123 (.Y (nx6124), .A (L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_4)) ;
    inv01 ix6125 (.Y (nx6126), .A (WindowDin_3__4__2)) ;
    mux21 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix149 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_4), .A0 (nx6128), .A1 (
          nx6130), .S0 (nx8372)) ;
    inv01 ix6127 (.Y (nx6128), .A (L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_5)) ;
    inv01 ix6129 (.Y (nx6130), .A (WindowDin_3__4__3)) ;
    mux21 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix157 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_5), .A0 (nx6132), .A1 (
          nx6134), .S0 (nx8372)) ;
    inv01 ix6131 (.Y (nx6132), .A (L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_6)) ;
    inv01 ix6133 (.Y (nx6134), .A (WindowDin_3__4__4)) ;
    mux21 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix165 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_6), .A0 (nx6136), .A1 (
          nx6138), .S0 (nx8372)) ;
    inv01 ix6135 (.Y (nx6136), .A (L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_7)) ;
    inv01 ix6137 (.Y (nx6138), .A (WindowDin_3__4__5)) ;
    mux21 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix173 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_7), .A0 (nx6140), .A1 (
          nx6142), .S0 (nx8374)) ;
    inv01 ix6139 (.Y (nx6140), .A (L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_8)) ;
    inv01 ix6141 (.Y (nx6142), .A (WindowDin_3__4__6)) ;
    mux21 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix181 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_8), .A0 (nx6144), .A1 (
          nx6146), .S0 (nx8374)) ;
    inv01 ix6143 (.Y (nx6144), .A (L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_9)) ;
    inv01 ix6145 (.Y (nx6146), .A (WindowDin_3__4__7)) ;
    nor02_2x L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix89 (.Y (
             L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_9), .A0 (nx8374), .A1 (
             nx6148)) ;
    inv01 ix6147 (.Y (nx6148), .A (L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_10)
          ) ;
    nor02_2x L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix93 (.Y (
             L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_10), .A0 (nx8374), .A1 (
             nx6150)) ;
    inv01 ix6149 (.Y (nx6150), .A (L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_11)
          ) ;
    nor02_2x L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix97 (.Y (
             L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_11), .A0 (nx8374), .A1 (
             nx6152)) ;
    inv01 ix6151 (.Y (nx6152), .A (L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_12)
          ) ;
    nor02_2x L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix101 (.Y (
             L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_12), .A0 (nx8374), .A1 (
             nx6154)) ;
    inv01 ix6153 (.Y (nx6154), .A (L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_13)
          ) ;
    nor02_2x L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix105 (.Y (
             L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_13), .A0 (nx8374), .A1 (
             nx6156)) ;
    inv01 ix6155 (.Y (nx6156), .A (L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_14)
          ) ;
    nor02_2x L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix109 (.Y (
             L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_14), .A0 (nx8376), .A1 (
             nx6158)) ;
    inv01 ix6157 (.Y (nx6158), .A (L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_15)
          ) ;
    nor02_2x L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix113 (.Y (
             L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_15), .A0 (nx8376), .A1 (
             nx6160)) ;
    inv01 ix6159 (.Y (nx6160), .A (L1_3_L2_4_G3_MINI_ALU_BoothPBeforeShift_16)
          ) ;
    nor02_2x L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix117 (.Y (
             L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_16), .A0 (nx8376), .A1 (
             nx6160)) ;
    mux21 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix189 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BoothOperand_0), .A0 (nx6162), .A1 (nx6164), .S0 (
          nx8364)) ;
    inv01 ix6161 (.Y (nx6162), .A (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_0)) ;
    inv01 ix6163 (.Y (nx6164), .A (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_0)) ;
    mux21 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix197 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BoothOperand_1), .A0 (nx6166), .A1 (nx6168), .S0 (
          nx8364)) ;
    inv01 ix6165 (.Y (nx6166), .A (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_1)) ;
    inv01 ix6167 (.Y (nx6168), .A (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_1)) ;
    mux21 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix205 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BoothOperand_2), .A0 (nx6170), .A1 (nx6172), .S0 (
          nx8364)) ;
    inv01 ix6169 (.Y (nx6170), .A (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_2)) ;
    inv01 ix6171 (.Y (nx6172), .A (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_2)) ;
    mux21 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix213 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BoothOperand_3), .A0 (nx6174), .A1 (nx6176), .S0 (
          nx8364)) ;
    inv01 ix6173 (.Y (nx6174), .A (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_3)) ;
    inv01 ix6175 (.Y (nx6176), .A (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_3)) ;
    mux21 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix221 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BoothOperand_4), .A0 (nx6178), .A1 (nx6180), .S0 (
          nx8364)) ;
    inv01 ix6177 (.Y (nx6178), .A (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_4)) ;
    inv01 ix6179 (.Y (nx6180), .A (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_4)) ;
    mux21 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix229 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BoothOperand_5), .A0 (nx6182), .A1 (nx6184), .S0 (
          nx8366)) ;
    inv01 ix6181 (.Y (nx6182), .A (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_5)) ;
    inv01 ix6183 (.Y (nx6184), .A (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_5)) ;
    mux21 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix237 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BoothOperand_6), .A0 (nx6186), .A1 (nx6188), .S0 (
          nx8366)) ;
    inv01 ix6185 (.Y (nx6186), .A (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_6)) ;
    inv01 ix6187 (.Y (nx6188), .A (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_6)) ;
    mux21 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix245 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BoothOperand_7), .A0 (nx6190), .A1 (nx6192), .S0 (
          nx8366)) ;
    inv01 ix6189 (.Y (nx6190), .A (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_7)) ;
    inv01 ix6191 (.Y (nx6192), .A (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_7)) ;
    mux21 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix253 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BoothOperand_8), .A0 (nx6194), .A1 (nx6196), .S0 (
          nx8366)) ;
    inv01 ix6193 (.Y (nx6194), .A (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_8)) ;
    inv01 ix6195 (.Y (nx6196), .A (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_8)) ;
    mux21 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix261 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BoothOperand_9), .A0 (nx6198), .A1 (nx6200), .S0 (
          nx8366)) ;
    inv01 ix6197 (.Y (nx6198), .A (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_9)) ;
    inv01 ix6199 (.Y (nx6200), .A (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_9)) ;
    mux21 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix269 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BoothOperand_10), .A0 (nx6202), .A1 (nx6204), .S0 (
          nx8366)) ;
    inv01 ix6201 (.Y (nx6202), .A (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_10)) ;
    inv01 ix6203 (.Y (nx6204), .A (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_10)) ;
    mux21 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix277 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BoothOperand_11), .A0 (nx6206), .A1 (nx6208), .S0 (
          nx8366)) ;
    inv01 ix6205 (.Y (nx6206), .A (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_11)) ;
    inv01 ix6207 (.Y (nx6208), .A (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_11)) ;
    mux21 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix285 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BoothOperand_12), .A0 (nx6210), .A1 (nx6212), .S0 (
          nx8368)) ;
    inv01 ix6209 (.Y (nx6210), .A (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_12)) ;
    inv01 ix6211 (.Y (nx6212), .A (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_12)) ;
    mux21 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix293 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BoothOperand_13), .A0 (nx6214), .A1 (nx6216), .S0 (
          nx8368)) ;
    inv01 ix6213 (.Y (nx6214), .A (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_13)) ;
    inv01 ix6215 (.Y (nx6216), .A (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_13)) ;
    mux21 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix301 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BoothOperand_14), .A0 (nx6218), .A1 (nx6220), .S0 (
          nx8368)) ;
    inv01 ix6217 (.Y (nx6218), .A (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_14)) ;
    inv01 ix6219 (.Y (nx6220), .A (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_14)) ;
    mux21 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix309 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BoothOperand_15), .A0 (nx6222), .A1 (nx6224), .S0 (
          nx8368)) ;
    inv01 ix6221 (.Y (nx6222), .A (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_15)) ;
    inv01 ix6223 (.Y (nx6224), .A (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_15)) ;
    mux21 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix317 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BoothOperand_16), .A0 (nx6226), .A1 (nx6228), .S0 (
          nx8368)) ;
    inv01 ix6225 (.Y (nx6226), .A (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_16)) ;
    inv01 ix6227 (.Y (nx6228), .A (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_16)) ;
    xnor2 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_ix321 (.Y (
          L1_3_L2_4_G3_MINI_ALU_AddPToBoothOperand), .A0 (nx8368), .A1 (nx6094)
          ) ;
    oai32 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix393 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .A0 (nx8710), .A1 (
          RST), .A2 (nx8378), .B0 (nx6164), .B1 (nx6232)) ;
    oai32 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix403 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .A0 (nx8710), .A1 (
          RST), .A2 (nx8378), .B0 (nx6168), .B1 (nx6232)) ;
    oai32 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix413 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .A0 (nx8710), .A1 (
          RST), .A2 (nx8378), .B0 (nx6172), .B1 (nx6232)) ;
    oai32 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix423 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .A0 (nx8710), .A1 (
          RST), .A2 (nx8378), .B0 (nx6176), .B1 (nx6232)) ;
    oai32 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix433 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .A0 (nx8710), .A1 (
          RST), .A2 (nx8378), .B0 (nx6180), .B1 (nx6232)) ;
    oai32 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix443 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .A0 (nx8710), .A1 (
          RST), .A2 (nx8378), .B0 (nx6184), .B1 (nx6232)) ;
    oai32 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix453 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .A0 (nx8710), .A1 (
          RST), .A2 (nx8380), .B0 (nx6188), .B1 (nx6232)) ;
    oai32 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix463 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .A0 (nx8712), .A1 (
          RST), .A2 (nx8380), .B0 (nx6192), .B1 (nx6234)) ;
    oai32 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix473 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .A0 (nx8712), .A1 (
          RST), .A2 (nx8380), .B0 (nx6196), .B1 (nx6234)) ;
    oai32 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix483 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .A0 (nx6236), .A1 (
          RST), .A2 (nx8380), .B0 (nx6200), .B1 (nx6234)) ;
    inv01 ix6235 (.Y (nx6236), .A (FilterDin_3__4__0)) ;
    oai32 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix493 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .A0 (nx6238), .A1 (
          RST), .A2 (nx8380), .B0 (nx6204), .B1 (nx6234)) ;
    inv01 ix6237 (.Y (nx6238), .A (FilterDin_3__4__1)) ;
    oai32 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix503 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .A0 (nx6240), .A1 (
          RST), .A2 (nx8380), .B0 (nx6208), .B1 (nx6234)) ;
    inv01 ix6239 (.Y (nx6240), .A (FilterDin_3__4__2)) ;
    oai32 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix513 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .A0 (nx6242), .A1 (
          RST), .A2 (nx8380), .B0 (nx6212), .B1 (nx6234)) ;
    inv01 ix6241 (.Y (nx6242), .A (FilterDin_3__4__3)) ;
    oai32 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix523 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .A0 (nx6244), .A1 (
          RST), .A2 (nx8382), .B0 (nx6216), .B1 (nx6234)) ;
    inv01 ix6243 (.Y (nx6244), .A (FilterDin_3__4__4)) ;
    oai32 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix533 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .A0 (nx6246), .A1 (
          RST), .A2 (nx8382), .B0 (nx6220), .B1 (nx6248)) ;
    inv01 ix6245 (.Y (nx6246), .A (FilterDin_3__4__5)) ;
    inv01 ix6247 (.Y (nx6248), .A (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566)) ;
    oai32 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix543 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .A0 (nx6250), .A1 (
          RST), .A2 (nx8382), .B0 (nx6224), .B1 (nx6248)) ;
    inv01 ix6249 (.Y (nx6250), .A (FilterDin_3__4__6)) ;
    oai32 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix553 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .A0 (nx6252), .A1 (
          RST), .A2 (nx8382), .B0 (nx6228), .B1 (nx6248)) ;
    inv01 ix6251 (.Y (nx6252), .A (FilterDin_3__4__7)) ;
    nand02_2x L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix633 (.Y (nx6232), .A0 (
              nx7608), .A1 (nx8382)) ;
    nand02_2x L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix635 (.Y (nx6234), .A0 (
              nx7608), .A1 (nx8382)) ;
    oai32 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix393 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .A0 (nx8712), .A1 (
          RST), .A2 (nx8384), .B0 (nx6162), .B1 (nx6254)) ;
    oai32 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix403 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .A0 (nx8712), .A1 (
          RST), .A2 (nx8384), .B0 (nx6166), .B1 (nx6254)) ;
    oai32 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix413 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .A0 (nx8712), .A1 (
          RST), .A2 (nx8384), .B0 (nx6170), .B1 (nx6254)) ;
    oai32 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix423 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .A0 (nx8712), .A1 (
          RST), .A2 (nx8384), .B0 (nx6174), .B1 (nx6254)) ;
    oai32 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix433 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .A0 (nx8712), .A1 (
          RST), .A2 (nx8384), .B0 (nx6178), .B1 (nx6254)) ;
    oai32 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix443 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .A0 (nx8714), .A1 (
          RST), .A2 (nx8384), .B0 (nx6182), .B1 (nx6254)) ;
    oai32 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix453 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .A0 (nx8714), .A1 (
          RST), .A2 (nx8386), .B0 (nx6186), .B1 (nx6254)) ;
    oai32 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix463 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .A0 (nx8714), .A1 (
          RST), .A2 (nx8386), .B0 (nx6190), .B1 (nx6256)) ;
    oai32 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix473 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .A0 (nx8714), .A1 (
          RST), .A2 (nx8386), .B0 (nx6194), .B1 (nx6256)) ;
    oai32 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix483 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .A0 (nx6236), .A1 (
          RST), .A2 (nx8386), .B0 (nx6198), .B1 (nx6256)) ;
    oai32 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix493 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .A0 (nx6258), .A1 (
          RST), .A2 (nx8386), .B0 (nx6202), .B1 (nx6256)) ;
    inv01 ix6257 (.Y (nx6258), .A (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_10)) ;
    oai32 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix503 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .A0 (nx6260), .A1 (
          RST), .A2 (nx8386), .B0 (nx6206), .B1 (nx6256)) ;
    inv01 ix6259 (.Y (nx6260), .A (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_11)) ;
    oai32 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix513 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .A0 (nx6262), .A1 (
          RST), .A2 (nx8386), .B0 (nx6210), .B1 (nx6256)) ;
    inv01 ix6261 (.Y (nx6262), .A (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_12)) ;
    oai32 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix523 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .A0 (nx6264), .A1 (
          RST), .A2 (nx8388), .B0 (nx6214), .B1 (nx6256)) ;
    inv01 ix6263 (.Y (nx6264), .A (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_13)) ;
    oai32 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix533 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .A0 (nx6266), .A1 (
          RST), .A2 (nx8388), .B0 (nx6218), .B1 (nx6268)) ;
    inv01 ix6265 (.Y (nx6266), .A (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_14)) ;
    inv01 ix6267 (.Y (nx6268), .A (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566)) ;
    oai32 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix543 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .A0 (nx6270), .A1 (
          RST), .A2 (nx8388), .B0 (nx6222), .B1 (nx6268)) ;
    inv01 ix6269 (.Y (nx6270), .A (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_15)) ;
    oai32 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix553 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .A0 (nx6272), .A1 (
          RST), .A2 (nx8388), .B0 (nx6226), .B1 (nx6268)) ;
    inv01 ix6271 (.Y (nx6272), .A (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_16)) ;
    nand02_2x L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix633 (.Y (nx6254), .A0 (
              nx7608), .A1 (nx8388)) ;
    nand02_2x L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix635 (.Y (nx6256), .A0 (
              nx7608), .A1 (nx8388)) ;
    oai32 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix393 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .A0 (nx6274), .A1 (
          RST), .A2 (nx8390), .B0 (L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_nx384), .B1 (
          nx6276)) ;
    inv01 ix6273 (.Y (nx6274), .A (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_0)) ;
    oai32 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix403 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .A0 (nx6278), .A1 (
          RST), .A2 (nx8390), .B0 (nx6094), .B1 (nx6276)) ;
    inv01 ix6277 (.Y (nx6278), .A (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_1)) ;
    oai32 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix413 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .A0 (nx6280), .A1 (
          RST), .A2 (nx8390), .B0 (L1_3_L2_4_G3_MINI_ALU_nx387), .B1 (nx6276)) ;
    inv01 ix6279 (.Y (nx6280), .A (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_2)) ;
    oai32 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix423 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .A0 (nx6282), .A1 (
          RST), .A2 (nx8390), .B0 (L1_3_L2_4_G3_MINI_ALU_nx399), .B1 (nx6276)) ;
    inv01 ix6281 (.Y (nx6282), .A (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_3)) ;
    oai32 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix433 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .A0 (nx6284), .A1 (
          RST), .A2 (nx8390), .B0 (L1_3_L2_4_G3_MINI_ALU_nx409), .B1 (nx6276)) ;
    inv01 ix6283 (.Y (nx6284), .A (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_4)) ;
    oai32 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix443 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .A0 (nx6286), .A1 (
          RST), .A2 (nx8390), .B0 (L1_3_L2_4_G3_MINI_ALU_nx419), .B1 (nx6276)) ;
    inv01 ix6285 (.Y (nx6286), .A (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_5)) ;
    oai32 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix453 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .A0 (nx6288), .A1 (
          RST), .A2 (nx8390), .B0 (L1_3_L2_4_G3_MINI_ALU_nx429), .B1 (nx6276)) ;
    inv01 ix6287 (.Y (nx6288), .A (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_6)) ;
    oai32 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix463 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .A0 (nx6290), .A1 (
          RST), .A2 (nx8392), .B0 (L1_3_L2_4_G3_MINI_ALU_nx439), .B1 (nx6292)) ;
    inv01 ix6289 (.Y (nx6290), .A (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_7)) ;
    oai32 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix473 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .A0 (nx6294), .A1 (
          RST), .A2 (nx8392), .B0 (L1_3_L2_4_G3_MINI_ALU_nx449), .B1 (nx6292)) ;
    inv01 ix6293 (.Y (nx6294), .A (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_8)) ;
    oai32 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix483 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .A0 (nx6296), .A1 (
          RST), .A2 (nx8392), .B0 (L1_3_L2_4_G3_MINI_ALU_nx469), .B1 (nx6292)) ;
    inv01 ix6295 (.Y (nx6296), .A (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_9)) ;
    oai32 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix493 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .A0 (nx6298), .A1 (
          RST), .A2 (nx8392), .B0 (L1_3_L2_4_G3_MINI_ALU_nx477), .B1 (nx6292)) ;
    inv01 ix6297 (.Y (nx6298), .A (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_10)) ;
    oai32 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix503 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .A0 (nx6300), .A1 (
          RST), .A2 (nx8392), .B0 (L1_3_L2_4_G3_MINI_ALU_nx485), .B1 (nx6292)) ;
    inv01 ix6299 (.Y (nx6300), .A (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_11)) ;
    oai32 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix513 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .A0 (nx6302), .A1 (
          RST), .A2 (nx8392), .B0 (L1_3_L2_4_G3_MINI_ALU_nx493), .B1 (nx6292)) ;
    inv01 ix6301 (.Y (nx6302), .A (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_12)) ;
    oai32 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix523 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .A0 (nx6304), .A1 (
          RST), .A2 (nx8392), .B0 (L1_3_L2_4_G3_MINI_ALU_nx501), .B1 (nx6292)) ;
    inv01 ix6303 (.Y (nx6304), .A (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_13)) ;
    oai32 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix533 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .A0 (nx6306), .A1 (
          RST), .A2 (nx8394), .B0 (L1_3_L2_4_G3_MINI_ALU_nx509), .B1 (nx6308)) ;
    inv01 ix6305 (.Y (nx6306), .A (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_14)) ;
    inv01 ix6307 (.Y (nx6308), .A (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566)) ;
    oai32 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix543 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .A0 (nx6310), .A1 (
          RST), .A2 (nx8394), .B0 (L1_3_L2_4_G3_MINI_ALU_nx517), .B1 (nx6308)) ;
    inv01 ix6309 (.Y (nx6310), .A (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_15)) ;
    oai32 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix553 (.Y (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .A0 (nx6312), .A1 (
          RST), .A2 (nx8394), .B0 (nx6110), .B1 (nx6308)) ;
    inv01 ix6311 (.Y (nx6312), .A (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_16)) ;
    nand02_2x L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix633 (.Y (nx6276), .A0 (
              nx7608), .A1 (nx8394)) ;
    nand02_2x L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix635 (.Y (nx6292), .A0 (
              nx7610), .A1 (nx8394)) ;
    mux21 L1_4_L2_0_G3_MINI_ALU_ix404 (.Y (L1_4_L2_0_G3_MINI_ALU_nx403), .A0 (
          nx6314), .A1 (L1_4_L2_0_G3_MINI_ALU_BoothP_2), .S0 (
          L1_4_L2_0_G3_MINI_ALU_nx395)) ;
    inv01 ix6313 (.Y (nx6314), .A (L1_4_L2_0_G3_MINI_ALU_nx391)) ;
    mux21 L1_4_L2_0_G3_MINI_ALU_ix414 (.Y (L1_4_L2_0_G3_MINI_ALU_nx413), .A0 (
          nx6316), .A1 (L1_4_L2_0_G3_MINI_ALU_BoothP_3), .S0 (
          L1_4_L2_0_G3_MINI_ALU_nx405)) ;
    inv01 ix6315 (.Y (nx6316), .A (L1_4_L2_0_G3_MINI_ALU_nx403)) ;
    mux21 L1_4_L2_0_G3_MINI_ALU_ix424 (.Y (L1_4_L2_0_G3_MINI_ALU_nx423), .A0 (
          nx6318), .A1 (L1_4_L2_0_G3_MINI_ALU_BoothP_4), .S0 (
          L1_4_L2_0_G3_MINI_ALU_nx415)) ;
    inv01 ix6317 (.Y (nx6318), .A (L1_4_L2_0_G3_MINI_ALU_nx413)) ;
    mux21 L1_4_L2_0_G3_MINI_ALU_ix434 (.Y (L1_4_L2_0_G3_MINI_ALU_nx433), .A0 (
          nx6320), .A1 (L1_4_L2_0_G3_MINI_ALU_BoothP_5), .S0 (
          L1_4_L2_0_G3_MINI_ALU_nx425)) ;
    inv01 ix6319 (.Y (nx6320), .A (L1_4_L2_0_G3_MINI_ALU_nx423)) ;
    mux21 L1_4_L2_0_G3_MINI_ALU_ix444 (.Y (L1_4_L2_0_G3_MINI_ALU_nx443), .A0 (
          nx6322), .A1 (L1_4_L2_0_G3_MINI_ALU_BoothP_6), .S0 (
          L1_4_L2_0_G3_MINI_ALU_nx435)) ;
    inv01 ix6321 (.Y (nx6322), .A (L1_4_L2_0_G3_MINI_ALU_nx433)) ;
    mux21 L1_4_L2_0_G3_MINI_ALU_ix454 (.Y (L1_4_L2_0_G3_MINI_ALU_nx453), .A0 (
          nx6324), .A1 (L1_4_L2_0_G3_MINI_ALU_BoothP_7), .S0 (
          L1_4_L2_0_G3_MINI_ALU_nx445)) ;
    inv01 ix6323 (.Y (nx6324), .A (L1_4_L2_0_G3_MINI_ALU_nx443)) ;
    mux21 L1_4_L2_0_G3_MINI_ALU_ix462 (.Y (L1_4_L2_0_G3_MINI_ALU_nx461), .A0 (
          nx6326), .A1 (L1_4_L2_0_G3_MINI_ALU_BoothP_8), .S0 (
          L1_4_L2_0_G3_MINI_ALU_nx455)) ;
    inv01 ix6325 (.Y (nx6326), .A (L1_4_L2_0_G3_MINI_ALU_nx453)) ;
    mux21 L1_4_L2_0_G3_MINI_ALU_ix468 (.Y (L1_4_L2_0_G3_MINI_ALU_nx467), .A0 (
          nx6328), .A1 (L1_4_L2_0_G3_MINI_ALU_BoothP_9), .S0 (
          L1_4_L2_0_G3_MINI_ALU_nx463)) ;
    inv01 ix6327 (.Y (nx6328), .A (L1_4_L2_0_G3_MINI_ALU_nx461)) ;
    mux21 L1_4_L2_0_G3_MINI_ALU_ix476 (.Y (L1_4_L2_0_G3_MINI_ALU_nx475), .A0 (
          nx6330), .A1 (L1_4_L2_0_G3_MINI_ALU_BoothP_10), .S0 (
          L1_4_L2_0_G3_MINI_ALU_nx471)) ;
    inv01 ix6329 (.Y (nx6330), .A (L1_4_L2_0_G3_MINI_ALU_nx467)) ;
    mux21 L1_4_L2_0_G3_MINI_ALU_ix484 (.Y (L1_4_L2_0_G3_MINI_ALU_nx483), .A0 (
          nx6332), .A1 (L1_4_L2_0_G3_MINI_ALU_BoothP_11), .S0 (
          L1_4_L2_0_G3_MINI_ALU_nx479)) ;
    inv01 ix6331 (.Y (nx6332), .A (L1_4_L2_0_G3_MINI_ALU_nx475)) ;
    mux21 L1_4_L2_0_G3_MINI_ALU_ix492 (.Y (L1_4_L2_0_G3_MINI_ALU_nx491), .A0 (
          nx6334), .A1 (L1_4_L2_0_G3_MINI_ALU_BoothP_12), .S0 (
          L1_4_L2_0_G3_MINI_ALU_nx487)) ;
    inv01 ix6333 (.Y (nx6334), .A (L1_4_L2_0_G3_MINI_ALU_nx483)) ;
    mux21 L1_4_L2_0_G3_MINI_ALU_ix500 (.Y (L1_4_L2_0_G3_MINI_ALU_nx499), .A0 (
          nx6336), .A1 (L1_4_L2_0_G3_MINI_ALU_BoothP_13), .S0 (
          L1_4_L2_0_G3_MINI_ALU_nx495)) ;
    inv01 ix6335 (.Y (nx6336), .A (L1_4_L2_0_G3_MINI_ALU_nx491)) ;
    mux21 L1_4_L2_0_G3_MINI_ALU_ix508 (.Y (L1_4_L2_0_G3_MINI_ALU_nx507), .A0 (
          nx6338), .A1 (L1_4_L2_0_G3_MINI_ALU_BoothP_14), .S0 (
          L1_4_L2_0_G3_MINI_ALU_nx503)) ;
    inv01 ix6337 (.Y (nx6338), .A (L1_4_L2_0_G3_MINI_ALU_nx499)) ;
    mux21 L1_4_L2_0_G3_MINI_ALU_ix516 (.Y (L1_4_L2_0_G3_MINI_ALU_nx515), .A0 (
          nx6340), .A1 (L1_4_L2_0_G3_MINI_ALU_BoothP_15), .S0 (
          L1_4_L2_0_G3_MINI_ALU_nx511)) ;
    inv01 ix6339 (.Y (nx6340), .A (L1_4_L2_0_G3_MINI_ALU_nx507)) ;
    mux21 L1_4_L2_0_G3_MINI_ALU_ix161 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_1), .A0 (nx6342), .A1 (
          L1_4_L2_0_G3_MINI_ALU_nx379), .S0 (nx8398)) ;
    inv01 ix6341 (.Y (nx6342), .A (L1_4_L2_0_G3_MINI_ALU_BoothP_1)) ;
    mux21 L1_4_L2_0_G3_MINI_ALU_ix181 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_2), .A0 (
          L1_4_L2_0_G3_MINI_ALU_nx387), .A1 (L1_4_L2_0_G3_MINI_ALU_nx389), .S0 (
          nx8398)) ;
    mux21 L1_4_L2_0_G3_MINI_ALU_ix201 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_3), .A0 (
          L1_4_L2_0_G3_MINI_ALU_nx399), .A1 (L1_4_L2_0_G3_MINI_ALU_nx401), .S0 (
          nx8398)) ;
    mux21 L1_4_L2_0_G3_MINI_ALU_ix221 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_4), .A0 (
          L1_4_L2_0_G3_MINI_ALU_nx409), .A1 (L1_4_L2_0_G3_MINI_ALU_nx411), .S0 (
          nx8398)) ;
    mux21 L1_4_L2_0_G3_MINI_ALU_ix241 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_5), .A0 (
          L1_4_L2_0_G3_MINI_ALU_nx419), .A1 (L1_4_L2_0_G3_MINI_ALU_nx421), .S0 (
          nx8398)) ;
    mux21 L1_4_L2_0_G3_MINI_ALU_ix261 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_6), .A0 (
          L1_4_L2_0_G3_MINI_ALU_nx429), .A1 (L1_4_L2_0_G3_MINI_ALU_nx431), .S0 (
          nx8398)) ;
    mux21 L1_4_L2_0_G3_MINI_ALU_ix281 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_7), .A0 (
          L1_4_L2_0_G3_MINI_ALU_nx439), .A1 (L1_4_L2_0_G3_MINI_ALU_nx441), .S0 (
          nx8398)) ;
    mux21 L1_4_L2_0_G3_MINI_ALU_ix301 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_8), .A0 (
          L1_4_L2_0_G3_MINI_ALU_nx449), .A1 (L1_4_L2_0_G3_MINI_ALU_nx451), .S0 (
          nx8400)) ;
    mux21 L1_4_L2_0_G3_MINI_ALU_ix321 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_9), .A0 (
          L1_4_L2_0_G3_MINI_ALU_nx469), .A1 (nx6344), .S0 (nx8400)) ;
    inv01 ix6343 (.Y (nx6344), .A (L1_4_L2_0_G3_MINI_ALU_nx316)) ;
    mux21 L1_4_L2_0_G3_MINI_ALU_ix341 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_10), .A0 (
          L1_4_L2_0_G3_MINI_ALU_nx477), .A1 (nx6346), .S0 (nx8400)) ;
    inv01 ix6345 (.Y (nx6346), .A (L1_4_L2_0_G3_MINI_ALU_nx336)) ;
    mux21 L1_4_L2_0_G3_MINI_ALU_ix361 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_11), .A0 (
          L1_4_L2_0_G3_MINI_ALU_nx485), .A1 (nx6348), .S0 (nx8400)) ;
    inv01 ix6347 (.Y (nx6348), .A (L1_4_L2_0_G3_MINI_ALU_nx356)) ;
    mux21 L1_4_L2_0_G3_MINI_ALU_ix381 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_12), .A0 (
          L1_4_L2_0_G3_MINI_ALU_nx493), .A1 (nx6350), .S0 (nx8400)) ;
    inv01 ix6349 (.Y (nx6350), .A (L1_4_L2_0_G3_MINI_ALU_nx376)) ;
    mux21 L1_4_L2_0_G3_MINI_ALU_ix401 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_13), .A0 (
          L1_4_L2_0_G3_MINI_ALU_nx501), .A1 (nx6352), .S0 (nx8400)) ;
    inv01 ix6351 (.Y (nx6352), .A (L1_4_L2_0_G3_MINI_ALU_nx396)) ;
    mux21 L1_4_L2_0_G3_MINI_ALU_ix421 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_14), .A0 (
          L1_4_L2_0_G3_MINI_ALU_nx509), .A1 (nx6354), .S0 (nx8400)) ;
    inv01 ix6353 (.Y (nx6354), .A (L1_4_L2_0_G3_MINI_ALU_nx416)) ;
    mux21 L1_4_L2_0_G3_MINI_ALU_ix441 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_15), .A0 (
          L1_4_L2_0_G3_MINI_ALU_nx517), .A1 (nx6356), .S0 (nx8402)) ;
    inv01 ix6355 (.Y (nx6356), .A (L1_4_L2_0_G3_MINI_ALU_nx436)) ;
    mux21 L1_4_L2_0_G3_MINI_ALU_ix461 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_16), .A0 (nx6358), .A1 (nx6360
          ), .S0 (nx8402)) ;
    inv01 ix6357 (.Y (nx6358), .A (L1_4_L2_0_G3_MINI_ALU_BoothP_16)) ;
    inv01 ix6359 (.Y (nx6360), .A (L1_4_L2_0_G3_MINI_ALU_nx456)) ;
    nor02_2x L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix319 (.Y (
             L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642), .A0 (Start), .A1 (
             CalculatingBooth_dup_1162)) ;
    nor02_2x L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix85 (.Y (
             L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_0), .A0 (nx8412), .A1 (
             nx6362)) ;
    inv01 ix6361 (.Y (nx6362), .A (L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_1)) ;
    mux21 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix125 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_1), .A0 (nx6364), .A1 (
          nx6366), .S0 (nx8412)) ;
    inv01 ix6363 (.Y (nx6364), .A (L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_2)) ;
    inv01 ix6365 (.Y (nx6366), .A (WindowDin_4__0__0)) ;
    mux21 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix133 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_2), .A0 (nx6368), .A1 (
          nx6370), .S0 (nx8412)) ;
    inv01 ix6367 (.Y (nx6368), .A (L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_3)) ;
    inv01 ix6369 (.Y (nx6370), .A (WindowDin_4__0__1)) ;
    mux21 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix141 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_3), .A0 (nx6372), .A1 (
          nx6374), .S0 (nx8412)) ;
    inv01 ix6371 (.Y (nx6372), .A (L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_4)) ;
    inv01 ix6373 (.Y (nx6374), .A (WindowDin_4__0__2)) ;
    mux21 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix149 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_4), .A0 (nx6376), .A1 (
          nx6378), .S0 (nx8412)) ;
    inv01 ix6375 (.Y (nx6376), .A (L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_5)) ;
    inv01 ix6377 (.Y (nx6378), .A (WindowDin_4__0__3)) ;
    mux21 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix157 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_5), .A0 (nx6380), .A1 (
          nx6382), .S0 (nx8412)) ;
    inv01 ix6379 (.Y (nx6380), .A (L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_6)) ;
    inv01 ix6381 (.Y (nx6382), .A (WindowDin_4__0__4)) ;
    mux21 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix165 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_6), .A0 (nx6384), .A1 (
          nx6386), .S0 (nx8412)) ;
    inv01 ix6383 (.Y (nx6384), .A (L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_7)) ;
    inv01 ix6385 (.Y (nx6386), .A (WindowDin_4__0__5)) ;
    mux21 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix173 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_7), .A0 (nx6388), .A1 (
          nx6390), .S0 (nx8414)) ;
    inv01 ix6387 (.Y (nx6388), .A (L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_8)) ;
    inv01 ix6389 (.Y (nx6390), .A (WindowDin_4__0__6)) ;
    mux21 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix181 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_8), .A0 (nx6392), .A1 (
          nx6394), .S0 (nx8414)) ;
    inv01 ix6391 (.Y (nx6392), .A (L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_9)) ;
    inv01 ix6393 (.Y (nx6394), .A (WindowDin_4__0__7)) ;
    nor02_2x L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix89 (.Y (
             L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_9), .A0 (nx8414), .A1 (
             nx6396)) ;
    inv01 ix6395 (.Y (nx6396), .A (L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_10)
          ) ;
    nor02_2x L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix93 (.Y (
             L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_10), .A0 (nx8414), .A1 (
             nx6398)) ;
    inv01 ix6397 (.Y (nx6398), .A (L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_11)
          ) ;
    nor02_2x L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix97 (.Y (
             L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_11), .A0 (nx8414), .A1 (
             nx6400)) ;
    inv01 ix6399 (.Y (nx6400), .A (L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_12)
          ) ;
    nor02_2x L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix101 (.Y (
             L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_12), .A0 (nx8414), .A1 (
             nx6402)) ;
    inv01 ix6401 (.Y (nx6402), .A (L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_13)
          ) ;
    nor02_2x L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix105 (.Y (
             L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_13), .A0 (nx8414), .A1 (
             nx6404)) ;
    inv01 ix6403 (.Y (nx6404), .A (L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_14)
          ) ;
    nor02_2x L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix109 (.Y (
             L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_14), .A0 (nx8416), .A1 (
             nx6406)) ;
    inv01 ix6405 (.Y (nx6406), .A (L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_15)
          ) ;
    nor02_2x L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix113 (.Y (
             L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_15), .A0 (nx8416), .A1 (
             nx6408)) ;
    inv01 ix6407 (.Y (nx6408), .A (L1_4_L2_0_G3_MINI_ALU_BoothPBeforeShift_16)
          ) ;
    nor02_2x L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix117 (.Y (
             L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_16), .A0 (nx8416), .A1 (
             nx6408)) ;
    mux21 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix189 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BoothOperand_0), .A0 (nx6410), .A1 (nx6412), .S0 (
          nx8404)) ;
    inv01 ix6409 (.Y (nx6410), .A (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_0)) ;
    inv01 ix6411 (.Y (nx6412), .A (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_0)) ;
    mux21 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix197 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BoothOperand_1), .A0 (nx6414), .A1 (nx6416), .S0 (
          nx8404)) ;
    inv01 ix6413 (.Y (nx6414), .A (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_1)) ;
    inv01 ix6415 (.Y (nx6416), .A (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_1)) ;
    mux21 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix205 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BoothOperand_2), .A0 (nx6418), .A1 (nx6420), .S0 (
          nx8404)) ;
    inv01 ix6417 (.Y (nx6418), .A (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_2)) ;
    inv01 ix6419 (.Y (nx6420), .A (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_2)) ;
    mux21 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix213 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BoothOperand_3), .A0 (nx6422), .A1 (nx6424), .S0 (
          nx8404)) ;
    inv01 ix6421 (.Y (nx6422), .A (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_3)) ;
    inv01 ix6423 (.Y (nx6424), .A (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_3)) ;
    mux21 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix221 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BoothOperand_4), .A0 (nx6426), .A1 (nx6428), .S0 (
          nx8404)) ;
    inv01 ix6425 (.Y (nx6426), .A (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_4)) ;
    inv01 ix6427 (.Y (nx6428), .A (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_4)) ;
    mux21 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix229 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BoothOperand_5), .A0 (nx6430), .A1 (nx6432), .S0 (
          nx8406)) ;
    inv01 ix6429 (.Y (nx6430), .A (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_5)) ;
    inv01 ix6431 (.Y (nx6432), .A (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_5)) ;
    mux21 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix237 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BoothOperand_6), .A0 (nx6434), .A1 (nx6436), .S0 (
          nx8406)) ;
    inv01 ix6433 (.Y (nx6434), .A (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_6)) ;
    inv01 ix6435 (.Y (nx6436), .A (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_6)) ;
    mux21 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix245 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BoothOperand_7), .A0 (nx6438), .A1 (nx6440), .S0 (
          nx8406)) ;
    inv01 ix6437 (.Y (nx6438), .A (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_7)) ;
    inv01 ix6439 (.Y (nx6440), .A (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_7)) ;
    mux21 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix253 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BoothOperand_8), .A0 (nx6442), .A1 (nx6444), .S0 (
          nx8406)) ;
    inv01 ix6441 (.Y (nx6442), .A (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_8)) ;
    inv01 ix6443 (.Y (nx6444), .A (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_8)) ;
    mux21 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix261 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BoothOperand_9), .A0 (nx6446), .A1 (nx6448), .S0 (
          nx8406)) ;
    inv01 ix6445 (.Y (nx6446), .A (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_9)) ;
    inv01 ix6447 (.Y (nx6448), .A (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_9)) ;
    mux21 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix269 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BoothOperand_10), .A0 (nx6450), .A1 (nx6452), .S0 (
          nx8406)) ;
    inv01 ix6449 (.Y (nx6450), .A (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_10)) ;
    inv01 ix6451 (.Y (nx6452), .A (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_10)) ;
    mux21 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix277 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BoothOperand_11), .A0 (nx6454), .A1 (nx6456), .S0 (
          nx8406)) ;
    inv01 ix6453 (.Y (nx6454), .A (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_11)) ;
    inv01 ix6455 (.Y (nx6456), .A (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_11)) ;
    mux21 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix285 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BoothOperand_12), .A0 (nx6458), .A1 (nx6460), .S0 (
          nx8408)) ;
    inv01 ix6457 (.Y (nx6458), .A (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_12)) ;
    inv01 ix6459 (.Y (nx6460), .A (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_12)) ;
    mux21 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix293 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BoothOperand_13), .A0 (nx6462), .A1 (nx6464), .S0 (
          nx8408)) ;
    inv01 ix6461 (.Y (nx6462), .A (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_13)) ;
    inv01 ix6463 (.Y (nx6464), .A (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_13)) ;
    mux21 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix301 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BoothOperand_14), .A0 (nx6466), .A1 (nx6468), .S0 (
          nx8408)) ;
    inv01 ix6465 (.Y (nx6466), .A (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_14)) ;
    inv01 ix6467 (.Y (nx6468), .A (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_14)) ;
    mux21 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix309 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BoothOperand_15), .A0 (nx6470), .A1 (nx6472), .S0 (
          nx8408)) ;
    inv01 ix6469 (.Y (nx6470), .A (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_15)) ;
    inv01 ix6471 (.Y (nx6472), .A (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_15)) ;
    mux21 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix317 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BoothOperand_16), .A0 (nx6474), .A1 (nx6476), .S0 (
          nx8408)) ;
    inv01 ix6473 (.Y (nx6474), .A (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_16)) ;
    inv01 ix6475 (.Y (nx6476), .A (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_16)) ;
    xnor2 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_ix321 (.Y (
          L1_4_L2_0_G3_MINI_ALU_AddPToBoothOperand), .A0 (nx8408), .A1 (nx6342)
          ) ;
    oai32 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix393 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .A0 (nx8716), .A1 (
          RST), .A2 (nx8418), .B0 (nx6412), .B1 (nx6480)) ;
    oai32 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix403 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .A0 (nx8716), .A1 (
          RST), .A2 (nx8418), .B0 (nx6416), .B1 (nx6480)) ;
    oai32 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix413 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .A0 (nx8716), .A1 (
          RST), .A2 (nx8418), .B0 (nx6420), .B1 (nx6480)) ;
    oai32 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix423 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .A0 (nx8716), .A1 (
          RST), .A2 (nx8418), .B0 (nx6424), .B1 (nx6480)) ;
    oai32 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix433 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .A0 (nx8716), .A1 (
          RST), .A2 (nx8418), .B0 (nx6428), .B1 (nx6480)) ;
    oai32 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix443 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .A0 (nx8716), .A1 (
          RST), .A2 (nx8418), .B0 (nx6432), .B1 (nx6480)) ;
    oai32 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix453 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .A0 (nx8716), .A1 (
          RST), .A2 (nx8420), .B0 (nx6436), .B1 (nx6480)) ;
    oai32 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix463 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .A0 (nx8718), .A1 (
          RST), .A2 (nx8420), .B0 (nx6440), .B1 (nx6482)) ;
    oai32 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix473 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .A0 (nx8718), .A1 (
          RST), .A2 (nx8420), .B0 (nx6444), .B1 (nx6482)) ;
    oai32 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix483 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .A0 (nx6484), .A1 (
          RST), .A2 (nx8420), .B0 (nx6448), .B1 (nx6482)) ;
    inv01 ix6483 (.Y (nx6484), .A (FilterDin_4__0__0)) ;
    oai32 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix493 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .A0 (nx6486), .A1 (
          RST), .A2 (nx8420), .B0 (nx6452), .B1 (nx6482)) ;
    inv01 ix6485 (.Y (nx6486), .A (FilterDin_4__0__1)) ;
    oai32 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix503 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .A0 (nx6488), .A1 (
          RST), .A2 (nx8420), .B0 (nx6456), .B1 (nx6482)) ;
    inv01 ix6487 (.Y (nx6488), .A (FilterDin_4__0__2)) ;
    oai32 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix513 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .A0 (nx6490), .A1 (
          RST), .A2 (nx8420), .B0 (nx6460), .B1 (nx6482)) ;
    inv01 ix6489 (.Y (nx6490), .A (FilterDin_4__0__3)) ;
    oai32 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix523 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .A0 (nx6492), .A1 (
          RST), .A2 (nx8422), .B0 (nx6464), .B1 (nx6482)) ;
    inv01 ix6491 (.Y (nx6492), .A (FilterDin_4__0__4)) ;
    oai32 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix533 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .A0 (nx6494), .A1 (
          RST), .A2 (nx8422), .B0 (nx6468), .B1 (nx6496)) ;
    inv01 ix6493 (.Y (nx6494), .A (FilterDin_4__0__5)) ;
    inv01 ix6495 (.Y (nx6496), .A (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566)) ;
    oai32 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix543 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .A0 (nx6498), .A1 (
          RST), .A2 (nx8422), .B0 (nx6472), .B1 (nx6496)) ;
    inv01 ix6497 (.Y (nx6498), .A (FilterDin_4__0__6)) ;
    oai32 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix553 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .A0 (nx6500), .A1 (
          RST), .A2 (nx8422), .B0 (nx6476), .B1 (nx6496)) ;
    inv01 ix6499 (.Y (nx6500), .A (FilterDin_4__0__7)) ;
    nand02_2x L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix633 (.Y (nx6480), .A0 (
              nx7610), .A1 (nx8422)) ;
    nand02_2x L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix635 (.Y (nx6482), .A0 (
              nx7610), .A1 (nx8422)) ;
    oai32 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix393 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .A0 (nx8718), .A1 (
          RST), .A2 (nx8424), .B0 (nx6410), .B1 (nx6502)) ;
    oai32 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix403 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .A0 (nx8718), .A1 (
          RST), .A2 (nx8424), .B0 (nx6414), .B1 (nx6502)) ;
    oai32 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix413 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .A0 (nx8718), .A1 (
          RST), .A2 (nx8424), .B0 (nx6418), .B1 (nx6502)) ;
    oai32 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix423 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .A0 (nx8718), .A1 (
          RST), .A2 (nx8424), .B0 (nx6422), .B1 (nx6502)) ;
    oai32 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix433 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .A0 (nx8718), .A1 (
          RST), .A2 (nx8424), .B0 (nx6426), .B1 (nx6502)) ;
    oai32 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix443 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .A0 (nx8720), .A1 (
          RST), .A2 (nx8424), .B0 (nx6430), .B1 (nx6502)) ;
    oai32 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix453 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .A0 (nx8720), .A1 (
          RST), .A2 (nx8426), .B0 (nx6434), .B1 (nx6502)) ;
    oai32 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix463 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .A0 (nx8720), .A1 (
          RST), .A2 (nx8426), .B0 (nx6438), .B1 (nx6504)) ;
    oai32 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix473 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .A0 (nx8720), .A1 (
          RST), .A2 (nx8426), .B0 (nx6442), .B1 (nx6504)) ;
    oai32 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix483 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .A0 (nx6484), .A1 (
          RST), .A2 (nx8426), .B0 (nx6446), .B1 (nx6504)) ;
    oai32 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix493 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .A0 (nx6506), .A1 (
          RST), .A2 (nx8426), .B0 (nx6450), .B1 (nx6504)) ;
    inv01 ix6505 (.Y (nx6506), .A (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_10)) ;
    oai32 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix503 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .A0 (nx6508), .A1 (
          RST), .A2 (nx8426), .B0 (nx6454), .B1 (nx6504)) ;
    inv01 ix6507 (.Y (nx6508), .A (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_11)) ;
    oai32 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix513 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .A0 (nx6510), .A1 (
          RST), .A2 (nx8426), .B0 (nx6458), .B1 (nx6504)) ;
    inv01 ix6509 (.Y (nx6510), .A (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_12)) ;
    oai32 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix523 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .A0 (nx6512), .A1 (
          RST), .A2 (nx8428), .B0 (nx6462), .B1 (nx6504)) ;
    inv01 ix6511 (.Y (nx6512), .A (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_13)) ;
    oai32 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix533 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .A0 (nx6514), .A1 (
          RST), .A2 (nx8428), .B0 (nx6466), .B1 (nx6516)) ;
    inv01 ix6513 (.Y (nx6514), .A (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_14)) ;
    inv01 ix6515 (.Y (nx6516), .A (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566)) ;
    oai32 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix543 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .A0 (nx6518), .A1 (
          RST), .A2 (nx8428), .B0 (nx6470), .B1 (nx6516)) ;
    inv01 ix6517 (.Y (nx6518), .A (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_15)) ;
    oai32 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix553 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .A0 (nx6520), .A1 (
          RST), .A2 (nx8428), .B0 (nx6474), .B1 (nx6516)) ;
    inv01 ix6519 (.Y (nx6520), .A (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_16)) ;
    nand02_2x L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix633 (.Y (nx6502), .A0 (
              nx7610), .A1 (nx8428)) ;
    nand02_2x L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix635 (.Y (nx6504), .A0 (
              nx7610), .A1 (nx8428)) ;
    oai32 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix393 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .A0 (nx6522), .A1 (
          RST), .A2 (nx8430), .B0 (L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_nx384), .B1 (
          nx6524)) ;
    inv01 ix6521 (.Y (nx6522), .A (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_0)) ;
    oai32 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix403 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .A0 (nx6526), .A1 (
          RST), .A2 (nx8430), .B0 (nx6342), .B1 (nx6524)) ;
    inv01 ix6525 (.Y (nx6526), .A (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_1)) ;
    oai32 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix413 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .A0 (nx6528), .A1 (
          RST), .A2 (nx8430), .B0 (L1_4_L2_0_G3_MINI_ALU_nx387), .B1 (nx6524)) ;
    inv01 ix6527 (.Y (nx6528), .A (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_2)) ;
    oai32 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix423 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .A0 (nx6530), .A1 (
          RST), .A2 (nx8430), .B0 (L1_4_L2_0_G3_MINI_ALU_nx399), .B1 (nx6524)) ;
    inv01 ix6529 (.Y (nx6530), .A (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_3)) ;
    oai32 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix433 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .A0 (nx6532), .A1 (
          RST), .A2 (nx8430), .B0 (L1_4_L2_0_G3_MINI_ALU_nx409), .B1 (nx6524)) ;
    inv01 ix6531 (.Y (nx6532), .A (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_4)) ;
    oai32 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix443 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .A0 (nx6534), .A1 (
          RST), .A2 (nx8430), .B0 (L1_4_L2_0_G3_MINI_ALU_nx419), .B1 (nx6524)) ;
    inv01 ix6533 (.Y (nx6534), .A (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_5)) ;
    oai32 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix453 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .A0 (nx6536), .A1 (
          RST), .A2 (nx8430), .B0 (L1_4_L2_0_G3_MINI_ALU_nx429), .B1 (nx6524)) ;
    inv01 ix6535 (.Y (nx6536), .A (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_6)) ;
    oai32 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix463 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .A0 (nx6538), .A1 (
          RST), .A2 (nx8432), .B0 (L1_4_L2_0_G3_MINI_ALU_nx439), .B1 (nx6540)) ;
    inv01 ix6537 (.Y (nx6538), .A (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_7)) ;
    oai32 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix473 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .A0 (nx6542), .A1 (
          RST), .A2 (nx8432), .B0 (L1_4_L2_0_G3_MINI_ALU_nx449), .B1 (nx6540)) ;
    inv01 ix6541 (.Y (nx6542), .A (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_8)) ;
    oai32 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix483 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .A0 (nx6544), .A1 (
          RST), .A2 (nx8432), .B0 (L1_4_L2_0_G3_MINI_ALU_nx469), .B1 (nx6540)) ;
    inv01 ix6543 (.Y (nx6544), .A (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_9)) ;
    oai32 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix493 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .A0 (nx6546), .A1 (
          RST), .A2 (nx8432), .B0 (L1_4_L2_0_G3_MINI_ALU_nx477), .B1 (nx6540)) ;
    inv01 ix6545 (.Y (nx6546), .A (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_10)) ;
    oai32 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix503 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .A0 (nx6548), .A1 (
          RST), .A2 (nx8432), .B0 (L1_4_L2_0_G3_MINI_ALU_nx485), .B1 (nx6540)) ;
    inv01 ix6547 (.Y (nx6548), .A (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_11)) ;
    oai32 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix513 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .A0 (nx6550), .A1 (
          RST), .A2 (nx8432), .B0 (L1_4_L2_0_G3_MINI_ALU_nx493), .B1 (nx6540)) ;
    inv01 ix6549 (.Y (nx6550), .A (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_12)) ;
    oai32 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix523 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .A0 (nx6552), .A1 (
          RST), .A2 (nx8432), .B0 (L1_4_L2_0_G3_MINI_ALU_nx501), .B1 (nx6540)) ;
    inv01 ix6551 (.Y (nx6552), .A (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_13)) ;
    oai32 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix533 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .A0 (nx6554), .A1 (
          RST), .A2 (nx8434), .B0 (L1_4_L2_0_G3_MINI_ALU_nx509), .B1 (nx6556)) ;
    inv01 ix6553 (.Y (nx6554), .A (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_14)) ;
    inv01 ix6555 (.Y (nx6556), .A (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566)) ;
    oai32 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix543 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .A0 (nx6558), .A1 (
          RST), .A2 (nx8434), .B0 (L1_4_L2_0_G3_MINI_ALU_nx517), .B1 (nx6556)) ;
    inv01 ix6557 (.Y (nx6558), .A (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_15)) ;
    oai32 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix553 (.Y (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .A0 (nx6560), .A1 (
          RST), .A2 (nx8434), .B0 (nx6358), .B1 (nx6556)) ;
    inv01 ix6559 (.Y (nx6560), .A (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_16)) ;
    nand02_2x L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix633 (.Y (nx6524), .A0 (
              nx7610), .A1 (nx8434)) ;
    nand02_2x L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix635 (.Y (nx6540), .A0 (
              nx7610), .A1 (nx8434)) ;
    mux21 L1_4_L2_1_G3_MINI_ALU_ix404 (.Y (L1_4_L2_1_G3_MINI_ALU_nx403), .A0 (
          nx6562), .A1 (L1_4_L2_1_G3_MINI_ALU_BoothP_2), .S0 (
          L1_4_L2_1_G3_MINI_ALU_nx395)) ;
    inv01 ix6561 (.Y (nx6562), .A (L1_4_L2_1_G3_MINI_ALU_nx391)) ;
    mux21 L1_4_L2_1_G3_MINI_ALU_ix414 (.Y (L1_4_L2_1_G3_MINI_ALU_nx413), .A0 (
          nx6564), .A1 (L1_4_L2_1_G3_MINI_ALU_BoothP_3), .S0 (
          L1_4_L2_1_G3_MINI_ALU_nx405)) ;
    inv01 ix6563 (.Y (nx6564), .A (L1_4_L2_1_G3_MINI_ALU_nx403)) ;
    mux21 L1_4_L2_1_G3_MINI_ALU_ix424 (.Y (L1_4_L2_1_G3_MINI_ALU_nx423), .A0 (
          nx6566), .A1 (L1_4_L2_1_G3_MINI_ALU_BoothP_4), .S0 (
          L1_4_L2_1_G3_MINI_ALU_nx415)) ;
    inv01 ix6565 (.Y (nx6566), .A (L1_4_L2_1_G3_MINI_ALU_nx413)) ;
    mux21 L1_4_L2_1_G3_MINI_ALU_ix434 (.Y (L1_4_L2_1_G3_MINI_ALU_nx433), .A0 (
          nx6568), .A1 (L1_4_L2_1_G3_MINI_ALU_BoothP_5), .S0 (
          L1_4_L2_1_G3_MINI_ALU_nx425)) ;
    inv01 ix6567 (.Y (nx6568), .A (L1_4_L2_1_G3_MINI_ALU_nx423)) ;
    mux21 L1_4_L2_1_G3_MINI_ALU_ix444 (.Y (L1_4_L2_1_G3_MINI_ALU_nx443), .A0 (
          nx6570), .A1 (L1_4_L2_1_G3_MINI_ALU_BoothP_6), .S0 (
          L1_4_L2_1_G3_MINI_ALU_nx435)) ;
    inv01 ix6569 (.Y (nx6570), .A (L1_4_L2_1_G3_MINI_ALU_nx433)) ;
    mux21 L1_4_L2_1_G3_MINI_ALU_ix454 (.Y (L1_4_L2_1_G3_MINI_ALU_nx453), .A0 (
          nx6572), .A1 (L1_4_L2_1_G3_MINI_ALU_BoothP_7), .S0 (
          L1_4_L2_1_G3_MINI_ALU_nx445)) ;
    inv01 ix6571 (.Y (nx6572), .A (L1_4_L2_1_G3_MINI_ALU_nx443)) ;
    mux21 L1_4_L2_1_G3_MINI_ALU_ix462 (.Y (L1_4_L2_1_G3_MINI_ALU_nx461), .A0 (
          nx6574), .A1 (L1_4_L2_1_G3_MINI_ALU_BoothP_8), .S0 (
          L1_4_L2_1_G3_MINI_ALU_nx455)) ;
    inv01 ix6573 (.Y (nx6574), .A (L1_4_L2_1_G3_MINI_ALU_nx453)) ;
    mux21 L1_4_L2_1_G3_MINI_ALU_ix468 (.Y (L1_4_L2_1_G3_MINI_ALU_nx467), .A0 (
          nx6576), .A1 (L1_4_L2_1_G3_MINI_ALU_BoothP_9), .S0 (
          L1_4_L2_1_G3_MINI_ALU_nx463)) ;
    inv01 ix6575 (.Y (nx6576), .A (L1_4_L2_1_G3_MINI_ALU_nx461)) ;
    mux21 L1_4_L2_1_G3_MINI_ALU_ix476 (.Y (L1_4_L2_1_G3_MINI_ALU_nx475), .A0 (
          nx6578), .A1 (L1_4_L2_1_G3_MINI_ALU_BoothP_10), .S0 (
          L1_4_L2_1_G3_MINI_ALU_nx471)) ;
    inv01 ix6577 (.Y (nx6578), .A (L1_4_L2_1_G3_MINI_ALU_nx467)) ;
    mux21 L1_4_L2_1_G3_MINI_ALU_ix484 (.Y (L1_4_L2_1_G3_MINI_ALU_nx483), .A0 (
          nx6580), .A1 (L1_4_L2_1_G3_MINI_ALU_BoothP_11), .S0 (
          L1_4_L2_1_G3_MINI_ALU_nx479)) ;
    inv01 ix6579 (.Y (nx6580), .A (L1_4_L2_1_G3_MINI_ALU_nx475)) ;
    mux21 L1_4_L2_1_G3_MINI_ALU_ix492 (.Y (L1_4_L2_1_G3_MINI_ALU_nx491), .A0 (
          nx6582), .A1 (L1_4_L2_1_G3_MINI_ALU_BoothP_12), .S0 (
          L1_4_L2_1_G3_MINI_ALU_nx487)) ;
    inv01 ix6581 (.Y (nx6582), .A (L1_4_L2_1_G3_MINI_ALU_nx483)) ;
    mux21 L1_4_L2_1_G3_MINI_ALU_ix500 (.Y (L1_4_L2_1_G3_MINI_ALU_nx499), .A0 (
          nx6584), .A1 (L1_4_L2_1_G3_MINI_ALU_BoothP_13), .S0 (
          L1_4_L2_1_G3_MINI_ALU_nx495)) ;
    inv01 ix6583 (.Y (nx6584), .A (L1_4_L2_1_G3_MINI_ALU_nx491)) ;
    mux21 L1_4_L2_1_G3_MINI_ALU_ix508 (.Y (L1_4_L2_1_G3_MINI_ALU_nx507), .A0 (
          nx6586), .A1 (L1_4_L2_1_G3_MINI_ALU_BoothP_14), .S0 (
          L1_4_L2_1_G3_MINI_ALU_nx503)) ;
    inv01 ix6585 (.Y (nx6586), .A (L1_4_L2_1_G3_MINI_ALU_nx499)) ;
    mux21 L1_4_L2_1_G3_MINI_ALU_ix516 (.Y (L1_4_L2_1_G3_MINI_ALU_nx515), .A0 (
          nx6588), .A1 (L1_4_L2_1_G3_MINI_ALU_BoothP_15), .S0 (
          L1_4_L2_1_G3_MINI_ALU_nx511)) ;
    inv01 ix6587 (.Y (nx6588), .A (L1_4_L2_1_G3_MINI_ALU_nx507)) ;
    mux21 L1_4_L2_1_G3_MINI_ALU_ix161 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_1), .A0 (nx6590), .A1 (
          L1_4_L2_1_G3_MINI_ALU_nx379), .S0 (nx8438)) ;
    inv01 ix6589 (.Y (nx6590), .A (L1_4_L2_1_G3_MINI_ALU_BoothP_1)) ;
    mux21 L1_4_L2_1_G3_MINI_ALU_ix181 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_2), .A0 (
          L1_4_L2_1_G3_MINI_ALU_nx387), .A1 (L1_4_L2_1_G3_MINI_ALU_nx389), .S0 (
          nx8438)) ;
    mux21 L1_4_L2_1_G3_MINI_ALU_ix201 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_3), .A0 (
          L1_4_L2_1_G3_MINI_ALU_nx399), .A1 (L1_4_L2_1_G3_MINI_ALU_nx401), .S0 (
          nx8438)) ;
    mux21 L1_4_L2_1_G3_MINI_ALU_ix221 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_4), .A0 (
          L1_4_L2_1_G3_MINI_ALU_nx409), .A1 (L1_4_L2_1_G3_MINI_ALU_nx411), .S0 (
          nx8438)) ;
    mux21 L1_4_L2_1_G3_MINI_ALU_ix241 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_5), .A0 (
          L1_4_L2_1_G3_MINI_ALU_nx419), .A1 (L1_4_L2_1_G3_MINI_ALU_nx421), .S0 (
          nx8438)) ;
    mux21 L1_4_L2_1_G3_MINI_ALU_ix261 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_6), .A0 (
          L1_4_L2_1_G3_MINI_ALU_nx429), .A1 (L1_4_L2_1_G3_MINI_ALU_nx431), .S0 (
          nx8438)) ;
    mux21 L1_4_L2_1_G3_MINI_ALU_ix281 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_7), .A0 (
          L1_4_L2_1_G3_MINI_ALU_nx439), .A1 (L1_4_L2_1_G3_MINI_ALU_nx441), .S0 (
          nx8438)) ;
    mux21 L1_4_L2_1_G3_MINI_ALU_ix301 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_8), .A0 (
          L1_4_L2_1_G3_MINI_ALU_nx449), .A1 (L1_4_L2_1_G3_MINI_ALU_nx451), .S0 (
          nx8440)) ;
    mux21 L1_4_L2_1_G3_MINI_ALU_ix321 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_9), .A0 (
          L1_4_L2_1_G3_MINI_ALU_nx469), .A1 (nx6592), .S0 (nx8440)) ;
    inv01 ix6591 (.Y (nx6592), .A (L1_4_L2_1_G3_MINI_ALU_nx316)) ;
    mux21 L1_4_L2_1_G3_MINI_ALU_ix341 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_10), .A0 (
          L1_4_L2_1_G3_MINI_ALU_nx477), .A1 (nx6594), .S0 (nx8440)) ;
    inv01 ix6593 (.Y (nx6594), .A (L1_4_L2_1_G3_MINI_ALU_nx336)) ;
    mux21 L1_4_L2_1_G3_MINI_ALU_ix361 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_11), .A0 (
          L1_4_L2_1_G3_MINI_ALU_nx485), .A1 (nx6596), .S0 (nx8440)) ;
    inv01 ix6595 (.Y (nx6596), .A (L1_4_L2_1_G3_MINI_ALU_nx356)) ;
    mux21 L1_4_L2_1_G3_MINI_ALU_ix381 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_12), .A0 (
          L1_4_L2_1_G3_MINI_ALU_nx493), .A1 (nx6598), .S0 (nx8440)) ;
    inv01 ix6597 (.Y (nx6598), .A (L1_4_L2_1_G3_MINI_ALU_nx376)) ;
    mux21 L1_4_L2_1_G3_MINI_ALU_ix401 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_13), .A0 (
          L1_4_L2_1_G3_MINI_ALU_nx501), .A1 (nx6600), .S0 (nx8440)) ;
    inv01 ix6599 (.Y (nx6600), .A (L1_4_L2_1_G3_MINI_ALU_nx396)) ;
    mux21 L1_4_L2_1_G3_MINI_ALU_ix421 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_14), .A0 (
          L1_4_L2_1_G3_MINI_ALU_nx509), .A1 (nx6602), .S0 (nx8440)) ;
    inv01 ix6601 (.Y (nx6602), .A (L1_4_L2_1_G3_MINI_ALU_nx416)) ;
    mux21 L1_4_L2_1_G3_MINI_ALU_ix441 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_15), .A0 (
          L1_4_L2_1_G3_MINI_ALU_nx517), .A1 (nx6604), .S0 (nx8442)) ;
    inv01 ix6603 (.Y (nx6604), .A (L1_4_L2_1_G3_MINI_ALU_nx436)) ;
    mux21 L1_4_L2_1_G3_MINI_ALU_ix461 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_16), .A0 (nx6606), .A1 (nx6608
          ), .S0 (nx8442)) ;
    inv01 ix6605 (.Y (nx6606), .A (L1_4_L2_1_G3_MINI_ALU_BoothP_16)) ;
    inv01 ix6607 (.Y (nx6608), .A (L1_4_L2_1_G3_MINI_ALU_nx456)) ;
    nor02_2x L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix319 (.Y (
             L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642), .A0 (Start), .A1 (
             CalculatingBooth_dup_1253)) ;
    nor02_2x L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix85 (.Y (
             L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_0), .A0 (nx8452), .A1 (
             nx6610)) ;
    inv01 ix6609 (.Y (nx6610), .A (L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_1)) ;
    mux21 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix125 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_1), .A0 (nx6612), .A1 (
          nx6614), .S0 (nx8452)) ;
    inv01 ix6611 (.Y (nx6612), .A (L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_2)) ;
    inv01 ix6613 (.Y (nx6614), .A (WindowDin_4__1__0)) ;
    mux21 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix133 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_2), .A0 (nx6616), .A1 (
          nx6618), .S0 (nx8452)) ;
    inv01 ix6615 (.Y (nx6616), .A (L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_3)) ;
    inv01 ix6617 (.Y (nx6618), .A (WindowDin_4__1__1)) ;
    mux21 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix141 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_3), .A0 (nx6620), .A1 (
          nx6622), .S0 (nx8452)) ;
    inv01 ix6619 (.Y (nx6620), .A (L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_4)) ;
    inv01 ix6621 (.Y (nx6622), .A (WindowDin_4__1__2)) ;
    mux21 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix149 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_4), .A0 (nx6624), .A1 (
          nx6626), .S0 (nx8452)) ;
    inv01 ix6623 (.Y (nx6624), .A (L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_5)) ;
    inv01 ix6625 (.Y (nx6626), .A (WindowDin_4__1__3)) ;
    mux21 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix157 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_5), .A0 (nx6628), .A1 (
          nx6630), .S0 (nx8452)) ;
    inv01 ix6627 (.Y (nx6628), .A (L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_6)) ;
    inv01 ix6629 (.Y (nx6630), .A (WindowDin_4__1__4)) ;
    mux21 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix165 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_6), .A0 (nx6632), .A1 (
          nx6634), .S0 (nx8452)) ;
    inv01 ix6631 (.Y (nx6632), .A (L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_7)) ;
    inv01 ix6633 (.Y (nx6634), .A (WindowDin_4__1__5)) ;
    mux21 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix173 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_7), .A0 (nx6636), .A1 (
          nx6638), .S0 (nx8454)) ;
    inv01 ix6635 (.Y (nx6636), .A (L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_8)) ;
    inv01 ix6637 (.Y (nx6638), .A (WindowDin_4__1__6)) ;
    mux21 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix181 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_8), .A0 (nx6640), .A1 (
          nx6642), .S0 (nx8454)) ;
    inv01 ix6639 (.Y (nx6640), .A (L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_9)) ;
    inv01 ix6641 (.Y (nx6642), .A (WindowDin_4__1__7)) ;
    nor02_2x L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix89 (.Y (
             L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_9), .A0 (nx8454), .A1 (
             nx6644)) ;
    inv01 ix6643 (.Y (nx6644), .A (L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_10)
          ) ;
    nor02_2x L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix93 (.Y (
             L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_10), .A0 (nx8454), .A1 (
             nx6646)) ;
    inv01 ix6645 (.Y (nx6646), .A (L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_11)
          ) ;
    nor02_2x L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix97 (.Y (
             L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_11), .A0 (nx8454), .A1 (
             nx6648)) ;
    inv01 ix6647 (.Y (nx6648), .A (L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_12)
          ) ;
    nor02_2x L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix101 (.Y (
             L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_12), .A0 (nx8454), .A1 (
             nx6650)) ;
    inv01 ix6649 (.Y (nx6650), .A (L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_13)
          ) ;
    nor02_2x L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix105 (.Y (
             L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_13), .A0 (nx8454), .A1 (
             nx6652)) ;
    inv01 ix6651 (.Y (nx6652), .A (L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_14)
          ) ;
    nor02_2x L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix109 (.Y (
             L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_14), .A0 (nx8456), .A1 (
             nx6654)) ;
    inv01 ix6653 (.Y (nx6654), .A (L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_15)
          ) ;
    nor02_2x L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix113 (.Y (
             L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_15), .A0 (nx8456), .A1 (
             nx6656)) ;
    inv01 ix6655 (.Y (nx6656), .A (L1_4_L2_1_G3_MINI_ALU_BoothPBeforeShift_16)
          ) ;
    nor02_2x L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix117 (.Y (
             L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_16), .A0 (nx8456), .A1 (
             nx6656)) ;
    mux21 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix189 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BoothOperand_0), .A0 (nx6658), .A1 (nx6660), .S0 (
          nx8444)) ;
    inv01 ix6657 (.Y (nx6658), .A (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_0)) ;
    inv01 ix6659 (.Y (nx6660), .A (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_0)) ;
    mux21 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix197 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BoothOperand_1), .A0 (nx6662), .A1 (nx6664), .S0 (
          nx8444)) ;
    inv01 ix6661 (.Y (nx6662), .A (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_1)) ;
    inv01 ix6663 (.Y (nx6664), .A (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_1)) ;
    mux21 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix205 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BoothOperand_2), .A0 (nx6666), .A1 (nx6668), .S0 (
          nx8444)) ;
    inv01 ix6665 (.Y (nx6666), .A (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_2)) ;
    inv01 ix6667 (.Y (nx6668), .A (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_2)) ;
    mux21 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix213 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BoothOperand_3), .A0 (nx6670), .A1 (nx6672), .S0 (
          nx8444)) ;
    inv01 ix6669 (.Y (nx6670), .A (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_3)) ;
    inv01 ix6671 (.Y (nx6672), .A (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_3)) ;
    mux21 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix221 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BoothOperand_4), .A0 (nx6674), .A1 (nx6676), .S0 (
          nx8444)) ;
    inv01 ix6673 (.Y (nx6674), .A (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_4)) ;
    inv01 ix6675 (.Y (nx6676), .A (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_4)) ;
    mux21 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix229 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BoothOperand_5), .A0 (nx6678), .A1 (nx6680), .S0 (
          nx8446)) ;
    inv01 ix6677 (.Y (nx6678), .A (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_5)) ;
    inv01 ix6679 (.Y (nx6680), .A (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_5)) ;
    mux21 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix237 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BoothOperand_6), .A0 (nx6682), .A1 (nx6684), .S0 (
          nx8446)) ;
    inv01 ix6681 (.Y (nx6682), .A (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_6)) ;
    inv01 ix6683 (.Y (nx6684), .A (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_6)) ;
    mux21 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix245 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BoothOperand_7), .A0 (nx6686), .A1 (nx6688), .S0 (
          nx8446)) ;
    inv01 ix6685 (.Y (nx6686), .A (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_7)) ;
    inv01 ix6687 (.Y (nx6688), .A (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_7)) ;
    mux21 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix253 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BoothOperand_8), .A0 (nx6690), .A1 (nx6692), .S0 (
          nx8446)) ;
    inv01 ix6689 (.Y (nx6690), .A (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_8)) ;
    inv01 ix6691 (.Y (nx6692), .A (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_8)) ;
    mux21 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix261 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BoothOperand_9), .A0 (nx6694), .A1 (nx6696), .S0 (
          nx8446)) ;
    inv01 ix6693 (.Y (nx6694), .A (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_9)) ;
    inv01 ix6695 (.Y (nx6696), .A (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_9)) ;
    mux21 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix269 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BoothOperand_10), .A0 (nx6698), .A1 (nx6700), .S0 (
          nx8446)) ;
    inv01 ix6697 (.Y (nx6698), .A (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_10)) ;
    inv01 ix6699 (.Y (nx6700), .A (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_10)) ;
    mux21 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix277 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BoothOperand_11), .A0 (nx6702), .A1 (nx6704), .S0 (
          nx8446)) ;
    inv01 ix6701 (.Y (nx6702), .A (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_11)) ;
    inv01 ix6703 (.Y (nx6704), .A (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_11)) ;
    mux21 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix285 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BoothOperand_12), .A0 (nx6706), .A1 (nx6708), .S0 (
          nx8448)) ;
    inv01 ix6705 (.Y (nx6706), .A (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_12)) ;
    inv01 ix6707 (.Y (nx6708), .A (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_12)) ;
    mux21 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix293 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BoothOperand_13), .A0 (nx6710), .A1 (nx6712), .S0 (
          nx8448)) ;
    inv01 ix6709 (.Y (nx6710), .A (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_13)) ;
    inv01 ix6711 (.Y (nx6712), .A (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_13)) ;
    mux21 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix301 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BoothOperand_14), .A0 (nx6714), .A1 (nx6716), .S0 (
          nx8448)) ;
    inv01 ix6713 (.Y (nx6714), .A (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_14)) ;
    inv01 ix6715 (.Y (nx6716), .A (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_14)) ;
    mux21 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix309 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BoothOperand_15), .A0 (nx6718), .A1 (nx6720), .S0 (
          nx8448)) ;
    inv01 ix6717 (.Y (nx6718), .A (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_15)) ;
    inv01 ix6719 (.Y (nx6720), .A (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_15)) ;
    mux21 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix317 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BoothOperand_16), .A0 (nx6722), .A1 (nx6724), .S0 (
          nx8448)) ;
    inv01 ix6721 (.Y (nx6722), .A (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDout_16)) ;
    inv01 ix6723 (.Y (nx6724), .A (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterADout_16)) ;
    xnor2 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_ix321 (.Y (
          L1_4_L2_1_G3_MINI_ALU_AddPToBoothOperand), .A0 (nx8448), .A1 (nx6590)
          ) ;
    oai32 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix393 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .A0 (nx8722), .A1 (
          RST), .A2 (nx8458), .B0 (nx6660), .B1 (nx6728)) ;
    oai32 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix403 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .A0 (nx8722), .A1 (
          RST), .A2 (nx8458), .B0 (nx6664), .B1 (nx6728)) ;
    oai32 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix413 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .A0 (nx8722), .A1 (
          RST), .A2 (nx8458), .B0 (nx6668), .B1 (nx6728)) ;
    oai32 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix423 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .A0 (nx8722), .A1 (
          RST), .A2 (nx8458), .B0 (nx6672), .B1 (nx6728)) ;
    oai32 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix433 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .A0 (nx8722), .A1 (
          RST), .A2 (nx8458), .B0 (nx6676), .B1 (nx6728)) ;
    oai32 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix443 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .A0 (nx8722), .A1 (
          RST), .A2 (nx8458), .B0 (nx6680), .B1 (nx6728)) ;
    oai32 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix453 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .A0 (nx8722), .A1 (
          RST), .A2 (nx8460), .B0 (nx6684), .B1 (nx6728)) ;
    oai32 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix463 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .A0 (nx8724), .A1 (
          RST), .A2 (nx8460), .B0 (nx6688), .B1 (nx6730)) ;
    oai32 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix473 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .A0 (nx8724), .A1 (
          RST), .A2 (nx8460), .B0 (nx6692), .B1 (nx6730)) ;
    oai32 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix483 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .A0 (nx6732), .A1 (
          RST), .A2 (nx8460), .B0 (nx6696), .B1 (nx6730)) ;
    inv01 ix6731 (.Y (nx6732), .A (FilterDin_4__1__0)) ;
    oai32 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix493 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .A0 (nx6734), .A1 (
          RST), .A2 (nx8460), .B0 (nx6700), .B1 (nx6730)) ;
    inv01 ix6733 (.Y (nx6734), .A (FilterDin_4__1__1)) ;
    oai32 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix503 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .A0 (nx6736), .A1 (
          RST), .A2 (nx8460), .B0 (nx6704), .B1 (nx6730)) ;
    inv01 ix6735 (.Y (nx6736), .A (FilterDin_4__1__2)) ;
    oai32 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix513 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .A0 (nx6738), .A1 (
          RST), .A2 (nx8460), .B0 (nx6708), .B1 (nx6730)) ;
    inv01 ix6737 (.Y (nx6738), .A (FilterDin_4__1__3)) ;
    oai32 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix523 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .A0 (nx6740), .A1 (
          RST), .A2 (nx8462), .B0 (nx6712), .B1 (nx6730)) ;
    inv01 ix6739 (.Y (nx6740), .A (FilterDin_4__1__4)) ;
    oai32 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix533 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .A0 (nx6742), .A1 (
          RST), .A2 (nx8462), .B0 (nx6716), .B1 (nx6744)) ;
    inv01 ix6741 (.Y (nx6742), .A (FilterDin_4__1__5)) ;
    inv01 ix6743 (.Y (nx6744), .A (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566)) ;
    oai32 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix543 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .A0 (nx6746), .A1 (
          RST), .A2 (nx8462), .B0 (nx6720), .B1 (nx6744)) ;
    inv01 ix6745 (.Y (nx6746), .A (FilterDin_4__1__6)) ;
    oai32 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix553 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .A0 (nx6748), .A1 (
          RST), .A2 (nx8462), .B0 (nx6724), .B1 (nx6744)) ;
    inv01 ix6747 (.Y (nx6748), .A (FilterDin_4__1__7)) ;
    nand02_2x L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix633 (.Y (nx6728), .A0 (
              nx7612), .A1 (nx8462)) ;
    nand02_2x L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix635 (.Y (nx6730), .A0 (
              nx7612), .A1 (nx8462)) ;
    oai32 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix393 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .A0 (nx8724), .A1 (
          RST), .A2 (nx8464), .B0 (nx6658), .B1 (nx6750)) ;
    oai32 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix403 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .A0 (nx8724), .A1 (
          RST), .A2 (nx8464), .B0 (nx6662), .B1 (nx6750)) ;
    oai32 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix413 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .A0 (nx8724), .A1 (
          RST), .A2 (nx8464), .B0 (nx6666), .B1 (nx6750)) ;
    oai32 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix423 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .A0 (nx8724), .A1 (
          RST), .A2 (nx8464), .B0 (nx6670), .B1 (nx6750)) ;
    oai32 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix433 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .A0 (nx8724), .A1 (
          RST), .A2 (nx8464), .B0 (nx6674), .B1 (nx6750)) ;
    oai32 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix443 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .A0 (nx8726), .A1 (
          RST), .A2 (nx8464), .B0 (nx6678), .B1 (nx6750)) ;
    oai32 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix453 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .A0 (nx8726), .A1 (
          RST), .A2 (nx8466), .B0 (nx6682), .B1 (nx6750)) ;
    oai32 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix463 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .A0 (nx8726), .A1 (
          RST), .A2 (nx8466), .B0 (nx6686), .B1 (nx6752)) ;
    oai32 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix473 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .A0 (nx8726), .A1 (
          RST), .A2 (nx8466), .B0 (nx6690), .B1 (nx6752)) ;
    oai32 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix483 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .A0 (nx6732), .A1 (
          RST), .A2 (nx8466), .B0 (nx6694), .B1 (nx6752)) ;
    oai32 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix493 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .A0 (nx6754), .A1 (
          RST), .A2 (nx8466), .B0 (nx6698), .B1 (nx6752)) ;
    inv01 ix6753 (.Y (nx6754), .A (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_10)) ;
    oai32 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix503 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .A0 (nx6756), .A1 (
          RST), .A2 (nx8466), .B0 (nx6702), .B1 (nx6752)) ;
    inv01 ix6755 (.Y (nx6756), .A (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_11)) ;
    oai32 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix513 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .A0 (nx6758), .A1 (
          RST), .A2 (nx8466), .B0 (nx6706), .B1 (nx6752)) ;
    inv01 ix6757 (.Y (nx6758), .A (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_12)) ;
    oai32 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix523 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .A0 (nx6760), .A1 (
          RST), .A2 (nx8468), .B0 (nx6710), .B1 (nx6752)) ;
    inv01 ix6759 (.Y (nx6760), .A (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_13)) ;
    oai32 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix533 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .A0 (nx6762), .A1 (
          RST), .A2 (nx8468), .B0 (nx6714), .B1 (nx6764)) ;
    inv01 ix6761 (.Y (nx6762), .A (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_14)) ;
    inv01 ix6763 (.Y (nx6764), .A (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566)) ;
    oai32 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix543 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .A0 (nx6766), .A1 (
          RST), .A2 (nx8468), .B0 (nx6718), .B1 (nx6764)) ;
    inv01 ix6765 (.Y (nx6766), .A (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_15)) ;
    oai32 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix553 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .A0 (nx6768), .A1 (
          RST), .A2 (nx8468), .B0 (nx6722), .B1 (nx6764)) ;
    inv01 ix6767 (.Y (nx6768), .A (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterSDin_16)) ;
    nand02_2x L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix633 (.Y (nx6750), .A0 (
              nx7612), .A1 (nx8468)) ;
    nand02_2x L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix635 (.Y (nx6752), .A0 (
              nx7612), .A1 (nx8468)) ;
    oai32 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix393 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .A0 (nx6770), .A1 (
          RST), .A2 (nx8470), .B0 (L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_nx384), .B1 (
          nx6772)) ;
    inv01 ix6769 (.Y (nx6770), .A (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_0)) ;
    oai32 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix403 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .A0 (nx6774), .A1 (
          RST), .A2 (nx8470), .B0 (nx6590), .B1 (nx6772)) ;
    inv01 ix6773 (.Y (nx6774), .A (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_1)) ;
    oai32 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix413 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .A0 (nx6776), .A1 (
          RST), .A2 (nx8470), .B0 (L1_4_L2_1_G3_MINI_ALU_nx387), .B1 (nx6772)) ;
    inv01 ix6775 (.Y (nx6776), .A (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_2)) ;
    oai32 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix423 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .A0 (nx6778), .A1 (
          RST), .A2 (nx8470), .B0 (L1_4_L2_1_G3_MINI_ALU_nx399), .B1 (nx6772)) ;
    inv01 ix6777 (.Y (nx6778), .A (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_3)) ;
    oai32 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix433 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .A0 (nx6780), .A1 (
          RST), .A2 (nx8470), .B0 (L1_4_L2_1_G3_MINI_ALU_nx409), .B1 (nx6772)) ;
    inv01 ix6779 (.Y (nx6780), .A (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_4)) ;
    oai32 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix443 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .A0 (nx6782), .A1 (
          RST), .A2 (nx8470), .B0 (L1_4_L2_1_G3_MINI_ALU_nx419), .B1 (nx6772)) ;
    inv01 ix6781 (.Y (nx6782), .A (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_5)) ;
    oai32 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix453 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .A0 (nx6784), .A1 (
          RST), .A2 (nx8470), .B0 (L1_4_L2_1_G3_MINI_ALU_nx429), .B1 (nx6772)) ;
    inv01 ix6783 (.Y (nx6784), .A (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_6)) ;
    oai32 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix463 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .A0 (nx6786), .A1 (
          RST), .A2 (nx8472), .B0 (L1_4_L2_1_G3_MINI_ALU_nx439), .B1 (nx6788)) ;
    inv01 ix6785 (.Y (nx6786), .A (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_7)) ;
    oai32 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix473 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .A0 (nx6790), .A1 (
          RST), .A2 (nx8472), .B0 (L1_4_L2_1_G3_MINI_ALU_nx449), .B1 (nx6788)) ;
    inv01 ix6789 (.Y (nx6790), .A (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_8)) ;
    oai32 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix483 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .A0 (nx6792), .A1 (
          RST), .A2 (nx8472), .B0 (L1_4_L2_1_G3_MINI_ALU_nx469), .B1 (nx6788)) ;
    inv01 ix6791 (.Y (nx6792), .A (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_9)) ;
    oai32 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix493 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .A0 (nx6794), .A1 (
          RST), .A2 (nx8472), .B0 (L1_4_L2_1_G3_MINI_ALU_nx477), .B1 (nx6788)) ;
    inv01 ix6793 (.Y (nx6794), .A (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_10)) ;
    oai32 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix503 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .A0 (nx6796), .A1 (
          RST), .A2 (nx8472), .B0 (L1_4_L2_1_G3_MINI_ALU_nx485), .B1 (nx6788)) ;
    inv01 ix6795 (.Y (nx6796), .A (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_11)) ;
    oai32 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix513 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .A0 (nx6798), .A1 (
          RST), .A2 (nx8472), .B0 (L1_4_L2_1_G3_MINI_ALU_nx493), .B1 (nx6788)) ;
    inv01 ix6797 (.Y (nx6798), .A (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_12)) ;
    oai32 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix523 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .A0 (nx6800), .A1 (
          RST), .A2 (nx8472), .B0 (L1_4_L2_1_G3_MINI_ALU_nx501), .B1 (nx6788)) ;
    inv01 ix6799 (.Y (nx6800), .A (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_13)) ;
    oai32 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix533 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .A0 (nx6802), .A1 (
          RST), .A2 (nx8474), .B0 (L1_4_L2_1_G3_MINI_ALU_nx509), .B1 (nx6804)) ;
    inv01 ix6801 (.Y (nx6802), .A (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_14)) ;
    inv01 ix6803 (.Y (nx6804), .A (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566)) ;
    oai32 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix543 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .A0 (nx6806), .A1 (
          RST), .A2 (nx8474), .B0 (L1_4_L2_1_G3_MINI_ALU_nx517), .B1 (nx6804)) ;
    inv01 ix6805 (.Y (nx6806), .A (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_15)) ;
    oai32 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix553 (.Y (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .A0 (nx6808), .A1 (
          RST), .A2 (nx8474), .B0 (nx6606), .B1 (nx6804)) ;
    inv01 ix6807 (.Y (nx6808), .A (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_RegisterPDin_16)) ;
    nand02_2x L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix633 (.Y (nx6772), .A0 (
              nx7612), .A1 (nx8474)) ;
    nand02_2x L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix635 (.Y (nx6788), .A0 (
              nx7612), .A1 (nx8474)) ;
    mux21 L1_4_L2_2_G4_MINI_ALU_ix404 (.Y (L1_4_L2_2_G4_MINI_ALU_nx403), .A0 (
          nx6810), .A1 (L1_4_L2_2_G4_MINI_ALU_BoothP_2), .S0 (
          L1_4_L2_2_G4_MINI_ALU_nx395)) ;
    inv01 ix6809 (.Y (nx6810), .A (L1_4_L2_2_G4_MINI_ALU_nx391)) ;
    mux21 L1_4_L2_2_G4_MINI_ALU_ix414 (.Y (L1_4_L2_2_G4_MINI_ALU_nx413), .A0 (
          nx6812), .A1 (L1_4_L2_2_G4_MINI_ALU_BoothP_3), .S0 (
          L1_4_L2_2_G4_MINI_ALU_nx405)) ;
    inv01 ix6811 (.Y (nx6812), .A (L1_4_L2_2_G4_MINI_ALU_nx403)) ;
    mux21 L1_4_L2_2_G4_MINI_ALU_ix424 (.Y (L1_4_L2_2_G4_MINI_ALU_nx423), .A0 (
          nx6814), .A1 (L1_4_L2_2_G4_MINI_ALU_BoothP_4), .S0 (
          L1_4_L2_2_G4_MINI_ALU_nx415)) ;
    inv01 ix6813 (.Y (nx6814), .A (L1_4_L2_2_G4_MINI_ALU_nx413)) ;
    mux21 L1_4_L2_2_G4_MINI_ALU_ix434 (.Y (L1_4_L2_2_G4_MINI_ALU_nx433), .A0 (
          nx6816), .A1 (L1_4_L2_2_G4_MINI_ALU_BoothP_5), .S0 (
          L1_4_L2_2_G4_MINI_ALU_nx425)) ;
    inv01 ix6815 (.Y (nx6816), .A (L1_4_L2_2_G4_MINI_ALU_nx423)) ;
    mux21 L1_4_L2_2_G4_MINI_ALU_ix444 (.Y (L1_4_L2_2_G4_MINI_ALU_nx443), .A0 (
          nx6818), .A1 (L1_4_L2_2_G4_MINI_ALU_BoothP_6), .S0 (
          L1_4_L2_2_G4_MINI_ALU_nx435)) ;
    inv01 ix6817 (.Y (nx6818), .A (L1_4_L2_2_G4_MINI_ALU_nx433)) ;
    mux21 L1_4_L2_2_G4_MINI_ALU_ix454 (.Y (L1_4_L2_2_G4_MINI_ALU_nx453), .A0 (
          nx6820), .A1 (L1_4_L2_2_G4_MINI_ALU_BoothP_7), .S0 (
          L1_4_L2_2_G4_MINI_ALU_nx445)) ;
    inv01 ix6819 (.Y (nx6820), .A (L1_4_L2_2_G4_MINI_ALU_nx443)) ;
    mux21 L1_4_L2_2_G4_MINI_ALU_ix462 (.Y (L1_4_L2_2_G4_MINI_ALU_nx461), .A0 (
          nx6822), .A1 (L1_4_L2_2_G4_MINI_ALU_BoothP_8), .S0 (
          L1_4_L2_2_G4_MINI_ALU_nx455)) ;
    inv01 ix6821 (.Y (nx6822), .A (L1_4_L2_2_G4_MINI_ALU_nx453)) ;
    mux21 L1_4_L2_2_G4_MINI_ALU_ix468 (.Y (L1_4_L2_2_G4_MINI_ALU_nx467), .A0 (
          nx6824), .A1 (L1_4_L2_2_G4_MINI_ALU_BoothP_9), .S0 (
          L1_4_L2_2_G4_MINI_ALU_nx463)) ;
    inv01 ix6823 (.Y (nx6824), .A (L1_4_L2_2_G4_MINI_ALU_nx461)) ;
    mux21 L1_4_L2_2_G4_MINI_ALU_ix476 (.Y (L1_4_L2_2_G4_MINI_ALU_nx475), .A0 (
          nx6826), .A1 (L1_4_L2_2_G4_MINI_ALU_BoothP_10), .S0 (
          L1_4_L2_2_G4_MINI_ALU_nx471)) ;
    inv01 ix6825 (.Y (nx6826), .A (L1_4_L2_2_G4_MINI_ALU_nx467)) ;
    mux21 L1_4_L2_2_G4_MINI_ALU_ix484 (.Y (L1_4_L2_2_G4_MINI_ALU_nx483), .A0 (
          nx6828), .A1 (L1_4_L2_2_G4_MINI_ALU_BoothP_11), .S0 (
          L1_4_L2_2_G4_MINI_ALU_nx479)) ;
    inv01 ix6827 (.Y (nx6828), .A (L1_4_L2_2_G4_MINI_ALU_nx475)) ;
    mux21 L1_4_L2_2_G4_MINI_ALU_ix492 (.Y (L1_4_L2_2_G4_MINI_ALU_nx491), .A0 (
          nx6830), .A1 (L1_4_L2_2_G4_MINI_ALU_BoothP_12), .S0 (
          L1_4_L2_2_G4_MINI_ALU_nx487)) ;
    inv01 ix6829 (.Y (nx6830), .A (L1_4_L2_2_G4_MINI_ALU_nx483)) ;
    mux21 L1_4_L2_2_G4_MINI_ALU_ix500 (.Y (L1_4_L2_2_G4_MINI_ALU_nx499), .A0 (
          nx6832), .A1 (L1_4_L2_2_G4_MINI_ALU_BoothP_13), .S0 (
          L1_4_L2_2_G4_MINI_ALU_nx495)) ;
    inv01 ix6831 (.Y (nx6832), .A (L1_4_L2_2_G4_MINI_ALU_nx491)) ;
    mux21 L1_4_L2_2_G4_MINI_ALU_ix508 (.Y (L1_4_L2_2_G4_MINI_ALU_nx507), .A0 (
          nx6834), .A1 (L1_4_L2_2_G4_MINI_ALU_BoothP_14), .S0 (
          L1_4_L2_2_G4_MINI_ALU_nx503)) ;
    inv01 ix6833 (.Y (nx6834), .A (L1_4_L2_2_G4_MINI_ALU_nx499)) ;
    mux21 L1_4_L2_2_G4_MINI_ALU_ix516 (.Y (L1_4_L2_2_G4_MINI_ALU_nx515), .A0 (
          nx6836), .A1 (L1_4_L2_2_G4_MINI_ALU_BoothP_15), .S0 (
          L1_4_L2_2_G4_MINI_ALU_nx511)) ;
    inv01 ix6835 (.Y (nx6836), .A (L1_4_L2_2_G4_MINI_ALU_nx507)) ;
    mux21 L1_4_L2_2_G4_MINI_ALU_ix161 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_1), .A0 (nx6838), .A1 (
          L1_4_L2_2_G4_MINI_ALU_nx379), .S0 (nx8478)) ;
    inv01 ix6837 (.Y (nx6838), .A (L1_4_L2_2_G4_MINI_ALU_BoothP_1)) ;
    mux21 L1_4_L2_2_G4_MINI_ALU_ix181 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_2), .A0 (
          L1_4_L2_2_G4_MINI_ALU_nx387), .A1 (L1_4_L2_2_G4_MINI_ALU_nx389), .S0 (
          nx8478)) ;
    mux21 L1_4_L2_2_G4_MINI_ALU_ix201 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_3), .A0 (
          L1_4_L2_2_G4_MINI_ALU_nx399), .A1 (L1_4_L2_2_G4_MINI_ALU_nx401), .S0 (
          nx8478)) ;
    mux21 L1_4_L2_2_G4_MINI_ALU_ix221 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_4), .A0 (
          L1_4_L2_2_G4_MINI_ALU_nx409), .A1 (L1_4_L2_2_G4_MINI_ALU_nx411), .S0 (
          nx8478)) ;
    mux21 L1_4_L2_2_G4_MINI_ALU_ix241 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_5), .A0 (
          L1_4_L2_2_G4_MINI_ALU_nx419), .A1 (L1_4_L2_2_G4_MINI_ALU_nx421), .S0 (
          nx8478)) ;
    mux21 L1_4_L2_2_G4_MINI_ALU_ix261 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_6), .A0 (
          L1_4_L2_2_G4_MINI_ALU_nx429), .A1 (L1_4_L2_2_G4_MINI_ALU_nx431), .S0 (
          nx8478)) ;
    mux21 L1_4_L2_2_G4_MINI_ALU_ix281 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_7), .A0 (
          L1_4_L2_2_G4_MINI_ALU_nx439), .A1 (L1_4_L2_2_G4_MINI_ALU_nx441), .S0 (
          nx8478)) ;
    mux21 L1_4_L2_2_G4_MINI_ALU_ix301 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_8), .A0 (
          L1_4_L2_2_G4_MINI_ALU_nx449), .A1 (L1_4_L2_2_G4_MINI_ALU_nx451), .S0 (
          nx8480)) ;
    mux21 L1_4_L2_2_G4_MINI_ALU_ix321 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_9), .A0 (
          L1_4_L2_2_G4_MINI_ALU_nx469), .A1 (nx6840), .S0 (nx8480)) ;
    inv01 ix6839 (.Y (nx6840), .A (L1_4_L2_2_G4_MINI_ALU_nx316)) ;
    mux21 L1_4_L2_2_G4_MINI_ALU_ix341 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_10), .A0 (
          L1_4_L2_2_G4_MINI_ALU_nx477), .A1 (nx6842), .S0 (nx8480)) ;
    inv01 ix6841 (.Y (nx6842), .A (L1_4_L2_2_G4_MINI_ALU_nx336)) ;
    mux21 L1_4_L2_2_G4_MINI_ALU_ix361 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_11), .A0 (
          L1_4_L2_2_G4_MINI_ALU_nx485), .A1 (nx6844), .S0 (nx8480)) ;
    inv01 ix6843 (.Y (nx6844), .A (L1_4_L2_2_G4_MINI_ALU_nx356)) ;
    mux21 L1_4_L2_2_G4_MINI_ALU_ix381 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_12), .A0 (
          L1_4_L2_2_G4_MINI_ALU_nx493), .A1 (nx6846), .S0 (nx8480)) ;
    inv01 ix6845 (.Y (nx6846), .A (L1_4_L2_2_G4_MINI_ALU_nx376)) ;
    mux21 L1_4_L2_2_G4_MINI_ALU_ix401 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_13), .A0 (
          L1_4_L2_2_G4_MINI_ALU_nx501), .A1 (nx6848), .S0 (nx8480)) ;
    inv01 ix6847 (.Y (nx6848), .A (L1_4_L2_2_G4_MINI_ALU_nx396)) ;
    mux21 L1_4_L2_2_G4_MINI_ALU_ix421 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_14), .A0 (
          L1_4_L2_2_G4_MINI_ALU_nx509), .A1 (nx6850), .S0 (nx8480)) ;
    inv01 ix6849 (.Y (nx6850), .A (L1_4_L2_2_G4_MINI_ALU_nx416)) ;
    mux21 L1_4_L2_2_G4_MINI_ALU_ix441 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_15), .A0 (
          L1_4_L2_2_G4_MINI_ALU_nx517), .A1 (nx6852), .S0 (nx8482)) ;
    inv01 ix6851 (.Y (nx6852), .A (L1_4_L2_2_G4_MINI_ALU_nx436)) ;
    mux21 L1_4_L2_2_G4_MINI_ALU_ix461 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_16), .A0 (nx6854), .A1 (nx6856
          ), .S0 (nx8482)) ;
    inv01 ix6853 (.Y (nx6854), .A (L1_4_L2_2_G4_MINI_ALU_BoothP_16)) ;
    inv01 ix6855 (.Y (nx6856), .A (L1_4_L2_2_G4_MINI_ALU_nx456)) ;
    nor02_2x L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix319 (.Y (
             L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642), .A0 (Start), .A1 (
             CalculatingBooth_dup_1253)) ;
    nor02_2x L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix85 (.Y (
             L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_0), .A0 (nx8492), .A1 (
             nx6858)) ;
    inv01 ix6857 (.Y (nx6858), .A (L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_1)) ;
    mux21 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix125 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_1), .A0 (nx6860), .A1 (
          nx6862), .S0 (nx8492)) ;
    inv01 ix6859 (.Y (nx6860), .A (L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_2)) ;
    inv01 ix6861 (.Y (nx6862), .A (WindowDin_4__2__0)) ;
    mux21 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix133 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_2), .A0 (nx6864), .A1 (
          nx6866), .S0 (nx8492)) ;
    inv01 ix6863 (.Y (nx6864), .A (L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_3)) ;
    inv01 ix6865 (.Y (nx6866), .A (WindowDin_4__2__1)) ;
    mux21 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix141 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_3), .A0 (nx6868), .A1 (
          nx6870), .S0 (nx8492)) ;
    inv01 ix6867 (.Y (nx6868), .A (L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_4)) ;
    inv01 ix6869 (.Y (nx6870), .A (WindowDin_4__2__2)) ;
    mux21 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix149 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_4), .A0 (nx6872), .A1 (
          nx6874), .S0 (nx8492)) ;
    inv01 ix6871 (.Y (nx6872), .A (L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_5)) ;
    inv01 ix6873 (.Y (nx6874), .A (WindowDin_4__2__3)) ;
    mux21 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix157 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_5), .A0 (nx6876), .A1 (
          nx6878), .S0 (nx8492)) ;
    inv01 ix6875 (.Y (nx6876), .A (L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_6)) ;
    inv01 ix6877 (.Y (nx6878), .A (WindowDin_4__2__4)) ;
    mux21 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix165 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_6), .A0 (nx6880), .A1 (
          nx6882), .S0 (nx8492)) ;
    inv01 ix6879 (.Y (nx6880), .A (L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_7)) ;
    inv01 ix6881 (.Y (nx6882), .A (WindowDin_4__2__5)) ;
    mux21 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix173 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_7), .A0 (nx6884), .A1 (
          nx6886), .S0 (nx8494)) ;
    inv01 ix6883 (.Y (nx6884), .A (L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_8)) ;
    inv01 ix6885 (.Y (nx6886), .A (WindowDin_4__2__6)) ;
    mux21 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix181 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_8), .A0 (nx6888), .A1 (
          nx6890), .S0 (nx8494)) ;
    inv01 ix6887 (.Y (nx6888), .A (L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_9)) ;
    inv01 ix6889 (.Y (nx6890), .A (WindowDin_4__2__7)) ;
    nor02_2x L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix89 (.Y (
             L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_9), .A0 (nx8494), .A1 (
             nx6892)) ;
    inv01 ix6891 (.Y (nx6892), .A (L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_10)
          ) ;
    nor02_2x L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix93 (.Y (
             L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_10), .A0 (nx8494), .A1 (
             nx6894)) ;
    inv01 ix6893 (.Y (nx6894), .A (L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_11)
          ) ;
    nor02_2x L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix97 (.Y (
             L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_11), .A0 (nx8494), .A1 (
             nx6896)) ;
    inv01 ix6895 (.Y (nx6896), .A (L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_12)
          ) ;
    nor02_2x L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix101 (.Y (
             L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_12), .A0 (nx8494), .A1 (
             nx6898)) ;
    inv01 ix6897 (.Y (nx6898), .A (L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_13)
          ) ;
    nor02_2x L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix105 (.Y (
             L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_13), .A0 (nx8494), .A1 (
             nx6900)) ;
    inv01 ix6899 (.Y (nx6900), .A (L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_14)
          ) ;
    nor02_2x L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix109 (.Y (
             L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_14), .A0 (nx8496), .A1 (
             nx6902)) ;
    inv01 ix6901 (.Y (nx6902), .A (L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_15)
          ) ;
    nor02_2x L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix113 (.Y (
             L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_15), .A0 (nx8496), .A1 (
             nx6904)) ;
    inv01 ix6903 (.Y (nx6904), .A (L1_4_L2_2_G4_MINI_ALU_BoothPBeforeShift_16)
          ) ;
    nor02_2x L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix117 (.Y (
             L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_16), .A0 (nx8496), .A1 (
             nx6904)) ;
    mux21 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix189 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BoothOperand_0), .A0 (nx6906), .A1 (nx6908), .S0 (
          nx8484)) ;
    inv01 ix6905 (.Y (nx6906), .A (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_0)) ;
    inv01 ix6907 (.Y (nx6908), .A (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_0)) ;
    mux21 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix197 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BoothOperand_1), .A0 (nx6910), .A1 (nx6912), .S0 (
          nx8484)) ;
    inv01 ix6909 (.Y (nx6910), .A (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_1)) ;
    inv01 ix6911 (.Y (nx6912), .A (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_1)) ;
    mux21 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix205 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BoothOperand_2), .A0 (nx6914), .A1 (nx6916), .S0 (
          nx8484)) ;
    inv01 ix6913 (.Y (nx6914), .A (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_2)) ;
    inv01 ix6915 (.Y (nx6916), .A (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_2)) ;
    mux21 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix213 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BoothOperand_3), .A0 (nx6918), .A1 (nx6920), .S0 (
          nx8484)) ;
    inv01 ix6917 (.Y (nx6918), .A (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_3)) ;
    inv01 ix6919 (.Y (nx6920), .A (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_3)) ;
    mux21 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix221 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BoothOperand_4), .A0 (nx6922), .A1 (nx6924), .S0 (
          nx8484)) ;
    inv01 ix6921 (.Y (nx6922), .A (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_4)) ;
    inv01 ix6923 (.Y (nx6924), .A (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_4)) ;
    mux21 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix229 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BoothOperand_5), .A0 (nx6926), .A1 (nx6928), .S0 (
          nx8486)) ;
    inv01 ix6925 (.Y (nx6926), .A (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_5)) ;
    inv01 ix6927 (.Y (nx6928), .A (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_5)) ;
    mux21 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix237 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BoothOperand_6), .A0 (nx6930), .A1 (nx6932), .S0 (
          nx8486)) ;
    inv01 ix6929 (.Y (nx6930), .A (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_6)) ;
    inv01 ix6931 (.Y (nx6932), .A (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_6)) ;
    mux21 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix245 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BoothOperand_7), .A0 (nx6934), .A1 (nx6936), .S0 (
          nx8486)) ;
    inv01 ix6933 (.Y (nx6934), .A (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_7)) ;
    inv01 ix6935 (.Y (nx6936), .A (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_7)) ;
    mux21 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix253 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BoothOperand_8), .A0 (nx6938), .A1 (nx6940), .S0 (
          nx8486)) ;
    inv01 ix6937 (.Y (nx6938), .A (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_8)) ;
    inv01 ix6939 (.Y (nx6940), .A (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_8)) ;
    mux21 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix261 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BoothOperand_9), .A0 (nx6942), .A1 (nx6944), .S0 (
          nx8486)) ;
    inv01 ix6941 (.Y (nx6942), .A (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_9)) ;
    inv01 ix6943 (.Y (nx6944), .A (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_9)) ;
    mux21 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix269 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BoothOperand_10), .A0 (nx6946), .A1 (nx6948), .S0 (
          nx8486)) ;
    inv01 ix6945 (.Y (nx6946), .A (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_10)) ;
    inv01 ix6947 (.Y (nx6948), .A (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_10)) ;
    mux21 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix277 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BoothOperand_11), .A0 (nx6950), .A1 (nx6952), .S0 (
          nx8486)) ;
    inv01 ix6949 (.Y (nx6950), .A (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_11)) ;
    inv01 ix6951 (.Y (nx6952), .A (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_11)) ;
    mux21 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix285 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BoothOperand_12), .A0 (nx6954), .A1 (nx6956), .S0 (
          nx8488)) ;
    inv01 ix6953 (.Y (nx6954), .A (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_12)) ;
    inv01 ix6955 (.Y (nx6956), .A (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_12)) ;
    mux21 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix293 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BoothOperand_13), .A0 (nx6958), .A1 (nx6960), .S0 (
          nx8488)) ;
    inv01 ix6957 (.Y (nx6958), .A (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_13)) ;
    inv01 ix6959 (.Y (nx6960), .A (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_13)) ;
    mux21 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix301 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BoothOperand_14), .A0 (nx6962), .A1 (nx6964), .S0 (
          nx8488)) ;
    inv01 ix6961 (.Y (nx6962), .A (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_14)) ;
    inv01 ix6963 (.Y (nx6964), .A (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_14)) ;
    mux21 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix309 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BoothOperand_15), .A0 (nx6966), .A1 (nx6968), .S0 (
          nx8488)) ;
    inv01 ix6965 (.Y (nx6966), .A (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_15)) ;
    inv01 ix6967 (.Y (nx6968), .A (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_15)) ;
    mux21 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix317 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BoothOperand_16), .A0 (nx6970), .A1 (nx6972), .S0 (
          nx8488)) ;
    inv01 ix6969 (.Y (nx6970), .A (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDout_16)) ;
    inv01 ix6971 (.Y (nx6972), .A (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterADout_16)) ;
    xnor2 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_ix321 (.Y (
          L1_4_L2_2_G4_MINI_ALU_AddPToBoothOperand), .A0 (nx8488), .A1 (nx6838)
          ) ;
    oai32 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix393 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .A0 (nx8728), .A1 (
          RST), .A2 (nx8498), .B0 (nx6908), .B1 (nx6976)) ;
    oai32 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix403 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .A0 (nx8728), .A1 (
          RST), .A2 (nx8498), .B0 (nx6912), .B1 (nx6976)) ;
    oai32 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix413 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .A0 (nx8728), .A1 (
          RST), .A2 (nx8498), .B0 (nx6916), .B1 (nx6976)) ;
    oai32 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix423 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .A0 (nx8728), .A1 (
          RST), .A2 (nx8498), .B0 (nx6920), .B1 (nx6976)) ;
    oai32 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix433 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .A0 (nx8728), .A1 (
          RST), .A2 (nx8498), .B0 (nx6924), .B1 (nx6976)) ;
    oai32 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix443 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .A0 (nx8728), .A1 (
          RST), .A2 (nx8498), .B0 (nx6928), .B1 (nx6976)) ;
    oai32 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix453 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .A0 (nx8728), .A1 (
          RST), .A2 (nx8500), .B0 (nx6932), .B1 (nx6976)) ;
    oai32 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix463 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .A0 (nx8730), .A1 (
          RST), .A2 (nx8500), .B0 (nx6936), .B1 (nx6978)) ;
    oai32 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix473 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .A0 (nx8730), .A1 (
          RST), .A2 (nx8500), .B0 (nx6940), .B1 (nx6978)) ;
    oai32 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix483 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .A0 (nx6980), .A1 (
          RST), .A2 (nx8500), .B0 (nx6944), .B1 (nx6978)) ;
    inv01 ix6979 (.Y (nx6980), .A (FilterDin_4__2__0)) ;
    oai32 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix493 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .A0 (nx6982), .A1 (
          RST), .A2 (nx8500), .B0 (nx6948), .B1 (nx6978)) ;
    inv01 ix6981 (.Y (nx6982), .A (FilterDin_4__2__1)) ;
    oai32 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix503 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .A0 (nx6984), .A1 (
          RST), .A2 (nx8500), .B0 (nx6952), .B1 (nx6978)) ;
    inv01 ix6983 (.Y (nx6984), .A (FilterDin_4__2__2)) ;
    oai32 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix513 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .A0 (nx6986), .A1 (
          RST), .A2 (nx8500), .B0 (nx6956), .B1 (nx6978)) ;
    inv01 ix6985 (.Y (nx6986), .A (FilterDin_4__2__3)) ;
    oai32 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix523 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .A0 (nx6988), .A1 (
          RST), .A2 (nx8502), .B0 (nx6960), .B1 (nx6978)) ;
    inv01 ix6987 (.Y (nx6988), .A (FilterDin_4__2__4)) ;
    oai32 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix533 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .A0 (nx6990), .A1 (
          RST), .A2 (nx8502), .B0 (nx6964), .B1 (nx6992)) ;
    inv01 ix6989 (.Y (nx6990), .A (FilterDin_4__2__5)) ;
    inv01 ix6991 (.Y (nx6992), .A (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566)) ;
    oai32 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix543 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .A0 (nx6994), .A1 (
          RST), .A2 (nx8502), .B0 (nx6968), .B1 (nx6992)) ;
    inv01 ix6993 (.Y (nx6994), .A (FilterDin_4__2__6)) ;
    oai32 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix553 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .A0 (nx6996), .A1 (
          RST), .A2 (nx8502), .B0 (nx6972), .B1 (nx6992)) ;
    inv01 ix6995 (.Y (nx6996), .A (FilterDin_4__2__7)) ;
    nand02_2x L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix633 (.Y (nx6976), .A0 (
              nx7612), .A1 (nx8502)) ;
    nand02_2x L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix635 (.Y (nx6978), .A0 (
              nx7614), .A1 (nx8502)) ;
    oai32 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix393 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .A0 (nx8730), .A1 (
          RST), .A2 (nx8504), .B0 (nx6906), .B1 (nx6998)) ;
    oai32 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix403 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .A0 (nx8730), .A1 (
          RST), .A2 (nx8504), .B0 (nx6910), .B1 (nx6998)) ;
    oai32 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix413 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .A0 (nx8730), .A1 (
          RST), .A2 (nx8504), .B0 (nx6914), .B1 (nx6998)) ;
    oai32 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix423 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .A0 (nx8730), .A1 (
          RST), .A2 (nx8504), .B0 (nx6918), .B1 (nx6998)) ;
    oai32 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix433 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .A0 (nx8730), .A1 (
          RST), .A2 (nx8504), .B0 (nx6922), .B1 (nx6998)) ;
    oai32 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix443 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .A0 (nx8732), .A1 (
          RST), .A2 (nx8504), .B0 (nx6926), .B1 (nx6998)) ;
    oai32 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix453 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .A0 (nx8732), .A1 (
          RST), .A2 (nx8506), .B0 (nx6930), .B1 (nx6998)) ;
    oai32 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix463 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .A0 (nx8732), .A1 (
          RST), .A2 (nx8506), .B0 (nx6934), .B1 (nx7000)) ;
    oai32 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix473 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .A0 (nx8732), .A1 (
          RST), .A2 (nx8506), .B0 (nx6938), .B1 (nx7000)) ;
    oai32 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix483 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .A0 (nx6980), .A1 (
          RST), .A2 (nx8506), .B0 (nx6942), .B1 (nx7000)) ;
    oai32 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix493 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .A0 (nx7002), .A1 (
          RST), .A2 (nx8506), .B0 (nx6946), .B1 (nx7000)) ;
    inv01 ix7001 (.Y (nx7002), .A (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDin_10)) ;
    oai32 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix503 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .A0 (nx7004), .A1 (
          RST), .A2 (nx8506), .B0 (nx6950), .B1 (nx7000)) ;
    inv01 ix7003 (.Y (nx7004), .A (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDin_11)) ;
    oai32 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix513 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .A0 (nx7006), .A1 (
          RST), .A2 (nx8506), .B0 (nx6954), .B1 (nx7000)) ;
    inv01 ix7005 (.Y (nx7006), .A (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDin_12)) ;
    oai32 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix523 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .A0 (nx7008), .A1 (
          RST), .A2 (nx8508), .B0 (nx6958), .B1 (nx7000)) ;
    inv01 ix7007 (.Y (nx7008), .A (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDin_13)) ;
    oai32 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix533 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .A0 (nx7010), .A1 (
          RST), .A2 (nx8508), .B0 (nx6962), .B1 (nx7012)) ;
    inv01 ix7009 (.Y (nx7010), .A (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDin_14)) ;
    inv01 ix7011 (.Y (nx7012), .A (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566)) ;
    oai32 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix543 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .A0 (nx7014), .A1 (
          RST), .A2 (nx8508), .B0 (nx6966), .B1 (nx7012)) ;
    inv01 ix7013 (.Y (nx7014), .A (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDin_15)) ;
    oai32 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix553 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .A0 (nx7016), .A1 (
          RST), .A2 (nx8508), .B0 (nx6970), .B1 (nx7012)) ;
    inv01 ix7015 (.Y (nx7016), .A (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterSDin_16)) ;
    nand02_2x L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix633 (.Y (nx6998), .A0 (
              nx7614), .A1 (nx8508)) ;
    nand02_2x L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix635 (.Y (nx7000), .A0 (
              nx7614), .A1 (nx8508)) ;
    oai32 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix393 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .A0 (nx7018), .A1 (
          RST), .A2 (nx8510), .B0 (L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_nx384), .B1 (
          nx7020)) ;
    inv01 ix7017 (.Y (nx7018), .A (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_0)) ;
    oai32 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix403 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .A0 (nx7022), .A1 (
          RST), .A2 (nx8510), .B0 (nx6838), .B1 (nx7020)) ;
    inv01 ix7021 (.Y (nx7022), .A (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_1)) ;
    oai32 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix413 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .A0 (nx7024), .A1 (
          RST), .A2 (nx8510), .B0 (L1_4_L2_2_G4_MINI_ALU_nx387), .B1 (nx7020)) ;
    inv01 ix7023 (.Y (nx7024), .A (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_2)) ;
    oai32 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix423 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .A0 (nx7026), .A1 (
          RST), .A2 (nx8510), .B0 (L1_4_L2_2_G4_MINI_ALU_nx399), .B1 (nx7020)) ;
    inv01 ix7025 (.Y (nx7026), .A (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_3)) ;
    oai32 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix433 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .A0 (nx7028), .A1 (
          RST), .A2 (nx8510), .B0 (L1_4_L2_2_G4_MINI_ALU_nx409), .B1 (nx7020)) ;
    inv01 ix7027 (.Y (nx7028), .A (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_4)) ;
    oai32 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix443 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .A0 (nx7030), .A1 (
          RST), .A2 (nx8510), .B0 (L1_4_L2_2_G4_MINI_ALU_nx419), .B1 (nx7020)) ;
    inv01 ix7029 (.Y (nx7030), .A (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_5)) ;
    oai32 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix453 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .A0 (nx7032), .A1 (
          RST), .A2 (nx8510), .B0 (L1_4_L2_2_G4_MINI_ALU_nx429), .B1 (nx7020)) ;
    inv01 ix7031 (.Y (nx7032), .A (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_6)) ;
    oai32 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix463 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .A0 (nx7034), .A1 (
          RST), .A2 (nx8512), .B0 (L1_4_L2_2_G4_MINI_ALU_nx439), .B1 (nx7036)) ;
    inv01 ix7033 (.Y (nx7034), .A (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_7)) ;
    oai32 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix473 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .A0 (nx7038), .A1 (
          RST), .A2 (nx8512), .B0 (L1_4_L2_2_G4_MINI_ALU_nx449), .B1 (nx7036)) ;
    inv01 ix7037 (.Y (nx7038), .A (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_8)) ;
    oai32 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix483 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .A0 (nx7040), .A1 (
          RST), .A2 (nx8512), .B0 (L1_4_L2_2_G4_MINI_ALU_nx469), .B1 (nx7036)) ;
    inv01 ix7039 (.Y (nx7040), .A (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_9)) ;
    oai32 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix493 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .A0 (nx7042), .A1 (
          RST), .A2 (nx8512), .B0 (L1_4_L2_2_G4_MINI_ALU_nx477), .B1 (nx7036)) ;
    inv01 ix7041 (.Y (nx7042), .A (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_10)) ;
    oai32 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix503 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .A0 (nx7044), .A1 (
          RST), .A2 (nx8512), .B0 (L1_4_L2_2_G4_MINI_ALU_nx485), .B1 (nx7036)) ;
    inv01 ix7043 (.Y (nx7044), .A (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_11)) ;
    oai32 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix513 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .A0 (nx7046), .A1 (
          RST), .A2 (nx8512), .B0 (L1_4_L2_2_G4_MINI_ALU_nx493), .B1 (nx7036)) ;
    inv01 ix7045 (.Y (nx7046), .A (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_12)) ;
    oai32 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix523 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .A0 (nx7048), .A1 (
          RST), .A2 (nx8512), .B0 (L1_4_L2_2_G4_MINI_ALU_nx501), .B1 (nx7036)) ;
    inv01 ix7047 (.Y (nx7048), .A (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_13)) ;
    oai32 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix533 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .A0 (nx7050), .A1 (
          RST), .A2 (nx8514), .B0 (L1_4_L2_2_G4_MINI_ALU_nx509), .B1 (nx7052)) ;
    inv01 ix7049 (.Y (nx7050), .A (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_14)) ;
    inv01 ix7051 (.Y (nx7052), .A (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566)) ;
    oai32 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix543 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .A0 (nx7054), .A1 (
          RST), .A2 (nx8514), .B0 (L1_4_L2_2_G4_MINI_ALU_nx517), .B1 (nx7052)) ;
    inv01 ix7053 (.Y (nx7054), .A (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_15)) ;
    oai32 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix553 (.Y (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .A0 (nx7056), .A1 (
          RST), .A2 (nx8514), .B0 (nx6854), .B1 (nx7052)) ;
    inv01 ix7055 (.Y (nx7056), .A (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_RegisterPDin_16)) ;
    nand02_2x L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix633 (.Y (nx7020), .A0 (
              nx7614), .A1 (nx8514)) ;
    nand02_2x L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix635 (.Y (nx7036), .A0 (
              nx7614), .A1 (nx8514)) ;
    mux21 L1_4_L2_3_G5_MINI_ALU_ix404 (.Y (L1_4_L2_3_G5_MINI_ALU_nx403), .A0 (
          nx7058), .A1 (L1_4_L2_3_G5_MINI_ALU_BoothP_2), .S0 (
          L1_4_L2_3_G5_MINI_ALU_nx395)) ;
    inv01 ix7057 (.Y (nx7058), .A (L1_4_L2_3_G5_MINI_ALU_nx391)) ;
    mux21 L1_4_L2_3_G5_MINI_ALU_ix414 (.Y (L1_4_L2_3_G5_MINI_ALU_nx413), .A0 (
          nx7060), .A1 (L1_4_L2_3_G5_MINI_ALU_BoothP_3), .S0 (
          L1_4_L2_3_G5_MINI_ALU_nx405)) ;
    inv01 ix7059 (.Y (nx7060), .A (L1_4_L2_3_G5_MINI_ALU_nx403)) ;
    mux21 L1_4_L2_3_G5_MINI_ALU_ix424 (.Y (L1_4_L2_3_G5_MINI_ALU_nx423), .A0 (
          nx7062), .A1 (L1_4_L2_3_G5_MINI_ALU_BoothP_4), .S0 (
          L1_4_L2_3_G5_MINI_ALU_nx415)) ;
    inv01 ix7061 (.Y (nx7062), .A (L1_4_L2_3_G5_MINI_ALU_nx413)) ;
    mux21 L1_4_L2_3_G5_MINI_ALU_ix434 (.Y (L1_4_L2_3_G5_MINI_ALU_nx433), .A0 (
          nx7064), .A1 (L1_4_L2_3_G5_MINI_ALU_BoothP_5), .S0 (
          L1_4_L2_3_G5_MINI_ALU_nx425)) ;
    inv01 ix7063 (.Y (nx7064), .A (L1_4_L2_3_G5_MINI_ALU_nx423)) ;
    mux21 L1_4_L2_3_G5_MINI_ALU_ix444 (.Y (L1_4_L2_3_G5_MINI_ALU_nx443), .A0 (
          nx7066), .A1 (L1_4_L2_3_G5_MINI_ALU_BoothP_6), .S0 (
          L1_4_L2_3_G5_MINI_ALU_nx435)) ;
    inv01 ix7065 (.Y (nx7066), .A (L1_4_L2_3_G5_MINI_ALU_nx433)) ;
    mux21 L1_4_L2_3_G5_MINI_ALU_ix454 (.Y (L1_4_L2_3_G5_MINI_ALU_nx453), .A0 (
          nx7068), .A1 (L1_4_L2_3_G5_MINI_ALU_BoothP_7), .S0 (
          L1_4_L2_3_G5_MINI_ALU_nx445)) ;
    inv01 ix7067 (.Y (nx7068), .A (L1_4_L2_3_G5_MINI_ALU_nx443)) ;
    mux21 L1_4_L2_3_G5_MINI_ALU_ix462 (.Y (L1_4_L2_3_G5_MINI_ALU_nx461), .A0 (
          nx7070), .A1 (L1_4_L2_3_G5_MINI_ALU_BoothP_8), .S0 (
          L1_4_L2_3_G5_MINI_ALU_nx455)) ;
    inv01 ix7069 (.Y (nx7070), .A (L1_4_L2_3_G5_MINI_ALU_nx453)) ;
    mux21 L1_4_L2_3_G5_MINI_ALU_ix468 (.Y (L1_4_L2_3_G5_MINI_ALU_nx467), .A0 (
          nx7072), .A1 (L1_4_L2_3_G5_MINI_ALU_BoothP_9), .S0 (
          L1_4_L2_3_G5_MINI_ALU_nx463)) ;
    inv01 ix7071 (.Y (nx7072), .A (L1_4_L2_3_G5_MINI_ALU_nx461)) ;
    mux21 L1_4_L2_3_G5_MINI_ALU_ix476 (.Y (L1_4_L2_3_G5_MINI_ALU_nx475), .A0 (
          nx7074), .A1 (L1_4_L2_3_G5_MINI_ALU_BoothP_10), .S0 (
          L1_4_L2_3_G5_MINI_ALU_nx471)) ;
    inv01 ix7073 (.Y (nx7074), .A (L1_4_L2_3_G5_MINI_ALU_nx467)) ;
    mux21 L1_4_L2_3_G5_MINI_ALU_ix484 (.Y (L1_4_L2_3_G5_MINI_ALU_nx483), .A0 (
          nx7076), .A1 (L1_4_L2_3_G5_MINI_ALU_BoothP_11), .S0 (
          L1_4_L2_3_G5_MINI_ALU_nx479)) ;
    inv01 ix7075 (.Y (nx7076), .A (L1_4_L2_3_G5_MINI_ALU_nx475)) ;
    mux21 L1_4_L2_3_G5_MINI_ALU_ix492 (.Y (L1_4_L2_3_G5_MINI_ALU_nx491), .A0 (
          nx7078), .A1 (L1_4_L2_3_G5_MINI_ALU_BoothP_12), .S0 (
          L1_4_L2_3_G5_MINI_ALU_nx487)) ;
    inv01 ix7077 (.Y (nx7078), .A (L1_4_L2_3_G5_MINI_ALU_nx483)) ;
    mux21 L1_4_L2_3_G5_MINI_ALU_ix500 (.Y (L1_4_L2_3_G5_MINI_ALU_nx499), .A0 (
          nx7080), .A1 (L1_4_L2_3_G5_MINI_ALU_BoothP_13), .S0 (
          L1_4_L2_3_G5_MINI_ALU_nx495)) ;
    inv01 ix7079 (.Y (nx7080), .A (L1_4_L2_3_G5_MINI_ALU_nx491)) ;
    mux21 L1_4_L2_3_G5_MINI_ALU_ix508 (.Y (L1_4_L2_3_G5_MINI_ALU_nx507), .A0 (
          nx7082), .A1 (L1_4_L2_3_G5_MINI_ALU_BoothP_14), .S0 (
          L1_4_L2_3_G5_MINI_ALU_nx503)) ;
    inv01 ix7081 (.Y (nx7082), .A (L1_4_L2_3_G5_MINI_ALU_nx499)) ;
    mux21 L1_4_L2_3_G5_MINI_ALU_ix516 (.Y (L1_4_L2_3_G5_MINI_ALU_nx515), .A0 (
          nx7084), .A1 (L1_4_L2_3_G5_MINI_ALU_BoothP_15), .S0 (
          L1_4_L2_3_G5_MINI_ALU_nx511)) ;
    inv01 ix7083 (.Y (nx7084), .A (L1_4_L2_3_G5_MINI_ALU_nx507)) ;
    mux21 L1_4_L2_3_G5_MINI_ALU_ix161 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_1), .A0 (nx7086), .A1 (
          L1_4_L2_3_G5_MINI_ALU_nx379), .S0 (nx8518)) ;
    inv01 ix7085 (.Y (nx7086), .A (L1_4_L2_3_G5_MINI_ALU_BoothP_1)) ;
    mux21 L1_4_L2_3_G5_MINI_ALU_ix181 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_2), .A0 (
          L1_4_L2_3_G5_MINI_ALU_nx387), .A1 (L1_4_L2_3_G5_MINI_ALU_nx389), .S0 (
          nx8518)) ;
    mux21 L1_4_L2_3_G5_MINI_ALU_ix201 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_3), .A0 (
          L1_4_L2_3_G5_MINI_ALU_nx399), .A1 (L1_4_L2_3_G5_MINI_ALU_nx401), .S0 (
          nx8518)) ;
    mux21 L1_4_L2_3_G5_MINI_ALU_ix221 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_4), .A0 (
          L1_4_L2_3_G5_MINI_ALU_nx409), .A1 (L1_4_L2_3_G5_MINI_ALU_nx411), .S0 (
          nx8518)) ;
    mux21 L1_4_L2_3_G5_MINI_ALU_ix241 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_5), .A0 (
          L1_4_L2_3_G5_MINI_ALU_nx419), .A1 (L1_4_L2_3_G5_MINI_ALU_nx421), .S0 (
          nx8518)) ;
    mux21 L1_4_L2_3_G5_MINI_ALU_ix261 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_6), .A0 (
          L1_4_L2_3_G5_MINI_ALU_nx429), .A1 (L1_4_L2_3_G5_MINI_ALU_nx431), .S0 (
          nx8518)) ;
    mux21 L1_4_L2_3_G5_MINI_ALU_ix281 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_7), .A0 (
          L1_4_L2_3_G5_MINI_ALU_nx439), .A1 (L1_4_L2_3_G5_MINI_ALU_nx441), .S0 (
          nx8518)) ;
    mux21 L1_4_L2_3_G5_MINI_ALU_ix301 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_8), .A0 (
          L1_4_L2_3_G5_MINI_ALU_nx449), .A1 (L1_4_L2_3_G5_MINI_ALU_nx451), .S0 (
          nx8520)) ;
    mux21 L1_4_L2_3_G5_MINI_ALU_ix321 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_9), .A0 (
          L1_4_L2_3_G5_MINI_ALU_nx469), .A1 (nx7088), .S0 (nx8520)) ;
    inv01 ix7087 (.Y (nx7088), .A (L1_4_L2_3_G5_MINI_ALU_nx316)) ;
    mux21 L1_4_L2_3_G5_MINI_ALU_ix341 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_10), .A0 (
          L1_4_L2_3_G5_MINI_ALU_nx477), .A1 (nx7090), .S0 (nx8520)) ;
    inv01 ix7089 (.Y (nx7090), .A (L1_4_L2_3_G5_MINI_ALU_nx336)) ;
    mux21 L1_4_L2_3_G5_MINI_ALU_ix361 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_11), .A0 (
          L1_4_L2_3_G5_MINI_ALU_nx485), .A1 (nx7092), .S0 (nx8520)) ;
    inv01 ix7091 (.Y (nx7092), .A (L1_4_L2_3_G5_MINI_ALU_nx356)) ;
    mux21 L1_4_L2_3_G5_MINI_ALU_ix381 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_12), .A0 (
          L1_4_L2_3_G5_MINI_ALU_nx493), .A1 (nx7094), .S0 (nx8520)) ;
    inv01 ix7093 (.Y (nx7094), .A (L1_4_L2_3_G5_MINI_ALU_nx376)) ;
    mux21 L1_4_L2_3_G5_MINI_ALU_ix401 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_13), .A0 (
          L1_4_L2_3_G5_MINI_ALU_nx501), .A1 (nx7096), .S0 (nx8520)) ;
    inv01 ix7095 (.Y (nx7096), .A (L1_4_L2_3_G5_MINI_ALU_nx396)) ;
    mux21 L1_4_L2_3_G5_MINI_ALU_ix421 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_14), .A0 (
          L1_4_L2_3_G5_MINI_ALU_nx509), .A1 (nx7098), .S0 (nx8520)) ;
    inv01 ix7097 (.Y (nx7098), .A (L1_4_L2_3_G5_MINI_ALU_nx416)) ;
    mux21 L1_4_L2_3_G5_MINI_ALU_ix441 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_15), .A0 (
          L1_4_L2_3_G5_MINI_ALU_nx517), .A1 (nx7100), .S0 (nx8522)) ;
    inv01 ix7099 (.Y (nx7100), .A (L1_4_L2_3_G5_MINI_ALU_nx436)) ;
    mux21 L1_4_L2_3_G5_MINI_ALU_ix461 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_16), .A0 (nx7102), .A1 (nx7104
          ), .S0 (nx8522)) ;
    inv01 ix7101 (.Y (nx7102), .A (L1_4_L2_3_G5_MINI_ALU_BoothP_16)) ;
    inv01 ix7103 (.Y (nx7104), .A (L1_4_L2_3_G5_MINI_ALU_nx456)) ;
    nor02_2x L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix319 (.Y (
             L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642), .A0 (Start), .A1 (
             CalculatingBooth_dup_1253)) ;
    nor02_2x L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix85 (.Y (
             L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_0), .A0 (nx8532), .A1 (
             nx7106)) ;
    inv01 ix7105 (.Y (nx7106), .A (L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_1)) ;
    mux21 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix125 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_1), .A0 (nx7108), .A1 (
          nx7110), .S0 (nx8532)) ;
    inv01 ix7107 (.Y (nx7108), .A (L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_2)) ;
    inv01 ix7109 (.Y (nx7110), .A (WindowDin_4__3__0)) ;
    mux21 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix133 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_2), .A0 (nx7112), .A1 (
          nx7114), .S0 (nx8532)) ;
    inv01 ix7111 (.Y (nx7112), .A (L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_3)) ;
    inv01 ix7113 (.Y (nx7114), .A (WindowDin_4__3__1)) ;
    mux21 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix141 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_3), .A0 (nx7116), .A1 (
          nx7118), .S0 (nx8532)) ;
    inv01 ix7115 (.Y (nx7116), .A (L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_4)) ;
    inv01 ix7117 (.Y (nx7118), .A (WindowDin_4__3__2)) ;
    mux21 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix149 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_4), .A0 (nx7120), .A1 (
          nx7122), .S0 (nx8532)) ;
    inv01 ix7119 (.Y (nx7120), .A (L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_5)) ;
    inv01 ix7121 (.Y (nx7122), .A (WindowDin_4__3__3)) ;
    mux21 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix157 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_5), .A0 (nx7124), .A1 (
          nx7126), .S0 (nx8532)) ;
    inv01 ix7123 (.Y (nx7124), .A (L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_6)) ;
    inv01 ix7125 (.Y (nx7126), .A (WindowDin_4__3__4)) ;
    mux21 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix165 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_6), .A0 (nx7128), .A1 (
          nx7130), .S0 (nx8532)) ;
    inv01 ix7127 (.Y (nx7128), .A (L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_7)) ;
    inv01 ix7129 (.Y (nx7130), .A (WindowDin_4__3__5)) ;
    mux21 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix173 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_7), .A0 (nx7132), .A1 (
          nx7134), .S0 (nx8534)) ;
    inv01 ix7131 (.Y (nx7132), .A (L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_8)) ;
    inv01 ix7133 (.Y (nx7134), .A (WindowDin_4__3__6)) ;
    mux21 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix181 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_8), .A0 (nx7136), .A1 (
          nx7138), .S0 (nx8534)) ;
    inv01 ix7135 (.Y (nx7136), .A (L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_9)) ;
    inv01 ix7137 (.Y (nx7138), .A (WindowDin_4__3__7)) ;
    nor02_2x L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix89 (.Y (
             L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_9), .A0 (nx8534), .A1 (
             nx7140)) ;
    inv01 ix7139 (.Y (nx7140), .A (L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_10)
          ) ;
    nor02_2x L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix93 (.Y (
             L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_10), .A0 (nx8534), .A1 (
             nx7142)) ;
    inv01 ix7141 (.Y (nx7142), .A (L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_11)
          ) ;
    nor02_2x L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix97 (.Y (
             L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_11), .A0 (nx8534), .A1 (
             nx7144)) ;
    inv01 ix7143 (.Y (nx7144), .A (L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_12)
          ) ;
    nor02_2x L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix101 (.Y (
             L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_12), .A0 (nx8534), .A1 (
             nx7146)) ;
    inv01 ix7145 (.Y (nx7146), .A (L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_13)
          ) ;
    nor02_2x L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix105 (.Y (
             L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_13), .A0 (nx8534), .A1 (
             nx7148)) ;
    inv01 ix7147 (.Y (nx7148), .A (L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_14)
          ) ;
    nor02_2x L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix109 (.Y (
             L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_14), .A0 (nx8536), .A1 (
             nx7150)) ;
    inv01 ix7149 (.Y (nx7150), .A (L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_15)
          ) ;
    nor02_2x L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix113 (.Y (
             L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_15), .A0 (nx8536), .A1 (
             nx7152)) ;
    inv01 ix7151 (.Y (nx7152), .A (L1_4_L2_3_G5_MINI_ALU_BoothPBeforeShift_16)
          ) ;
    nor02_2x L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix117 (.Y (
             L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_16), .A0 (nx8536), .A1 (
             nx7152)) ;
    mux21 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix189 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BoothOperand_0), .A0 (nx7154), .A1 (nx7156), .S0 (
          nx8524)) ;
    inv01 ix7153 (.Y (nx7154), .A (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_0)) ;
    inv01 ix7155 (.Y (nx7156), .A (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_0)) ;
    mux21 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix197 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BoothOperand_1), .A0 (nx7158), .A1 (nx7160), .S0 (
          nx8524)) ;
    inv01 ix7157 (.Y (nx7158), .A (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_1)) ;
    inv01 ix7159 (.Y (nx7160), .A (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_1)) ;
    mux21 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix205 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BoothOperand_2), .A0 (nx7162), .A1 (nx7164), .S0 (
          nx8524)) ;
    inv01 ix7161 (.Y (nx7162), .A (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_2)) ;
    inv01 ix7163 (.Y (nx7164), .A (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_2)) ;
    mux21 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix213 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BoothOperand_3), .A0 (nx7166), .A1 (nx7168), .S0 (
          nx8524)) ;
    inv01 ix7165 (.Y (nx7166), .A (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_3)) ;
    inv01 ix7167 (.Y (nx7168), .A (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_3)) ;
    mux21 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix221 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BoothOperand_4), .A0 (nx7170), .A1 (nx7172), .S0 (
          nx8524)) ;
    inv01 ix7169 (.Y (nx7170), .A (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_4)) ;
    inv01 ix7171 (.Y (nx7172), .A (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_4)) ;
    mux21 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix229 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BoothOperand_5), .A0 (nx7174), .A1 (nx7176), .S0 (
          nx8526)) ;
    inv01 ix7173 (.Y (nx7174), .A (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_5)) ;
    inv01 ix7175 (.Y (nx7176), .A (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_5)) ;
    mux21 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix237 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BoothOperand_6), .A0 (nx7178), .A1 (nx7180), .S0 (
          nx8526)) ;
    inv01 ix7177 (.Y (nx7178), .A (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_6)) ;
    inv01 ix7179 (.Y (nx7180), .A (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_6)) ;
    mux21 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix245 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BoothOperand_7), .A0 (nx7182), .A1 (nx7184), .S0 (
          nx8526)) ;
    inv01 ix7181 (.Y (nx7182), .A (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_7)) ;
    inv01 ix7183 (.Y (nx7184), .A (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_7)) ;
    mux21 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix253 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BoothOperand_8), .A0 (nx7186), .A1 (nx7188), .S0 (
          nx8526)) ;
    inv01 ix7185 (.Y (nx7186), .A (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_8)) ;
    inv01 ix7187 (.Y (nx7188), .A (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_8)) ;
    mux21 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix261 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BoothOperand_9), .A0 (nx7190), .A1 (nx7192), .S0 (
          nx8526)) ;
    inv01 ix7189 (.Y (nx7190), .A (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_9)) ;
    inv01 ix7191 (.Y (nx7192), .A (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_9)) ;
    mux21 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix269 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BoothOperand_10), .A0 (nx7194), .A1 (nx7196), .S0 (
          nx8526)) ;
    inv01 ix7193 (.Y (nx7194), .A (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_10)) ;
    inv01 ix7195 (.Y (nx7196), .A (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_10)) ;
    mux21 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix277 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BoothOperand_11), .A0 (nx7198), .A1 (nx7200), .S0 (
          nx8526)) ;
    inv01 ix7197 (.Y (nx7198), .A (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_11)) ;
    inv01 ix7199 (.Y (nx7200), .A (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_11)) ;
    mux21 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix285 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BoothOperand_12), .A0 (nx7202), .A1 (nx7204), .S0 (
          nx8528)) ;
    inv01 ix7201 (.Y (nx7202), .A (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_12)) ;
    inv01 ix7203 (.Y (nx7204), .A (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_12)) ;
    mux21 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix293 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BoothOperand_13), .A0 (nx7206), .A1 (nx7208), .S0 (
          nx8528)) ;
    inv01 ix7205 (.Y (nx7206), .A (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_13)) ;
    inv01 ix7207 (.Y (nx7208), .A (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_13)) ;
    mux21 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix301 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BoothOperand_14), .A0 (nx7210), .A1 (nx7212), .S0 (
          nx8528)) ;
    inv01 ix7209 (.Y (nx7210), .A (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_14)) ;
    inv01 ix7211 (.Y (nx7212), .A (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_14)) ;
    mux21 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix309 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BoothOperand_15), .A0 (nx7214), .A1 (nx7216), .S0 (
          nx8528)) ;
    inv01 ix7213 (.Y (nx7214), .A (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_15)) ;
    inv01 ix7215 (.Y (nx7216), .A (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_15)) ;
    mux21 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix317 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BoothOperand_16), .A0 (nx7218), .A1 (nx7220), .S0 (
          nx8528)) ;
    inv01 ix7217 (.Y (nx7218), .A (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_16)) ;
    inv01 ix7219 (.Y (nx7220), .A (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_16)) ;
    xnor2 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_ix321 (.Y (
          L1_4_L2_3_G5_MINI_ALU_AddPToBoothOperand), .A0 (nx8528), .A1 (nx7086)
          ) ;
    oai32 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix393 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .A0 (nx8734), .A1 (
          RST), .A2 (nx8538), .B0 (nx7156), .B1 (nx7224)) ;
    oai32 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix403 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .A0 (nx8734), .A1 (
          RST), .A2 (nx8538), .B0 (nx7160), .B1 (nx7224)) ;
    oai32 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix413 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .A0 (nx8734), .A1 (
          RST), .A2 (nx8538), .B0 (nx7164), .B1 (nx7224)) ;
    oai32 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix423 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .A0 (nx8734), .A1 (
          RST), .A2 (nx8538), .B0 (nx7168), .B1 (nx7224)) ;
    oai32 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix433 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .A0 (nx8734), .A1 (
          RST), .A2 (nx8538), .B0 (nx7172), .B1 (nx7224)) ;
    oai32 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix443 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .A0 (nx8734), .A1 (
          RST), .A2 (nx8538), .B0 (nx7176), .B1 (nx7224)) ;
    oai32 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix453 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .A0 (nx8734), .A1 (
          RST), .A2 (nx8540), .B0 (nx7180), .B1 (nx7224)) ;
    oai32 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix463 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .A0 (nx8736), .A1 (
          RST), .A2 (nx8540), .B0 (nx7184), .B1 (nx7226)) ;
    oai32 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix473 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .A0 (nx8736), .A1 (
          RST), .A2 (nx8540), .B0 (nx7188), .B1 (nx7226)) ;
    oai32 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix483 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .A0 (nx7228), .A1 (
          RST), .A2 (nx8540), .B0 (nx7192), .B1 (nx7226)) ;
    inv01 ix7227 (.Y (nx7228), .A (FilterDin_4__3__0)) ;
    oai32 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix493 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .A0 (nx7230), .A1 (
          RST), .A2 (nx8540), .B0 (nx7196), .B1 (nx7226)) ;
    inv01 ix7229 (.Y (nx7230), .A (FilterDin_4__3__1)) ;
    oai32 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix503 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .A0 (nx7232), .A1 (
          RST), .A2 (nx8540), .B0 (nx7200), .B1 (nx7226)) ;
    inv01 ix7231 (.Y (nx7232), .A (FilterDin_4__3__2)) ;
    oai32 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix513 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .A0 (nx7234), .A1 (
          RST), .A2 (nx8540), .B0 (nx7204), .B1 (nx7226)) ;
    inv01 ix7233 (.Y (nx7234), .A (FilterDin_4__3__3)) ;
    oai32 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix523 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .A0 (nx7236), .A1 (
          RST), .A2 (nx8542), .B0 (nx7208), .B1 (nx7226)) ;
    inv01 ix7235 (.Y (nx7236), .A (FilterDin_4__3__4)) ;
    oai32 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix533 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .A0 (nx7238), .A1 (
          RST), .A2 (nx8542), .B0 (nx7212), .B1 (nx7240)) ;
    inv01 ix7237 (.Y (nx7238), .A (FilterDin_4__3__5)) ;
    inv01 ix7239 (.Y (nx7240), .A (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566)) ;
    oai32 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix543 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .A0 (nx7242), .A1 (
          RST), .A2 (nx8542), .B0 (nx7216), .B1 (nx7240)) ;
    inv01 ix7241 (.Y (nx7242), .A (FilterDin_4__3__6)) ;
    oai32 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix553 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .A0 (nx7244), .A1 (
          RST), .A2 (nx8542), .B0 (nx7220), .B1 (nx7240)) ;
    inv01 ix7243 (.Y (nx7244), .A (FilterDin_4__3__7)) ;
    nand02_2x L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix633 (.Y (nx7224), .A0 (
              nx7614), .A1 (nx8542)) ;
    nand02_2x L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix635 (.Y (nx7226), .A0 (
              nx7614), .A1 (nx8542)) ;
    oai32 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix393 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .A0 (nx8736), .A1 (
          RST), .A2 (nx8544), .B0 (nx7154), .B1 (nx7246)) ;
    oai32 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix403 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .A0 (nx8736), .A1 (
          RST), .A2 (nx8544), .B0 (nx7158), .B1 (nx7246)) ;
    oai32 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix413 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .A0 (nx8736), .A1 (
          RST), .A2 (nx8544), .B0 (nx7162), .B1 (nx7246)) ;
    oai32 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix423 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .A0 (nx8736), .A1 (
          RST), .A2 (nx8544), .B0 (nx7166), .B1 (nx7246)) ;
    oai32 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix433 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .A0 (nx8736), .A1 (
          RST), .A2 (nx8544), .B0 (nx7170), .B1 (nx7246)) ;
    oai32 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix443 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .A0 (nx8738), .A1 (
          RST), .A2 (nx8544), .B0 (nx7174), .B1 (nx7246)) ;
    oai32 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix453 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .A0 (nx8738), .A1 (
          RST), .A2 (nx8546), .B0 (nx7178), .B1 (nx7246)) ;
    oai32 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix463 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .A0 (nx8738), .A1 (
          RST), .A2 (nx8546), .B0 (nx7182), .B1 (nx7248)) ;
    oai32 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix473 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .A0 (nx8738), .A1 (
          RST), .A2 (nx8546), .B0 (nx7186), .B1 (nx7248)) ;
    oai32 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix483 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .A0 (nx7228), .A1 (
          RST), .A2 (nx8546), .B0 (nx7190), .B1 (nx7248)) ;
    oai32 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix493 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .A0 (nx7250), .A1 (
          RST), .A2 (nx8546), .B0 (nx7194), .B1 (nx7248)) ;
    inv01 ix7249 (.Y (nx7250), .A (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_10)) ;
    oai32 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix503 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .A0 (nx7252), .A1 (
          RST), .A2 (nx8546), .B0 (nx7198), .B1 (nx7248)) ;
    inv01 ix7251 (.Y (nx7252), .A (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_11)) ;
    oai32 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix513 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .A0 (nx7254), .A1 (
          RST), .A2 (nx8546), .B0 (nx7202), .B1 (nx7248)) ;
    inv01 ix7253 (.Y (nx7254), .A (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_12)) ;
    oai32 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix523 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .A0 (nx7256), .A1 (
          RST), .A2 (nx8548), .B0 (nx7206), .B1 (nx7248)) ;
    inv01 ix7255 (.Y (nx7256), .A (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_13)) ;
    oai32 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix533 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .A0 (nx7258), .A1 (
          RST), .A2 (nx8548), .B0 (nx7210), .B1 (nx7260)) ;
    inv01 ix7257 (.Y (nx7258), .A (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_14)) ;
    inv01 ix7259 (.Y (nx7260), .A (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566)) ;
    oai32 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix543 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .A0 (nx7262), .A1 (
          RST), .A2 (nx8548), .B0 (nx7214), .B1 (nx7260)) ;
    inv01 ix7261 (.Y (nx7262), .A (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_15)) ;
    oai32 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix553 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .A0 (nx7264), .A1 (
          RST), .A2 (nx8548), .B0 (nx7218), .B1 (nx7260)) ;
    inv01 ix7263 (.Y (nx7264), .A (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_16)) ;
    nand02_2x L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix633 (.Y (nx7246), .A0 (
              nx7616), .A1 (nx8548)) ;
    nand02_2x L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix635 (.Y (nx7248), .A0 (
              nx7616), .A1 (nx8548)) ;
    oai32 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix393 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .A0 (nx7266), .A1 (
          RST), .A2 (nx8550), .B0 (L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_nx384), .B1 (
          nx7268)) ;
    inv01 ix7265 (.Y (nx7266), .A (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_0)) ;
    oai32 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix403 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .A0 (nx7270), .A1 (
          RST), .A2 (nx8550), .B0 (nx7086), .B1 (nx7268)) ;
    inv01 ix7269 (.Y (nx7270), .A (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_1)) ;
    oai32 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix413 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .A0 (nx7272), .A1 (
          RST), .A2 (nx8550), .B0 (L1_4_L2_3_G5_MINI_ALU_nx387), .B1 (nx7268)) ;
    inv01 ix7271 (.Y (nx7272), .A (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_2)) ;
    oai32 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix423 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .A0 (nx7274), .A1 (
          RST), .A2 (nx8550), .B0 (L1_4_L2_3_G5_MINI_ALU_nx399), .B1 (nx7268)) ;
    inv01 ix7273 (.Y (nx7274), .A (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_3)) ;
    oai32 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix433 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .A0 (nx7276), .A1 (
          RST), .A2 (nx8550), .B0 (L1_4_L2_3_G5_MINI_ALU_nx409), .B1 (nx7268)) ;
    inv01 ix7275 (.Y (nx7276), .A (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_4)) ;
    oai32 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix443 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .A0 (nx7278), .A1 (
          RST), .A2 (nx8550), .B0 (L1_4_L2_3_G5_MINI_ALU_nx419), .B1 (nx7268)) ;
    inv01 ix7277 (.Y (nx7278), .A (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_5)) ;
    oai32 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix453 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .A0 (nx7280), .A1 (
          RST), .A2 (nx8550), .B0 (L1_4_L2_3_G5_MINI_ALU_nx429), .B1 (nx7268)) ;
    inv01 ix7279 (.Y (nx7280), .A (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_6)) ;
    oai32 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix463 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .A0 (nx7282), .A1 (
          RST), .A2 (nx8552), .B0 (L1_4_L2_3_G5_MINI_ALU_nx439), .B1 (nx7284)) ;
    inv01 ix7281 (.Y (nx7282), .A (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_7)) ;
    oai32 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix473 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .A0 (nx7286), .A1 (
          RST), .A2 (nx8552), .B0 (L1_4_L2_3_G5_MINI_ALU_nx449), .B1 (nx7284)) ;
    inv01 ix7285 (.Y (nx7286), .A (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_8)) ;
    oai32 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix483 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .A0 (nx7288), .A1 (
          RST), .A2 (nx8552), .B0 (L1_4_L2_3_G5_MINI_ALU_nx469), .B1 (nx7284)) ;
    inv01 ix7287 (.Y (nx7288), .A (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_9)) ;
    oai32 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix493 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .A0 (nx7290), .A1 (
          RST), .A2 (nx8552), .B0 (L1_4_L2_3_G5_MINI_ALU_nx477), .B1 (nx7284)) ;
    inv01 ix7289 (.Y (nx7290), .A (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_10)) ;
    oai32 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix503 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .A0 (nx7292), .A1 (
          RST), .A2 (nx8552), .B0 (L1_4_L2_3_G5_MINI_ALU_nx485), .B1 (nx7284)) ;
    inv01 ix7291 (.Y (nx7292), .A (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_11)) ;
    oai32 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix513 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .A0 (nx7294), .A1 (
          RST), .A2 (nx8552), .B0 (L1_4_L2_3_G5_MINI_ALU_nx493), .B1 (nx7284)) ;
    inv01 ix7293 (.Y (nx7294), .A (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_12)) ;
    oai32 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix523 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .A0 (nx7296), .A1 (
          RST), .A2 (nx8552), .B0 (L1_4_L2_3_G5_MINI_ALU_nx501), .B1 (nx7284)) ;
    inv01 ix7295 (.Y (nx7296), .A (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_13)) ;
    oai32 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix533 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .A0 (nx7298), .A1 (
          RST), .A2 (nx8554), .B0 (L1_4_L2_3_G5_MINI_ALU_nx509), .B1 (nx7300)) ;
    inv01 ix7297 (.Y (nx7298), .A (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_14)) ;
    inv01 ix7299 (.Y (nx7300), .A (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566)) ;
    oai32 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix543 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .A0 (nx7302), .A1 (
          RST), .A2 (nx8554), .B0 (L1_4_L2_3_G5_MINI_ALU_nx517), .B1 (nx7300)) ;
    inv01 ix7301 (.Y (nx7302), .A (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_15)) ;
    oai32 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix553 (.Y (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .A0 (nx7304), .A1 (
          RST), .A2 (nx8554), .B0 (nx7102), .B1 (nx7300)) ;
    inv01 ix7303 (.Y (nx7304), .A (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_16)) ;
    nand02_2x L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix633 (.Y (nx7268), .A0 (
              nx7616), .A1 (nx8554)) ;
    nand02_2x L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix635 (.Y (nx7284), .A0 (
              nx7616), .A1 (nx8554)) ;
    mux21 L1_4_L2_4_G5_MINI_ALU_ix404 (.Y (L1_4_L2_4_G5_MINI_ALU_nx403), .A0 (
          nx7306), .A1 (L1_4_L2_4_G5_MINI_ALU_BoothP_2), .S0 (
          L1_4_L2_4_G5_MINI_ALU_nx395)) ;
    inv01 ix7305 (.Y (nx7306), .A (L1_4_L2_4_G5_MINI_ALU_nx391)) ;
    mux21 L1_4_L2_4_G5_MINI_ALU_ix414 (.Y (L1_4_L2_4_G5_MINI_ALU_nx413), .A0 (
          nx7308), .A1 (L1_4_L2_4_G5_MINI_ALU_BoothP_3), .S0 (
          L1_4_L2_4_G5_MINI_ALU_nx405)) ;
    inv01 ix7307 (.Y (nx7308), .A (L1_4_L2_4_G5_MINI_ALU_nx403)) ;
    mux21 L1_4_L2_4_G5_MINI_ALU_ix424 (.Y (L1_4_L2_4_G5_MINI_ALU_nx423), .A0 (
          nx7310), .A1 (L1_4_L2_4_G5_MINI_ALU_BoothP_4), .S0 (
          L1_4_L2_4_G5_MINI_ALU_nx415)) ;
    inv01 ix7309 (.Y (nx7310), .A (L1_4_L2_4_G5_MINI_ALU_nx413)) ;
    mux21 L1_4_L2_4_G5_MINI_ALU_ix434 (.Y (L1_4_L2_4_G5_MINI_ALU_nx433), .A0 (
          nx7312), .A1 (L1_4_L2_4_G5_MINI_ALU_BoothP_5), .S0 (
          L1_4_L2_4_G5_MINI_ALU_nx425)) ;
    inv01 ix7311 (.Y (nx7312), .A (L1_4_L2_4_G5_MINI_ALU_nx423)) ;
    mux21 L1_4_L2_4_G5_MINI_ALU_ix444 (.Y (L1_4_L2_4_G5_MINI_ALU_nx443), .A0 (
          nx7314), .A1 (L1_4_L2_4_G5_MINI_ALU_BoothP_6), .S0 (
          L1_4_L2_4_G5_MINI_ALU_nx435)) ;
    inv01 ix7313 (.Y (nx7314), .A (L1_4_L2_4_G5_MINI_ALU_nx433)) ;
    mux21 L1_4_L2_4_G5_MINI_ALU_ix454 (.Y (L1_4_L2_4_G5_MINI_ALU_nx453), .A0 (
          nx7316), .A1 (L1_4_L2_4_G5_MINI_ALU_BoothP_7), .S0 (
          L1_4_L2_4_G5_MINI_ALU_nx445)) ;
    inv01 ix7315 (.Y (nx7316), .A (L1_4_L2_4_G5_MINI_ALU_nx443)) ;
    mux21 L1_4_L2_4_G5_MINI_ALU_ix462 (.Y (L1_4_L2_4_G5_MINI_ALU_nx461), .A0 (
          nx7318), .A1 (L1_4_L2_4_G5_MINI_ALU_BoothP_8), .S0 (
          L1_4_L2_4_G5_MINI_ALU_nx455)) ;
    inv01 ix7317 (.Y (nx7318), .A (L1_4_L2_4_G5_MINI_ALU_nx453)) ;
    mux21 L1_4_L2_4_G5_MINI_ALU_ix468 (.Y (L1_4_L2_4_G5_MINI_ALU_nx467), .A0 (
          nx7320), .A1 (L1_4_L2_4_G5_MINI_ALU_BoothP_9), .S0 (
          L1_4_L2_4_G5_MINI_ALU_nx463)) ;
    inv01 ix7319 (.Y (nx7320), .A (L1_4_L2_4_G5_MINI_ALU_nx461)) ;
    mux21 L1_4_L2_4_G5_MINI_ALU_ix476 (.Y (L1_4_L2_4_G5_MINI_ALU_nx475), .A0 (
          nx7322), .A1 (L1_4_L2_4_G5_MINI_ALU_BoothP_10), .S0 (
          L1_4_L2_4_G5_MINI_ALU_nx471)) ;
    inv01 ix7321 (.Y (nx7322), .A (L1_4_L2_4_G5_MINI_ALU_nx467)) ;
    mux21 L1_4_L2_4_G5_MINI_ALU_ix484 (.Y (L1_4_L2_4_G5_MINI_ALU_nx483), .A0 (
          nx7324), .A1 (L1_4_L2_4_G5_MINI_ALU_BoothP_11), .S0 (
          L1_4_L2_4_G5_MINI_ALU_nx479)) ;
    inv01 ix7323 (.Y (nx7324), .A (L1_4_L2_4_G5_MINI_ALU_nx475)) ;
    mux21 L1_4_L2_4_G5_MINI_ALU_ix492 (.Y (L1_4_L2_4_G5_MINI_ALU_nx491), .A0 (
          nx7326), .A1 (L1_4_L2_4_G5_MINI_ALU_BoothP_12), .S0 (
          L1_4_L2_4_G5_MINI_ALU_nx487)) ;
    inv01 ix7325 (.Y (nx7326), .A (L1_4_L2_4_G5_MINI_ALU_nx483)) ;
    mux21 L1_4_L2_4_G5_MINI_ALU_ix500 (.Y (L1_4_L2_4_G5_MINI_ALU_nx499), .A0 (
          nx7328), .A1 (L1_4_L2_4_G5_MINI_ALU_BoothP_13), .S0 (
          L1_4_L2_4_G5_MINI_ALU_nx495)) ;
    inv01 ix7327 (.Y (nx7328), .A (L1_4_L2_4_G5_MINI_ALU_nx491)) ;
    mux21 L1_4_L2_4_G5_MINI_ALU_ix508 (.Y (L1_4_L2_4_G5_MINI_ALU_nx507), .A0 (
          nx7330), .A1 (L1_4_L2_4_G5_MINI_ALU_BoothP_14), .S0 (
          L1_4_L2_4_G5_MINI_ALU_nx503)) ;
    inv01 ix7329 (.Y (nx7330), .A (L1_4_L2_4_G5_MINI_ALU_nx499)) ;
    mux21 L1_4_L2_4_G5_MINI_ALU_ix516 (.Y (L1_4_L2_4_G5_MINI_ALU_nx515), .A0 (
          nx7332), .A1 (L1_4_L2_4_G5_MINI_ALU_BoothP_15), .S0 (
          L1_4_L2_4_G5_MINI_ALU_nx511)) ;
    inv01 ix7331 (.Y (nx7332), .A (L1_4_L2_4_G5_MINI_ALU_nx507)) ;
    mux21 L1_4_L2_4_G5_MINI_ALU_ix161 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_1), .A0 (nx7334), .A1 (
          L1_4_L2_4_G5_MINI_ALU_nx379), .S0 (nx8558)) ;
    inv01 ix7333 (.Y (nx7334), .A (L1_4_L2_4_G5_MINI_ALU_BoothP_1)) ;
    mux21 L1_4_L2_4_G5_MINI_ALU_ix181 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_2), .A0 (
          L1_4_L2_4_G5_MINI_ALU_nx387), .A1 (L1_4_L2_4_G5_MINI_ALU_nx389), .S0 (
          nx8558)) ;
    mux21 L1_4_L2_4_G5_MINI_ALU_ix201 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_3), .A0 (
          L1_4_L2_4_G5_MINI_ALU_nx399), .A1 (L1_4_L2_4_G5_MINI_ALU_nx401), .S0 (
          nx8558)) ;
    mux21 L1_4_L2_4_G5_MINI_ALU_ix221 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_4), .A0 (
          L1_4_L2_4_G5_MINI_ALU_nx409), .A1 (L1_4_L2_4_G5_MINI_ALU_nx411), .S0 (
          nx8558)) ;
    mux21 L1_4_L2_4_G5_MINI_ALU_ix241 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_5), .A0 (
          L1_4_L2_4_G5_MINI_ALU_nx419), .A1 (L1_4_L2_4_G5_MINI_ALU_nx421), .S0 (
          nx8558)) ;
    mux21 L1_4_L2_4_G5_MINI_ALU_ix261 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_6), .A0 (
          L1_4_L2_4_G5_MINI_ALU_nx429), .A1 (L1_4_L2_4_G5_MINI_ALU_nx431), .S0 (
          nx8558)) ;
    mux21 L1_4_L2_4_G5_MINI_ALU_ix281 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_7), .A0 (
          L1_4_L2_4_G5_MINI_ALU_nx439), .A1 (L1_4_L2_4_G5_MINI_ALU_nx441), .S0 (
          nx8558)) ;
    mux21 L1_4_L2_4_G5_MINI_ALU_ix301 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_8), .A0 (
          L1_4_L2_4_G5_MINI_ALU_nx449), .A1 (L1_4_L2_4_G5_MINI_ALU_nx451), .S0 (
          nx8560)) ;
    mux21 L1_4_L2_4_G5_MINI_ALU_ix321 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_9), .A0 (
          L1_4_L2_4_G5_MINI_ALU_nx469), .A1 (nx7336), .S0 (nx8560)) ;
    inv01 ix7335 (.Y (nx7336), .A (L1_4_L2_4_G5_MINI_ALU_nx316)) ;
    mux21 L1_4_L2_4_G5_MINI_ALU_ix341 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_10), .A0 (
          L1_4_L2_4_G5_MINI_ALU_nx477), .A1 (nx7338), .S0 (nx8560)) ;
    inv01 ix7337 (.Y (nx7338), .A (L1_4_L2_4_G5_MINI_ALU_nx336)) ;
    mux21 L1_4_L2_4_G5_MINI_ALU_ix361 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_11), .A0 (
          L1_4_L2_4_G5_MINI_ALU_nx485), .A1 (nx7340), .S0 (nx8560)) ;
    inv01 ix7339 (.Y (nx7340), .A (L1_4_L2_4_G5_MINI_ALU_nx356)) ;
    mux21 L1_4_L2_4_G5_MINI_ALU_ix381 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_12), .A0 (
          L1_4_L2_4_G5_MINI_ALU_nx493), .A1 (nx7342), .S0 (nx8560)) ;
    inv01 ix7341 (.Y (nx7342), .A (L1_4_L2_4_G5_MINI_ALU_nx376)) ;
    mux21 L1_4_L2_4_G5_MINI_ALU_ix401 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_13), .A0 (
          L1_4_L2_4_G5_MINI_ALU_nx501), .A1 (nx7344), .S0 (nx8560)) ;
    inv01 ix7343 (.Y (nx7344), .A (L1_4_L2_4_G5_MINI_ALU_nx396)) ;
    mux21 L1_4_L2_4_G5_MINI_ALU_ix421 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_14), .A0 (
          L1_4_L2_4_G5_MINI_ALU_nx509), .A1 (nx7346), .S0 (nx8560)) ;
    inv01 ix7345 (.Y (nx7346), .A (L1_4_L2_4_G5_MINI_ALU_nx416)) ;
    mux21 L1_4_L2_4_G5_MINI_ALU_ix441 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_15), .A0 (
          L1_4_L2_4_G5_MINI_ALU_nx517), .A1 (nx7348), .S0 (nx8562)) ;
    inv01 ix7347 (.Y (nx7348), .A (L1_4_L2_4_G5_MINI_ALU_nx436)) ;
    mux21 L1_4_L2_4_G5_MINI_ALU_ix461 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_16), .A0 (nx7350), .A1 (nx7352
          ), .S0 (nx8562)) ;
    inv01 ix7349 (.Y (nx7350), .A (L1_4_L2_4_G5_MINI_ALU_BoothP_16)) ;
    inv01 ix7351 (.Y (nx7352), .A (L1_4_L2_4_G5_MINI_ALU_nx456)) ;
    nor02_2x L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix319 (.Y (
             L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx642), .A0 (Start), .A1 (
             CalculatingBooth_dup_1253)) ;
    nor02_2x L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix85 (.Y (
             L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_0), .A0 (nx8572), .A1 (
             nx7354)) ;
    inv01 ix7353 (.Y (nx7354), .A (L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_1)) ;
    mux21 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix125 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_1), .A0 (nx7356), .A1 (
          nx7358), .S0 (nx8572)) ;
    inv01 ix7355 (.Y (nx7356), .A (L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_2)) ;
    inv01 ix7357 (.Y (nx7358), .A (WindowDin_4__4__0)) ;
    mux21 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix133 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_2), .A0 (nx7360), .A1 (
          nx7362), .S0 (nx8572)) ;
    inv01 ix7359 (.Y (nx7360), .A (L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_3)) ;
    inv01 ix7361 (.Y (nx7362), .A (WindowDin_4__4__1)) ;
    mux21 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix141 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_3), .A0 (nx7364), .A1 (
          nx7366), .S0 (nx8572)) ;
    inv01 ix7363 (.Y (nx7364), .A (L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_4)) ;
    inv01 ix7365 (.Y (nx7366), .A (WindowDin_4__4__2)) ;
    mux21 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix149 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_4), .A0 (nx7368), .A1 (
          nx7370), .S0 (nx8572)) ;
    inv01 ix7367 (.Y (nx7368), .A (L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_5)) ;
    inv01 ix7369 (.Y (nx7370), .A (WindowDin_4__4__3)) ;
    mux21 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix157 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_5), .A0 (nx7372), .A1 (
          nx7374), .S0 (nx8572)) ;
    inv01 ix7371 (.Y (nx7372), .A (L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_6)) ;
    inv01 ix7373 (.Y (nx7374), .A (WindowDin_4__4__4)) ;
    mux21 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix165 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_6), .A0 (nx7376), .A1 (
          nx7378), .S0 (nx8572)) ;
    inv01 ix7375 (.Y (nx7376), .A (L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_7)) ;
    inv01 ix7377 (.Y (nx7378), .A (WindowDin_4__4__5)) ;
    mux21 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix173 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_7), .A0 (nx7380), .A1 (
          nx7382), .S0 (nx8574)) ;
    inv01 ix7379 (.Y (nx7380), .A (L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_8)) ;
    inv01 ix7381 (.Y (nx7382), .A (WindowDin_4__4__6)) ;
    mux21 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix181 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_8), .A0 (nx7384), .A1 (
          nx7386), .S0 (nx8574)) ;
    inv01 ix7383 (.Y (nx7384), .A (L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_9)) ;
    inv01 ix7385 (.Y (nx7386), .A (WindowDin_4__4__7)) ;
    nor02_2x L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix89 (.Y (
             L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_9), .A0 (nx8574), .A1 (
             nx7388)) ;
    inv01 ix7387 (.Y (nx7388), .A (L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_10)
          ) ;
    nor02_2x L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix93 (.Y (
             L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_10), .A0 (nx8574), .A1 (
             nx7390)) ;
    inv01 ix7389 (.Y (nx7390), .A (L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_11)
          ) ;
    nor02_2x L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix97 (.Y (
             L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_11), .A0 (nx8574), .A1 (
             nx7392)) ;
    inv01 ix7391 (.Y (nx7392), .A (L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_12)
          ) ;
    nor02_2x L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix101 (.Y (
             L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_12), .A0 (nx8574), .A1 (
             nx7394)) ;
    inv01 ix7393 (.Y (nx7394), .A (L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_13)
          ) ;
    nor02_2x L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix105 (.Y (
             L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_13), .A0 (nx8574), .A1 (
             nx7396)) ;
    inv01 ix7395 (.Y (nx7396), .A (L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_14)
          ) ;
    nor02_2x L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix109 (.Y (
             L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_14), .A0 (nx8576), .A1 (
             nx7398)) ;
    inv01 ix7397 (.Y (nx7398), .A (L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_15)
          ) ;
    nor02_2x L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix113 (.Y (
             L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_15), .A0 (nx8576), .A1 (
             nx7400)) ;
    inv01 ix7399 (.Y (nx7400), .A (L1_4_L2_4_G5_MINI_ALU_BoothPBeforeShift_16)
          ) ;
    nor02_2x L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix117 (.Y (
             L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_16), .A0 (nx8576), .A1 (
             nx7400)) ;
    mux21 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix189 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BoothOperand_0), .A0 (nx7402), .A1 (nx7404), .S0 (
          nx8564)) ;
    inv01 ix7401 (.Y (nx7402), .A (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_0)) ;
    inv01 ix7403 (.Y (nx7404), .A (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_0)) ;
    mux21 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix197 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BoothOperand_1), .A0 (nx7406), .A1 (nx7408), .S0 (
          nx8564)) ;
    inv01 ix7405 (.Y (nx7406), .A (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_1)) ;
    inv01 ix7407 (.Y (nx7408), .A (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_1)) ;
    mux21 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix205 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BoothOperand_2), .A0 (nx7410), .A1 (nx7412), .S0 (
          nx8564)) ;
    inv01 ix7409 (.Y (nx7410), .A (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_2)) ;
    inv01 ix7411 (.Y (nx7412), .A (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_2)) ;
    mux21 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix213 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BoothOperand_3), .A0 (nx7414), .A1 (nx7416), .S0 (
          nx8564)) ;
    inv01 ix7413 (.Y (nx7414), .A (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_3)) ;
    inv01 ix7415 (.Y (nx7416), .A (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_3)) ;
    mux21 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix221 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BoothOperand_4), .A0 (nx7418), .A1 (nx7420), .S0 (
          nx8564)) ;
    inv01 ix7417 (.Y (nx7418), .A (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_4)) ;
    inv01 ix7419 (.Y (nx7420), .A (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_4)) ;
    mux21 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix229 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BoothOperand_5), .A0 (nx7422), .A1 (nx7424), .S0 (
          nx8566)) ;
    inv01 ix7421 (.Y (nx7422), .A (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_5)) ;
    inv01 ix7423 (.Y (nx7424), .A (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_5)) ;
    mux21 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix237 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BoothOperand_6), .A0 (nx7426), .A1 (nx7428), .S0 (
          nx8566)) ;
    inv01 ix7425 (.Y (nx7426), .A (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_6)) ;
    inv01 ix7427 (.Y (nx7428), .A (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_6)) ;
    mux21 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix245 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BoothOperand_7), .A0 (nx7430), .A1 (nx7432), .S0 (
          nx8566)) ;
    inv01 ix7429 (.Y (nx7430), .A (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_7)) ;
    inv01 ix7431 (.Y (nx7432), .A (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_7)) ;
    mux21 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix253 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BoothOperand_8), .A0 (nx7434), .A1 (nx7436), .S0 (
          nx8566)) ;
    inv01 ix7433 (.Y (nx7434), .A (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_8)) ;
    inv01 ix7435 (.Y (nx7436), .A (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_8)) ;
    mux21 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix261 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BoothOperand_9), .A0 (nx7438), .A1 (nx7440), .S0 (
          nx8566)) ;
    inv01 ix7437 (.Y (nx7438), .A (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_9)) ;
    inv01 ix7439 (.Y (nx7440), .A (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_9)) ;
    mux21 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix269 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BoothOperand_10), .A0 (nx7442), .A1 (nx7444), .S0 (
          nx8566)) ;
    inv01 ix7441 (.Y (nx7442), .A (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_10)) ;
    inv01 ix7443 (.Y (nx7444), .A (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_10)) ;
    mux21 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix277 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BoothOperand_11), .A0 (nx7446), .A1 (nx7448), .S0 (
          nx8566)) ;
    inv01 ix7445 (.Y (nx7446), .A (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_11)) ;
    inv01 ix7447 (.Y (nx7448), .A (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_11)) ;
    mux21 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix285 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BoothOperand_12), .A0 (nx7450), .A1 (nx7452), .S0 (
          nx8568)) ;
    inv01 ix7449 (.Y (nx7450), .A (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_12)) ;
    inv01 ix7451 (.Y (nx7452), .A (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_12)) ;
    mux21 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix293 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BoothOperand_13), .A0 (nx7454), .A1 (nx7456), .S0 (
          nx8568)) ;
    inv01 ix7453 (.Y (nx7454), .A (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_13)) ;
    inv01 ix7455 (.Y (nx7456), .A (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_13)) ;
    mux21 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix301 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BoothOperand_14), .A0 (nx7458), .A1 (nx7460), .S0 (
          nx8568)) ;
    inv01 ix7457 (.Y (nx7458), .A (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_14)) ;
    inv01 ix7459 (.Y (nx7460), .A (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_14)) ;
    mux21 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix309 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BoothOperand_15), .A0 (nx7462), .A1 (nx7464), .S0 (
          nx8568)) ;
    inv01 ix7461 (.Y (nx7462), .A (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_15)) ;
    inv01 ix7463 (.Y (nx7464), .A (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_15)) ;
    mux21 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix317 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BoothOperand_16), .A0 (nx7466), .A1 (nx7468), .S0 (
          nx8568)) ;
    inv01 ix7465 (.Y (nx7466), .A (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDout_16)) ;
    inv01 ix7467 (.Y (nx7468), .A (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterADout_16)) ;
    xnor2 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_ix321 (.Y (
          L1_4_L2_4_G5_MINI_ALU_AddPToBoothOperand), .A0 (nx8568), .A1 (nx7334)
          ) ;
    oai32 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix393 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx392), .A0 (nx8740), .A1 (
          RST), .A2 (nx8578), .B0 (nx7404), .B1 (nx7472)) ;
    oai32 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix403 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx402), .A0 (nx8740), .A1 (
          RST), .A2 (nx8578), .B0 (nx7408), .B1 (nx7472)) ;
    oai32 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix413 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx412), .A0 (nx8740), .A1 (
          RST), .A2 (nx8578), .B0 (nx7412), .B1 (nx7472)) ;
    oai32 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix423 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx422), .A0 (nx8740), .A1 (
          RST), .A2 (nx8578), .B0 (nx7416), .B1 (nx7472)) ;
    oai32 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix433 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx432), .A0 (nx8740), .A1 (
          RST), .A2 (nx8578), .B0 (nx7420), .B1 (nx7472)) ;
    oai32 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix443 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx442), .A0 (nx8740), .A1 (
          RST), .A2 (nx8578), .B0 (nx7424), .B1 (nx7472)) ;
    oai32 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix453 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx452), .A0 (nx8740), .A1 (
          RST), .A2 (nx8580), .B0 (nx7428), .B1 (nx7472)) ;
    oai32 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix463 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx462), .A0 (nx8742), .A1 (
          RST), .A2 (nx8580), .B0 (nx7432), .B1 (nx7474)) ;
    oai32 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix473 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx472), .A0 (nx8742), .A1 (
          RST), .A2 (nx8580), .B0 (nx7436), .B1 (nx7474)) ;
    oai32 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix483 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx482), .A0 (nx7476), .A1 (
          RST), .A2 (nx8580), .B0 (nx7440), .B1 (nx7474)) ;
    inv01 ix7475 (.Y (nx7476), .A (FilterDin_4__4__0)) ;
    oai32 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix493 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx492), .A0 (nx7478), .A1 (
          RST), .A2 (nx8580), .B0 (nx7444), .B1 (nx7474)) ;
    inv01 ix7477 (.Y (nx7478), .A (FilterDin_4__4__1)) ;
    oai32 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix503 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx502), .A0 (nx7480), .A1 (
          RST), .A2 (nx8580), .B0 (nx7448), .B1 (nx7474)) ;
    inv01 ix7479 (.Y (nx7480), .A (FilterDin_4__4__2)) ;
    oai32 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix513 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx512), .A0 (nx7482), .A1 (
          RST), .A2 (nx8580), .B0 (nx7452), .B1 (nx7474)) ;
    inv01 ix7481 (.Y (nx7482), .A (FilterDin_4__4__3)) ;
    oai32 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix523 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx522), .A0 (nx7484), .A1 (
          RST), .A2 (nx8582), .B0 (nx7456), .B1 (nx7474)) ;
    inv01 ix7483 (.Y (nx7484), .A (FilterDin_4__4__4)) ;
    oai32 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix533 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx532), .A0 (nx7486), .A1 (
          RST), .A2 (nx8582), .B0 (nx7460), .B1 (nx7488)) ;
    inv01 ix7485 (.Y (nx7486), .A (FilterDin_4__4__5)) ;
    inv01 ix7487 (.Y (nx7488), .A (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx566)) ;
    oai32 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix543 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx542), .A0 (nx7490), .A1 (
          RST), .A2 (nx8582), .B0 (nx7464), .B1 (nx7488)) ;
    inv01 ix7489 (.Y (nx7490), .A (FilterDin_4__4__6)) ;
    oai32 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix553 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx552), .A0 (nx7492), .A1 (
          RST), .A2 (nx8582), .B0 (nx7468), .B1 (nx7488)) ;
    inv01 ix7491 (.Y (nx7492), .A (FilterDin_4__4__7)) ;
    nand02_2x L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix633 (.Y (nx7472), .A0 (
              nx7616), .A1 (nx8582)) ;
    nand02_2x L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix635 (.Y (nx7474), .A0 (
              nx7616), .A1 (nx8582)) ;
    oai32 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix393 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx392), .A0 (nx8742), .A1 (
          RST), .A2 (nx8584), .B0 (nx7402), .B1 (nx7494)) ;
    oai32 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix403 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx402), .A0 (nx8742), .A1 (
          RST), .A2 (nx8584), .B0 (nx7406), .B1 (nx7494)) ;
    oai32 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix413 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx412), .A0 (nx8742), .A1 (
          RST), .A2 (nx8584), .B0 (nx7410), .B1 (nx7494)) ;
    oai32 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix423 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx422), .A0 (nx8742), .A1 (
          RST), .A2 (nx8584), .B0 (nx7414), .B1 (nx7494)) ;
    oai32 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix433 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx432), .A0 (nx8742), .A1 (
          RST), .A2 (nx8584), .B0 (nx7418), .B1 (nx7494)) ;
    oai32 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix443 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx442), .A0 (nx8744), .A1 (
          RST), .A2 (nx8584), .B0 (nx7422), .B1 (nx7494)) ;
    oai32 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix453 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx452), .A0 (nx8744), .A1 (
          RST), .A2 (nx8586), .B0 (nx7426), .B1 (nx7494)) ;
    oai32 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix463 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx462), .A0 (nx8744), .A1 (
          RST), .A2 (nx8586), .B0 (nx7430), .B1 (nx7496)) ;
    oai32 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix473 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx472), .A0 (nx8744), .A1 (
          RST), .A2 (nx8586), .B0 (nx7434), .B1 (nx7496)) ;
    oai32 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix483 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx482), .A0 (nx7476), .A1 (
          RST), .A2 (nx8586), .B0 (nx7438), .B1 (nx7496)) ;
    oai32 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix493 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx492), .A0 (nx7498), .A1 (
          RST), .A2 (nx8586), .B0 (nx7442), .B1 (nx7496)) ;
    inv01 ix7497 (.Y (nx7498), .A (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_10)) ;
    oai32 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix503 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx502), .A0 (nx7500), .A1 (
          RST), .A2 (nx8586), .B0 (nx7446), .B1 (nx7496)) ;
    inv01 ix7499 (.Y (nx7500), .A (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_11)) ;
    oai32 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix513 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx512), .A0 (nx7502), .A1 (
          RST), .A2 (nx8586), .B0 (nx7450), .B1 (nx7496)) ;
    inv01 ix7501 (.Y (nx7502), .A (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_12)) ;
    oai32 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix523 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx522), .A0 (nx7504), .A1 (
          RST), .A2 (nx8588), .B0 (nx7454), .B1 (nx7496)) ;
    inv01 ix7503 (.Y (nx7504), .A (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_13)) ;
    oai32 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix533 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx532), .A0 (nx7506), .A1 (
          RST), .A2 (nx8588), .B0 (nx7458), .B1 (nx7508)) ;
    inv01 ix7505 (.Y (nx7506), .A (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_14)) ;
    inv01 ix7507 (.Y (nx7508), .A (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx566)) ;
    oai32 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix543 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx542), .A0 (nx7510), .A1 (
          RST), .A2 (nx8588), .B0 (nx7462), .B1 (nx7508)) ;
    inv01 ix7509 (.Y (nx7510), .A (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_15)) ;
    oai32 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix553 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_nx552), .A0 (nx7512), .A1 (
          RST), .A2 (nx8588), .B0 (nx7466), .B1 (nx7508)) ;
    inv01 ix7511 (.Y (nx7512), .A (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterSDin_16)) ;
    nand02_2x L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix633 (.Y (nx7494), .A0 (
              nx7616), .A1 (nx8588)) ;
    nand02_2x L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_S_ix635 (.Y (nx7496), .A0 (
              L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx564), .A1 (nx8588)
              ) ;
    oai32 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix393 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx392), .A0 (nx7514), .A1 (
          RST), .A2 (nx8590), .B0 (L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_nx384), .B1 (
          nx7516)) ;
    inv01 ix7513 (.Y (nx7514), .A (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_0)) ;
    oai32 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix403 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx402), .A0 (nx7518), .A1 (
          RST), .A2 (nx8590), .B0 (nx7334), .B1 (nx7516)) ;
    inv01 ix7517 (.Y (nx7518), .A (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_1)) ;
    oai32 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix413 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx412), .A0 (nx7520), .A1 (
          RST), .A2 (nx8590), .B0 (L1_4_L2_4_G5_MINI_ALU_nx387), .B1 (nx7516)) ;
    inv01 ix7519 (.Y (nx7520), .A (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_2)) ;
    oai32 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix423 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx422), .A0 (nx7522), .A1 (
          RST), .A2 (nx8590), .B0 (L1_4_L2_4_G5_MINI_ALU_nx399), .B1 (nx7516)) ;
    inv01 ix7521 (.Y (nx7522), .A (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_3)) ;
    oai32 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix433 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx432), .A0 (nx7524), .A1 (
          RST), .A2 (nx8590), .B0 (L1_4_L2_4_G5_MINI_ALU_nx409), .B1 (nx7516)) ;
    inv01 ix7523 (.Y (nx7524), .A (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_4)) ;
    oai32 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix443 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx442), .A0 (nx7526), .A1 (
          RST), .A2 (nx8590), .B0 (L1_4_L2_4_G5_MINI_ALU_nx419), .B1 (nx7516)) ;
    inv01 ix7525 (.Y (nx7526), .A (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_5)) ;
    oai32 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix453 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx452), .A0 (nx7528), .A1 (
          RST), .A2 (nx8590), .B0 (L1_4_L2_4_G5_MINI_ALU_nx429), .B1 (nx7516)) ;
    inv01 ix7527 (.Y (nx7528), .A (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_6)) ;
    oai32 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix463 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx462), .A0 (nx7530), .A1 (
          RST), .A2 (nx8592), .B0 (L1_4_L2_4_G5_MINI_ALU_nx439), .B1 (nx7532)) ;
    inv01 ix7529 (.Y (nx7530), .A (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_7)) ;
    oai32 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix473 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx472), .A0 (nx7534), .A1 (
          RST), .A2 (nx8592), .B0 (L1_4_L2_4_G5_MINI_ALU_nx449), .B1 (nx7532)) ;
    inv01 ix7533 (.Y (nx7534), .A (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_8)) ;
    oai32 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix483 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx482), .A0 (nx7536), .A1 (
          RST), .A2 (nx8592), .B0 (L1_4_L2_4_G5_MINI_ALU_nx469), .B1 (nx7532)) ;
    inv01 ix7535 (.Y (nx7536), .A (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_9)) ;
    oai32 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix493 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx492), .A0 (nx7538), .A1 (
          RST), .A2 (nx8592), .B0 (L1_4_L2_4_G5_MINI_ALU_nx477), .B1 (nx7532)) ;
    inv01 ix7537 (.Y (nx7538), .A (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_10)) ;
    oai32 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix503 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx502), .A0 (nx7540), .A1 (
          RST), .A2 (nx8592), .B0 (L1_4_L2_4_G5_MINI_ALU_nx485), .B1 (nx7532)) ;
    inv01 ix7539 (.Y (nx7540), .A (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_11)) ;
    oai32 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix513 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx512), .A0 (nx7542), .A1 (
          RST), .A2 (nx8592), .B0 (L1_4_L2_4_G5_MINI_ALU_nx493), .B1 (nx7532)) ;
    inv01 ix7541 (.Y (nx7542), .A (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_12)) ;
    oai32 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix523 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx522), .A0 (nx7544), .A1 (
          RST), .A2 (nx8592), .B0 (L1_4_L2_4_G5_MINI_ALU_nx501), .B1 (nx7532)) ;
    inv01 ix7543 (.Y (nx7544), .A (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_13)) ;
    oai32 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix533 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx532), .A0 (nx7546), .A1 (
          RST), .A2 (nx8594), .B0 (L1_4_L2_4_G5_MINI_ALU_nx509), .B1 (nx7548)) ;
    inv01 ix7545 (.Y (nx7546), .A (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_14)) ;
    inv01 ix7547 (.Y (nx7548), .A (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx566)) ;
    oai32 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix543 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx542), .A0 (nx7550), .A1 (
          RST), .A2 (nx8594), .B0 (L1_4_L2_4_G5_MINI_ALU_nx517), .B1 (nx7548)) ;
    inv01 ix7549 (.Y (nx7550), .A (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_15)) ;
    oai32 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix553 (.Y (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx552), .A0 (nx7552), .A1 (
          RST), .A2 (nx8594), .B0 (nx7350), .B1 (nx7548)) ;
    inv01 ix7551 (.Y (nx7552), .A (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_RegisterPDin_16)) ;
    nand02_2x L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix633 (.Y (nx7516), .A0 (
              L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx564), .A1 (nx8594)
              ) ;
    nand02_2x L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_ix635 (.Y (nx7532), .A0 (
              L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_nx564), .A1 (nx8594)
              ) ;
    inv01 ix7553 (.Y (nx7554), .A (L1_0_L2_0_G1_MINI_ALU_AddPToBoothOperand)) ;
    inv02 ix7555 (.Y (nx7556), .A (nx7554)) ;
    inv02 ix7557 (.Y (nx7558), .A (nx7554)) ;
    inv02 ix7559 (.Y (nx7560), .A (nx7554)) ;
    inv02 ix7561 (.Y (nx7562), .A (L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix7563 (.Y (nx7564), .A (L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix7565 (.Y (nx7566), .A (L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv01 ix7567 (.Y (nx7568), .A (L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx80)) ;
    inv02 ix7569 (.Y (nx7570), .A (nx7568)) ;
    inv02 ix7571 (.Y (nx7572), .A (nx7568)) ;
    inv02 ix7573 (.Y (nx7574), .A (nx7568)) ;
    inv02 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix565_rep_1 (.Y (nx7576), 
          .A (RST)) ;
    inv02 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix565_rep_2 (.Y (nx7578), 
          .A (RST)) ;
    inv02 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix565_rep_3 (.Y (nx7580), 
          .A (RST)) ;
    inv02 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix565_rep_4 (.Y (nx7582), 
          .A (RST)) ;
    inv02 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix565_rep_5 (.Y (nx7584), 
          .A (RST)) ;
    inv02 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix565_rep_6 (.Y (nx7586), 
          .A (RST)) ;
    inv02 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix565_rep_7 (.Y (nx7588), 
          .A (RST)) ;
    inv02 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix565_rep_8 (.Y (nx7590), 
          .A (RST)) ;
    inv02 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix565_rep_9 (.Y (nx7592), 
          .A (RST)) ;
    inv02 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix565_rep_10 (.Y (nx7594)
          , .A (RST)) ;
    inv02 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix565_rep_11 (.Y (nx7596)
          , .A (RST)) ;
    inv02 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix565_rep_12 (.Y (nx7598)
          , .A (RST)) ;
    inv02 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix565_rep_13 (.Y (nx7600)
          , .A (RST)) ;
    inv02 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix565_rep_14 (.Y (nx7602)
          , .A (RST)) ;
    inv02 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix565_rep_15 (.Y (nx7604)
          , .A (RST)) ;
    inv02 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix565_rep_16 (.Y (nx7606)
          , .A (RST)) ;
    inv02 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix565_rep_17 (.Y (nx7608)
          , .A (RST)) ;
    inv02 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix565_rep_18 (.Y (nx7610)
          , .A (RST)) ;
    inv02 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix565_rep_19 (.Y (nx7612)
          , .A (RST)) ;
    inv02 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix565_rep_20 (.Y (nx7614)
          , .A (RST)) ;
    inv02 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_A_ix565_rep_21 (.Y (nx7616)
          , .A (RST)) ;
    inv02 ix7617 (.Y (nx7618), .A (Start)) ;
    inv02 ix7619 (.Y (nx7620), .A (Start)) ;
    inv02 ix7621 (.Y (nx7622), .A (Start)) ;
    inv02 ix7623 (.Y (nx7624), .A (Start)) ;
    inv02 ix7625 (.Y (nx7626), .A (Start)) ;
    inv02 ix7627 (.Y (nx7628), .A (Start)) ;
    inv02 ix7629 (.Y (nx7630), .A (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix7631 (.Y (nx7632), .A (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix7633 (.Y (nx7634), .A (
          L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv01 ix7635 (.Y (nx7636), .A (L1_0_L2_1_G1_MINI_ALU_AddPToBoothOperand)) ;
    inv02 ix7637 (.Y (nx7638), .A (nx7636)) ;
    inv02 ix7639 (.Y (nx7640), .A (nx7636)) ;
    inv02 ix7641 (.Y (nx7642), .A (nx7636)) ;
    inv02 ix7643 (.Y (nx7644), .A (L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix7645 (.Y (nx7646), .A (L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix7647 (.Y (nx7648), .A (L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv01 ix7649 (.Y (nx7650), .A (L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx80)) ;
    inv02 ix7651 (.Y (nx7652), .A (nx7650)) ;
    inv02 ix7653 (.Y (nx7654), .A (nx7650)) ;
    inv02 ix7655 (.Y (nx7656), .A (nx7650)) ;
    inv02 ix7657 (.Y (nx7658), .A (Start)) ;
    inv02 ix7659 (.Y (nx7660), .A (Start)) ;
    inv02 ix7661 (.Y (nx7662), .A (Start)) ;
    inv02 ix7663 (.Y (nx7664), .A (Start)) ;
    inv02 ix7665 (.Y (nx7666), .A (Start)) ;
    inv02 ix7667 (.Y (nx7668), .A (Start)) ;
    inv02 ix7669 (.Y (nx7670), .A (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix7671 (.Y (nx7672), .A (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix7673 (.Y (nx7674), .A (
          L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv01 ix7675 (.Y (nx7676), .A (L1_0_L2_2_G1_MINI_ALU_AddPToBoothOperand)) ;
    inv02 ix7677 (.Y (nx7678), .A (nx7676)) ;
    inv02 ix7679 (.Y (nx7680), .A (nx7676)) ;
    inv02 ix7681 (.Y (nx7682), .A (nx7676)) ;
    inv02 ix7683 (.Y (nx7684), .A (L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix7685 (.Y (nx7686), .A (L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix7687 (.Y (nx7688), .A (L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv01 ix7689 (.Y (nx7690), .A (L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx80)) ;
    inv02 ix7691 (.Y (nx7692), .A (nx7690)) ;
    inv02 ix7693 (.Y (nx7694), .A (nx7690)) ;
    inv02 ix7695 (.Y (nx7696), .A (nx7690)) ;
    inv02 ix7697 (.Y (nx7698), .A (Start)) ;
    inv02 ix7699 (.Y (nx7700), .A (Start)) ;
    inv02 ix7701 (.Y (nx7702), .A (Start)) ;
    inv02 ix7703 (.Y (nx7704), .A (Start)) ;
    inv02 ix7705 (.Y (nx7706), .A (Start)) ;
    inv02 ix7707 (.Y (nx7708), .A (Start)) ;
    inv02 ix7709 (.Y (nx7710), .A (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix7711 (.Y (nx7712), .A (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix7713 (.Y (nx7714), .A (
          L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv01 ix7715 (.Y (nx7716), .A (L1_0_L2_3_G1_MINI_ALU_AddPToBoothOperand)) ;
    inv02 ix7717 (.Y (nx7718), .A (nx7716)) ;
    inv02 ix7719 (.Y (nx7720), .A (nx7716)) ;
    inv02 ix7721 (.Y (nx7722), .A (nx7716)) ;
    inv02 ix7723 (.Y (nx7724), .A (L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix7725 (.Y (nx7726), .A (L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix7727 (.Y (nx7728), .A (L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv01 ix7729 (.Y (nx7730), .A (L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx80)) ;
    inv02 ix7731 (.Y (nx7732), .A (nx7730)) ;
    inv02 ix7733 (.Y (nx7734), .A (nx7730)) ;
    inv02 ix7735 (.Y (nx7736), .A (nx7730)) ;
    inv02 ix7737 (.Y (nx7738), .A (Start)) ;
    inv02 ix7739 (.Y (nx7740), .A (Start)) ;
    inv02 ix7741 (.Y (nx7742), .A (Start)) ;
    inv02 ix7743 (.Y (nx7744), .A (Start)) ;
    inv02 ix7745 (.Y (nx7746), .A (Start)) ;
    inv02 ix7747 (.Y (nx7748), .A (Start)) ;
    inv02 ix7749 (.Y (nx7750), .A (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix7751 (.Y (nx7752), .A (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix7753 (.Y (nx7754), .A (
          L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv01 ix7755 (.Y (nx7756), .A (L1_0_L2_4_G1_MINI_ALU_AddPToBoothOperand)) ;
    inv02 ix7757 (.Y (nx7758), .A (nx7756)) ;
    inv02 ix7759 (.Y (nx7760), .A (nx7756)) ;
    inv02 ix7761 (.Y (nx7762), .A (nx7756)) ;
    inv02 ix7763 (.Y (nx7764), .A (L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix7765 (.Y (nx7766), .A (L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix7767 (.Y (nx7768), .A (L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv01 ix7769 (.Y (nx7770), .A (L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx80)) ;
    inv02 ix7771 (.Y (nx7772), .A (nx7770)) ;
    inv02 ix7773 (.Y (nx7774), .A (nx7770)) ;
    inv02 ix7775 (.Y (nx7776), .A (nx7770)) ;
    inv02 ix7777 (.Y (nx7778), .A (Start)) ;
    inv02 ix7779 (.Y (nx7780), .A (Start)) ;
    inv02 ix7781 (.Y (nx7782), .A (Start)) ;
    inv02 ix7783 (.Y (nx7784), .A (Start)) ;
    inv02 ix7785 (.Y (nx7786), .A (Start)) ;
    inv02 ix7787 (.Y (nx7788), .A (Start)) ;
    inv02 ix7789 (.Y (nx7790), .A (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix7791 (.Y (nx7792), .A (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix7793 (.Y (nx7794), .A (
          L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv01 ix7795 (.Y (nx7796), .A (L1_1_L2_0_G1_MINI_ALU_AddPToBoothOperand)) ;
    inv02 ix7797 (.Y (nx7798), .A (nx7796)) ;
    inv02 ix7799 (.Y (nx7800), .A (nx7796)) ;
    inv02 ix7801 (.Y (nx7802), .A (nx7796)) ;
    inv02 ix7803 (.Y (nx7804), .A (L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix7805 (.Y (nx7806), .A (L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix7807 (.Y (nx7808), .A (L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv01 ix7809 (.Y (nx7810), .A (L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx80)) ;
    inv02 ix7811 (.Y (nx7812), .A (nx7810)) ;
    inv02 ix7813 (.Y (nx7814), .A (nx7810)) ;
    inv02 ix7815 (.Y (nx7816), .A (nx7810)) ;
    inv02 ix7817 (.Y (nx7818), .A (Start)) ;
    inv02 ix7819 (.Y (nx7820), .A (Start)) ;
    inv02 ix7821 (.Y (nx7822), .A (Start)) ;
    inv02 ix7823 (.Y (nx7824), .A (Start)) ;
    inv02 ix7825 (.Y (nx7826), .A (Start)) ;
    inv02 ix7827 (.Y (nx7828), .A (Start)) ;
    inv02 ix7829 (.Y (nx7830), .A (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix7831 (.Y (nx7832), .A (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix7833 (.Y (nx7834), .A (
          L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv01 ix7835 (.Y (nx7836), .A (L1_1_L2_1_G1_MINI_ALU_AddPToBoothOperand)) ;
    inv02 ix7837 (.Y (nx7838), .A (nx7836)) ;
    inv02 ix7839 (.Y (nx7840), .A (nx7836)) ;
    inv02 ix7841 (.Y (nx7842), .A (nx7836)) ;
    inv02 ix7843 (.Y (nx7844), .A (L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix7845 (.Y (nx7846), .A (L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix7847 (.Y (nx7848), .A (L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv01 ix7849 (.Y (nx7850), .A (L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx80)) ;
    inv02 ix7851 (.Y (nx7852), .A (nx7850)) ;
    inv02 ix7853 (.Y (nx7854), .A (nx7850)) ;
    inv02 ix7855 (.Y (nx7856), .A (nx7850)) ;
    inv02 ix7857 (.Y (nx7858), .A (Start)) ;
    inv02 ix7859 (.Y (nx7860), .A (Start)) ;
    inv02 ix7861 (.Y (nx7862), .A (Start)) ;
    inv02 ix7863 (.Y (nx7864), .A (Start)) ;
    inv02 ix7865 (.Y (nx7866), .A (Start)) ;
    inv02 ix7867 (.Y (nx7868), .A (Start)) ;
    inv02 ix7869 (.Y (nx7870), .A (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix7871 (.Y (nx7872), .A (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix7873 (.Y (nx7874), .A (
          L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv01 ix7875 (.Y (nx7876), .A (L1_1_L2_2_G1_MINI_ALU_AddPToBoothOperand)) ;
    inv02 ix7877 (.Y (nx7878), .A (nx7876)) ;
    inv02 ix7879 (.Y (nx7880), .A (nx7876)) ;
    inv02 ix7881 (.Y (nx7882), .A (nx7876)) ;
    inv02 ix7883 (.Y (nx7884), .A (L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix7885 (.Y (nx7886), .A (L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix7887 (.Y (nx7888), .A (L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv01 ix7889 (.Y (nx7890), .A (L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx80)) ;
    inv02 ix7891 (.Y (nx7892), .A (nx7890)) ;
    inv02 ix7893 (.Y (nx7894), .A (nx7890)) ;
    inv02 ix7895 (.Y (nx7896), .A (nx7890)) ;
    inv02 ix7897 (.Y (nx7898), .A (Start)) ;
    inv02 ix7899 (.Y (nx7900), .A (Start)) ;
    inv02 ix7901 (.Y (nx7902), .A (Start)) ;
    inv02 ix7903 (.Y (nx7904), .A (Start)) ;
    inv02 ix7905 (.Y (nx7906), .A (Start)) ;
    inv02 ix7907 (.Y (nx7908), .A (Start)) ;
    inv02 ix7909 (.Y (nx7910), .A (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix7911 (.Y (nx7912), .A (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix7913 (.Y (nx7914), .A (
          L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv01 ix7915 (.Y (nx7916), .A (L1_1_L2_3_G1_MINI_ALU_AddPToBoothOperand)) ;
    inv02 ix7917 (.Y (nx7918), .A (nx7916)) ;
    inv02 ix7919 (.Y (nx7920), .A (nx7916)) ;
    inv02 ix7921 (.Y (nx7922), .A (nx7916)) ;
    inv02 ix7923 (.Y (nx7924), .A (L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix7925 (.Y (nx7926), .A (L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix7927 (.Y (nx7928), .A (L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv01 ix7929 (.Y (nx7930), .A (L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_nx80)) ;
    inv02 ix7931 (.Y (nx7932), .A (nx7930)) ;
    inv02 ix7933 (.Y (nx7934), .A (nx7930)) ;
    inv02 ix7935 (.Y (nx7936), .A (nx7930)) ;
    inv02 ix7937 (.Y (nx7938), .A (Start)) ;
    inv02 ix7939 (.Y (nx7940), .A (Start)) ;
    inv02 ix7941 (.Y (nx7942), .A (Start)) ;
    inv02 ix7943 (.Y (nx7944), .A (Start)) ;
    inv02 ix7945 (.Y (nx7946), .A (Start)) ;
    inv02 ix7947 (.Y (nx7948), .A (Start)) ;
    inv02 ix7949 (.Y (nx7950), .A (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix7951 (.Y (nx7952), .A (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix7953 (.Y (nx7954), .A (
          L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv01 ix7955 (.Y (nx7956), .A (L1_1_L2_4_G1_MINI_ALU_AddPToBoothOperand)) ;
    inv02 ix7957 (.Y (nx7958), .A (nx7956)) ;
    inv02 ix7959 (.Y (nx7960), .A (nx7956)) ;
    inv02 ix7961 (.Y (nx7962), .A (nx7956)) ;
    inv02 ix7963 (.Y (nx7964), .A (L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix7965 (.Y (nx7966), .A (L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix7967 (.Y (nx7968), .A (L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv01 ix7969 (.Y (nx7970), .A (L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_nx80)) ;
    inv02 ix7971 (.Y (nx7972), .A (nx7970)) ;
    inv02 ix7973 (.Y (nx7974), .A (nx7970)) ;
    inv02 ix7975 (.Y (nx7976), .A (nx7970)) ;
    inv02 ix7977 (.Y (nx7978), .A (Start)) ;
    inv02 ix7979 (.Y (nx7980), .A (Start)) ;
    inv02 ix7981 (.Y (nx7982), .A (Start)) ;
    inv02 ix7983 (.Y (nx7984), .A (Start)) ;
    inv02 ix7985 (.Y (nx7986), .A (Start)) ;
    inv02 ix7987 (.Y (nx7988), .A (Start)) ;
    inv02 ix7989 (.Y (nx7990), .A (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix7991 (.Y (nx7992), .A (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix7993 (.Y (nx7994), .A (
          L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv01 ix7995 (.Y (nx7996), .A (L1_2_L2_0_G1_MINI_ALU_AddPToBoothOperand)) ;
    inv02 ix7997 (.Y (nx7998), .A (nx7996)) ;
    inv02 ix7999 (.Y (nx8000), .A (nx7996)) ;
    inv02 ix8001 (.Y (nx8002), .A (nx7996)) ;
    inv02 ix8003 (.Y (nx8004), .A (L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix8005 (.Y (nx8006), .A (L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix8007 (.Y (nx8008), .A (L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv01 ix8009 (.Y (nx8010), .A (L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_nx80)) ;
    inv02 ix8011 (.Y (nx8012), .A (nx8010)) ;
    inv02 ix8013 (.Y (nx8014), .A (nx8010)) ;
    inv02 ix8015 (.Y (nx8016), .A (nx8010)) ;
    inv02 ix8017 (.Y (nx8018), .A (Start)) ;
    inv02 ix8019 (.Y (nx8020), .A (Start)) ;
    inv02 ix8021 (.Y (nx8022), .A (Start)) ;
    inv02 ix8023 (.Y (nx8024), .A (Start)) ;
    inv02 ix8025 (.Y (nx8026), .A (Start)) ;
    inv02 ix8027 (.Y (nx8028), .A (Start)) ;
    inv02 ix8029 (.Y (nx8030), .A (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix8031 (.Y (nx8032), .A (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix8033 (.Y (nx8034), .A (
          L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv01 ix8035 (.Y (nx8036), .A (L1_2_L2_1_G1_MINI_ALU_AddPToBoothOperand)) ;
    inv02 ix8037 (.Y (nx8038), .A (nx8036)) ;
    inv02 ix8039 (.Y (nx8040), .A (nx8036)) ;
    inv02 ix8041 (.Y (nx8042), .A (nx8036)) ;
    inv02 ix8043 (.Y (nx8044), .A (L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix8045 (.Y (nx8046), .A (L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix8047 (.Y (nx8048), .A (L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv01 ix8049 (.Y (nx8050), .A (L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_nx80)) ;
    inv02 ix8051 (.Y (nx8052), .A (nx8050)) ;
    inv02 ix8053 (.Y (nx8054), .A (nx8050)) ;
    inv02 ix8055 (.Y (nx8056), .A (nx8050)) ;
    inv02 ix8057 (.Y (nx8058), .A (Start)) ;
    inv02 ix8059 (.Y (nx8060), .A (Start)) ;
    inv02 ix8061 (.Y (nx8062), .A (Start)) ;
    inv02 ix8063 (.Y (nx8064), .A (Start)) ;
    inv02 ix8065 (.Y (nx8066), .A (Start)) ;
    inv02 ix8067 (.Y (nx8068), .A (Start)) ;
    inv02 ix8069 (.Y (nx8070), .A (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix8071 (.Y (nx8072), .A (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix8073 (.Y (nx8074), .A (
          L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv01 ix8075 (.Y (nx8076), .A (L1_2_L2_2_G1_MINI_ALU_AddPToBoothOperand)) ;
    inv02 ix8077 (.Y (nx8078), .A (nx8076)) ;
    inv02 ix8079 (.Y (nx8080), .A (nx8076)) ;
    inv02 ix8081 (.Y (nx8082), .A (nx8076)) ;
    inv02 ix8083 (.Y (nx8084), .A (L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix8085 (.Y (nx8086), .A (L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix8087 (.Y (nx8088), .A (L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv01 ix8089 (.Y (nx8090), .A (L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_nx80)) ;
    inv02 ix8091 (.Y (nx8092), .A (nx8090)) ;
    inv02 ix8093 (.Y (nx8094), .A (nx8090)) ;
    inv02 ix8095 (.Y (nx8096), .A (nx8090)) ;
    inv02 ix8097 (.Y (nx8098), .A (Start)) ;
    inv02 ix8099 (.Y (nx8100), .A (Start)) ;
    inv02 ix8101 (.Y (nx8102), .A (Start)) ;
    inv02 ix8103 (.Y (nx8104), .A (Start)) ;
    inv02 ix8105 (.Y (nx8106), .A (Start)) ;
    inv02 ix8107 (.Y (nx8108), .A (Start)) ;
    inv02 ix8109 (.Y (nx8110), .A (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix8111 (.Y (nx8112), .A (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix8113 (.Y (nx8114), .A (
          L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv01 ix8115 (.Y (nx8116), .A (L1_2_L2_3_G2_MINI_ALU_AddPToBoothOperand)) ;
    inv02 ix8117 (.Y (nx8118), .A (nx8116)) ;
    inv02 ix8119 (.Y (nx8120), .A (nx8116)) ;
    inv02 ix8121 (.Y (nx8122), .A (nx8116)) ;
    inv02 ix8123 (.Y (nx8124), .A (L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix8125 (.Y (nx8126), .A (L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix8127 (.Y (nx8128), .A (L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv01 ix8129 (.Y (nx8130), .A (L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx80)) ;
    inv02 ix8131 (.Y (nx8132), .A (nx8130)) ;
    inv02 ix8133 (.Y (nx8134), .A (nx8130)) ;
    inv02 ix8135 (.Y (nx8136), .A (nx8130)) ;
    inv02 ix8137 (.Y (nx8138), .A (Start)) ;
    inv02 ix8139 (.Y (nx8140), .A (Start)) ;
    inv02 ix8141 (.Y (nx8142), .A (Start)) ;
    inv02 ix8143 (.Y (nx8144), .A (Start)) ;
    inv02 ix8145 (.Y (nx8146), .A (Start)) ;
    inv02 ix8147 (.Y (nx8148), .A (Start)) ;
    inv02 ix8149 (.Y (nx8150), .A (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix8151 (.Y (nx8152), .A (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix8153 (.Y (nx8154), .A (
          L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv01 ix8155 (.Y (nx8156), .A (L1_2_L2_4_G2_MINI_ALU_AddPToBoothOperand)) ;
    inv02 ix8157 (.Y (nx8158), .A (nx8156)) ;
    inv02 ix8159 (.Y (nx8160), .A (nx8156)) ;
    inv02 ix8161 (.Y (nx8162), .A (nx8156)) ;
    inv02 ix8163 (.Y (nx8164), .A (L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix8165 (.Y (nx8166), .A (L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix8167 (.Y (nx8168), .A (L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv01 ix8169 (.Y (nx8170), .A (L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_nx80)) ;
    inv02 ix8171 (.Y (nx8172), .A (nx8170)) ;
    inv02 ix8173 (.Y (nx8174), .A (nx8170)) ;
    inv02 ix8175 (.Y (nx8176), .A (nx8170)) ;
    inv02 ix8177 (.Y (nx8178), .A (Start)) ;
    inv02 ix8179 (.Y (nx8180), .A (Start)) ;
    inv02 ix8181 (.Y (nx8182), .A (Start)) ;
    inv02 ix8183 (.Y (nx8184), .A (Start)) ;
    inv02 ix8185 (.Y (nx8186), .A (Start)) ;
    inv02 ix8187 (.Y (nx8188), .A (Start)) ;
    inv02 ix8189 (.Y (nx8190), .A (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix8191 (.Y (nx8192), .A (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix8193 (.Y (nx8194), .A (
          L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv01 ix8195 (.Y (nx8196), .A (L1_3_L2_0_G2_MINI_ALU_AddPToBoothOperand)) ;
    inv02 ix8197 (.Y (nx8198), .A (nx8196)) ;
    inv02 ix8199 (.Y (nx8200), .A (nx8196)) ;
    inv02 ix8201 (.Y (nx8202), .A (nx8196)) ;
    inv02 ix8203 (.Y (nx8204), .A (L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix8205 (.Y (nx8206), .A (L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix8207 (.Y (nx8208), .A (L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv01 ix8209 (.Y (nx8210), .A (L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_nx80)) ;
    inv02 ix8211 (.Y (nx8212), .A (nx8210)) ;
    inv02 ix8213 (.Y (nx8214), .A (nx8210)) ;
    inv02 ix8215 (.Y (nx8216), .A (nx8210)) ;
    inv02 ix8217 (.Y (nx8218), .A (Start)) ;
    inv02 ix8219 (.Y (nx8220), .A (Start)) ;
    inv02 ix8221 (.Y (nx8222), .A (Start)) ;
    inv02 ix8223 (.Y (nx8224), .A (Start)) ;
    inv02 ix8225 (.Y (nx8226), .A (Start)) ;
    inv02 ix8227 (.Y (nx8228), .A (Start)) ;
    inv02 ix8229 (.Y (nx8230), .A (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix8231 (.Y (nx8232), .A (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix8233 (.Y (nx8234), .A (
          L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv01 ix8235 (.Y (nx8236), .A (L1_3_L2_1_G2_MINI_ALU_AddPToBoothOperand)) ;
    inv02 ix8237 (.Y (nx8238), .A (nx8236)) ;
    inv02 ix8239 (.Y (nx8240), .A (nx8236)) ;
    inv02 ix8241 (.Y (nx8242), .A (nx8236)) ;
    inv02 ix8243 (.Y (nx8244), .A (L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix8245 (.Y (nx8246), .A (L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix8247 (.Y (nx8248), .A (L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv01 ix8249 (.Y (nx8250), .A (L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_nx80)) ;
    inv02 ix8251 (.Y (nx8252), .A (nx8250)) ;
    inv02 ix8253 (.Y (nx8254), .A (nx8250)) ;
    inv02 ix8255 (.Y (nx8256), .A (nx8250)) ;
    inv02 ix8257 (.Y (nx8258), .A (Start)) ;
    inv02 ix8259 (.Y (nx8260), .A (Start)) ;
    inv02 ix8261 (.Y (nx8262), .A (Start)) ;
    inv02 ix8263 (.Y (nx8264), .A (Start)) ;
    inv02 ix8265 (.Y (nx8266), .A (Start)) ;
    inv02 ix8267 (.Y (nx8268), .A (Start)) ;
    inv02 ix8269 (.Y (nx8270), .A (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix8271 (.Y (nx8272), .A (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix8273 (.Y (nx8274), .A (
          L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv01 ix8275 (.Y (nx8276), .A (L1_3_L2_2_G2_MINI_ALU_AddPToBoothOperand)) ;
    inv02 ix8277 (.Y (nx8278), .A (nx8276)) ;
    inv02 ix8279 (.Y (nx8280), .A (nx8276)) ;
    inv02 ix8281 (.Y (nx8282), .A (nx8276)) ;
    inv02 ix8283 (.Y (nx8284), .A (L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix8285 (.Y (nx8286), .A (L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix8287 (.Y (nx8288), .A (L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv01 ix8289 (.Y (nx8290), .A (L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_nx80)) ;
    inv02 ix8291 (.Y (nx8292), .A (nx8290)) ;
    inv02 ix8293 (.Y (nx8294), .A (nx8290)) ;
    inv02 ix8295 (.Y (nx8296), .A (nx8290)) ;
    inv02 ix8297 (.Y (nx8298), .A (Start)) ;
    inv02 ix8299 (.Y (nx8300), .A (Start)) ;
    inv02 ix8301 (.Y (nx8302), .A (Start)) ;
    inv02 ix8303 (.Y (nx8304), .A (Start)) ;
    inv02 ix8305 (.Y (nx8306), .A (Start)) ;
    inv02 ix8307 (.Y (nx8308), .A (Start)) ;
    inv02 ix8309 (.Y (nx8310), .A (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix8311 (.Y (nx8312), .A (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix8313 (.Y (nx8314), .A (
          L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv01 ix8315 (.Y (nx8316), .A (L1_3_L2_3_G2_MINI_ALU_AddPToBoothOperand)) ;
    inv02 ix8317 (.Y (nx8318), .A (nx8316)) ;
    inv02 ix8319 (.Y (nx8320), .A (nx8316)) ;
    inv02 ix8321 (.Y (nx8322), .A (nx8316)) ;
    inv02 ix8323 (.Y (nx8324), .A (L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix8325 (.Y (nx8326), .A (L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix8327 (.Y (nx8328), .A (L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv01 ix8329 (.Y (nx8330), .A (L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_nx80)) ;
    inv02 ix8331 (.Y (nx8332), .A (nx8330)) ;
    inv02 ix8333 (.Y (nx8334), .A (nx8330)) ;
    inv02 ix8335 (.Y (nx8336), .A (nx8330)) ;
    inv02 ix8337 (.Y (nx8338), .A (Start)) ;
    inv02 ix8339 (.Y (nx8340), .A (Start)) ;
    inv02 ix8341 (.Y (nx8342), .A (Start)) ;
    inv02 ix8343 (.Y (nx8344), .A (Start)) ;
    inv02 ix8345 (.Y (nx8346), .A (Start)) ;
    inv02 ix8347 (.Y (nx8348), .A (Start)) ;
    inv02 ix8349 (.Y (nx8350), .A (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix8351 (.Y (nx8352), .A (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix8353 (.Y (nx8354), .A (
          L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv01 ix8355 (.Y (nx8356), .A (L1_3_L2_4_G3_MINI_ALU_AddPToBoothOperand)) ;
    inv02 ix8357 (.Y (nx8358), .A (nx8356)) ;
    inv02 ix8359 (.Y (nx8360), .A (nx8356)) ;
    inv02 ix8361 (.Y (nx8362), .A (nx8356)) ;
    inv02 ix8363 (.Y (nx8364), .A (L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix8365 (.Y (nx8366), .A (L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix8367 (.Y (nx8368), .A (L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv01 ix8369 (.Y (nx8370), .A (L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_nx80)) ;
    inv02 ix8371 (.Y (nx8372), .A (nx8370)) ;
    inv02 ix8373 (.Y (nx8374), .A (nx8370)) ;
    inv02 ix8375 (.Y (nx8376), .A (nx8370)) ;
    inv02 ix8377 (.Y (nx8378), .A (Start)) ;
    inv02 ix8379 (.Y (nx8380), .A (Start)) ;
    inv02 ix8381 (.Y (nx8382), .A (Start)) ;
    inv02 ix8383 (.Y (nx8384), .A (Start)) ;
    inv02 ix8385 (.Y (nx8386), .A (Start)) ;
    inv02 ix8387 (.Y (nx8388), .A (Start)) ;
    inv02 ix8389 (.Y (nx8390), .A (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix8391 (.Y (nx8392), .A (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix8393 (.Y (nx8394), .A (
          L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv01 ix8395 (.Y (nx8396), .A (L1_4_L2_0_G3_MINI_ALU_AddPToBoothOperand)) ;
    inv02 ix8397 (.Y (nx8398), .A (nx8396)) ;
    inv02 ix8399 (.Y (nx8400), .A (nx8396)) ;
    inv02 ix8401 (.Y (nx8402), .A (nx8396)) ;
    inv02 ix8403 (.Y (nx8404), .A (L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix8405 (.Y (nx8406), .A (L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix8407 (.Y (nx8408), .A (L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv01 ix8409 (.Y (nx8410), .A (L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_nx80)) ;
    inv02 ix8411 (.Y (nx8412), .A (nx8410)) ;
    inv02 ix8413 (.Y (nx8414), .A (nx8410)) ;
    inv02 ix8415 (.Y (nx8416), .A (nx8410)) ;
    inv02 ix8417 (.Y (nx8418), .A (Start)) ;
    inv02 ix8419 (.Y (nx8420), .A (Start)) ;
    inv02 ix8421 (.Y (nx8422), .A (Start)) ;
    inv02 ix8423 (.Y (nx8424), .A (Start)) ;
    inv02 ix8425 (.Y (nx8426), .A (Start)) ;
    inv02 ix8427 (.Y (nx8428), .A (Start)) ;
    inv02 ix8429 (.Y (nx8430), .A (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix8431 (.Y (nx8432), .A (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix8433 (.Y (nx8434), .A (
          L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv01 ix8435 (.Y (nx8436), .A (L1_4_L2_1_G3_MINI_ALU_AddPToBoothOperand)) ;
    inv02 ix8437 (.Y (nx8438), .A (nx8436)) ;
    inv02 ix8439 (.Y (nx8440), .A (nx8436)) ;
    inv02 ix8441 (.Y (nx8442), .A (nx8436)) ;
    inv02 ix8443 (.Y (nx8444), .A (L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix8445 (.Y (nx8446), .A (L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix8447 (.Y (nx8448), .A (L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv01 ix8449 (.Y (nx8450), .A (L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_nx80)) ;
    inv02 ix8451 (.Y (nx8452), .A (nx8450)) ;
    inv02 ix8453 (.Y (nx8454), .A (nx8450)) ;
    inv02 ix8455 (.Y (nx8456), .A (nx8450)) ;
    inv02 ix8457 (.Y (nx8458), .A (Start)) ;
    inv02 ix8459 (.Y (nx8460), .A (Start)) ;
    inv02 ix8461 (.Y (nx8462), .A (Start)) ;
    inv02 ix8463 (.Y (nx8464), .A (Start)) ;
    inv02 ix8465 (.Y (nx8466), .A (Start)) ;
    inv02 ix8467 (.Y (nx8468), .A (Start)) ;
    inv02 ix8469 (.Y (nx8470), .A (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix8471 (.Y (nx8472), .A (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix8473 (.Y (nx8474), .A (
          L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv01 ix8475 (.Y (nx8476), .A (L1_4_L2_2_G4_MINI_ALU_AddPToBoothOperand)) ;
    inv02 ix8477 (.Y (nx8478), .A (nx8476)) ;
    inv02 ix8479 (.Y (nx8480), .A (nx8476)) ;
    inv02 ix8481 (.Y (nx8482), .A (nx8476)) ;
    inv02 ix8483 (.Y (nx8484), .A (L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix8485 (.Y (nx8486), .A (L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix8487 (.Y (nx8488), .A (L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv01 ix8489 (.Y (nx8490), .A (L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_nx80)) ;
    inv02 ix8491 (.Y (nx8492), .A (nx8490)) ;
    inv02 ix8493 (.Y (nx8494), .A (nx8490)) ;
    inv02 ix8495 (.Y (nx8496), .A (nx8490)) ;
    inv02 ix8497 (.Y (nx8498), .A (Start)) ;
    inv02 ix8499 (.Y (nx8500), .A (Start)) ;
    inv02 ix8501 (.Y (nx8502), .A (Start)) ;
    inv02 ix8503 (.Y (nx8504), .A (Start)) ;
    inv02 ix8505 (.Y (nx8506), .A (Start)) ;
    inv02 ix8507 (.Y (nx8508), .A (Start)) ;
    inv02 ix8509 (.Y (nx8510), .A (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix8511 (.Y (nx8512), .A (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix8513 (.Y (nx8514), .A (
          L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv01 ix8515 (.Y (nx8516), .A (L1_4_L2_3_G5_MINI_ALU_AddPToBoothOperand)) ;
    inv02 ix8517 (.Y (nx8518), .A (nx8516)) ;
    inv02 ix8519 (.Y (nx8520), .A (nx8516)) ;
    inv02 ix8521 (.Y (nx8522), .A (nx8516)) ;
    inv02 ix8523 (.Y (nx8524), .A (L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix8525 (.Y (nx8526), .A (L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix8527 (.Y (nx8528), .A (L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv01 ix8529 (.Y (nx8530), .A (L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_nx80)) ;
    inv02 ix8531 (.Y (nx8532), .A (nx8530)) ;
    inv02 ix8533 (.Y (nx8534), .A (nx8530)) ;
    inv02 ix8535 (.Y (nx8536), .A (nx8530)) ;
    inv02 ix8537 (.Y (nx8538), .A (Start)) ;
    inv02 ix8539 (.Y (nx8540), .A (Start)) ;
    inv02 ix8541 (.Y (nx8542), .A (Start)) ;
    inv02 ix8543 (.Y (nx8544), .A (Start)) ;
    inv02 ix8545 (.Y (nx8546), .A (Start)) ;
    inv02 ix8547 (.Y (nx8548), .A (Start)) ;
    inv02 ix8549 (.Y (nx8550), .A (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix8551 (.Y (nx8552), .A (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix8553 (.Y (nx8554), .A (
          L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv01 ix8555 (.Y (nx8556), .A (L1_4_L2_4_G5_MINI_ALU_AddPToBoothOperand)) ;
    inv02 ix8557 (.Y (nx8558), .A (nx8556)) ;
    inv02 ix8559 (.Y (nx8560), .A (nx8556)) ;
    inv02 ix8561 (.Y (nx8562), .A (nx8556)) ;
    inv02 ix8563 (.Y (nx8564), .A (L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix8565 (.Y (nx8566), .A (L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv02 ix8567 (.Y (nx8568), .A (L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_nx384)) ;
    inv01 ix8569 (.Y (nx8570), .A (L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_nx80)) ;
    inv02 ix8571 (.Y (nx8572), .A (nx8570)) ;
    inv02 ix8573 (.Y (nx8574), .A (nx8570)) ;
    inv02 ix8575 (.Y (nx8576), .A (nx8570)) ;
    inv02 ix8577 (.Y (nx8578), .A (Start)) ;
    inv02 ix8579 (.Y (nx8580), .A (Start)) ;
    inv02 ix8581 (.Y (nx8582), .A (Start)) ;
    inv02 ix8583 (.Y (nx8584), .A (Start)) ;
    inv02 ix8585 (.Y (nx8586), .A (Start)) ;
    inv02 ix8587 (.Y (nx8588), .A (Start)) ;
    inv02 ix8589 (.Y (nx8590), .A (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix8591 (.Y (nx8592), .A (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix8593 (.Y (nx8594), .A (
          L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT_REGISTER_P_nx644)) ;
    inv02 ix8595 (.Y (nx8596), .A (
          L1_0_L2_0_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8597 (.Y (nx8598), .A (
          L1_0_L2_0_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8599 (.Y (nx8600), .A (
          L1_0_L2_0_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8601 (.Y (nx8602), .A (
          L1_0_L2_1_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8603 (.Y (nx8604), .A (
          L1_0_L2_1_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8605 (.Y (nx8606), .A (
          L1_0_L2_1_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8607 (.Y (nx8608), .A (
          L1_0_L2_2_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8609 (.Y (nx8610), .A (
          L1_0_L2_2_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8611 (.Y (nx8612), .A (
          L1_0_L2_2_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8613 (.Y (nx8614), .A (
          L1_0_L2_3_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8615 (.Y (nx8616), .A (
          L1_0_L2_3_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8617 (.Y (nx8618), .A (
          L1_0_L2_3_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8619 (.Y (nx8620), .A (
          L1_0_L2_4_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8621 (.Y (nx8622), .A (
          L1_0_L2_4_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8623 (.Y (nx8624), .A (
          L1_0_L2_4_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8625 (.Y (nx8626), .A (
          L1_1_L2_0_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8627 (.Y (nx8628), .A (
          L1_1_L2_0_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8629 (.Y (nx8630), .A (
          L1_1_L2_0_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8631 (.Y (nx8632), .A (
          L1_1_L2_1_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8633 (.Y (nx8634), .A (
          L1_1_L2_1_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8635 (.Y (nx8636), .A (
          L1_1_L2_1_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8637 (.Y (nx8638), .A (
          L1_1_L2_2_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8639 (.Y (nx8640), .A (
          L1_1_L2_2_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8641 (.Y (nx8642), .A (
          L1_1_L2_2_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8643 (.Y (nx8644), .A (
          L1_1_L2_3_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8645 (.Y (nx8646), .A (
          L1_1_L2_3_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8647 (.Y (nx8648), .A (
          L1_1_L2_3_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8649 (.Y (nx8650), .A (
          L1_1_L2_4_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8651 (.Y (nx8652), .A (
          L1_1_L2_4_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8653 (.Y (nx8654), .A (
          L1_1_L2_4_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8655 (.Y (nx8656), .A (
          L1_2_L2_0_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8657 (.Y (nx8658), .A (
          L1_2_L2_0_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8659 (.Y (nx8660), .A (
          L1_2_L2_0_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8661 (.Y (nx8662), .A (
          L1_2_L2_1_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8663 (.Y (nx8664), .A (
          L1_2_L2_1_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8665 (.Y (nx8666), .A (
          L1_2_L2_1_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8667 (.Y (nx8668), .A (
          L1_2_L2_2_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8669 (.Y (nx8670), .A (
          L1_2_L2_2_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8671 (.Y (nx8672), .A (
          L1_2_L2_2_G1_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8673 (.Y (nx8674), .A (
          L1_2_L2_3_G2_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8675 (.Y (nx8676), .A (
          L1_2_L2_3_G2_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8677 (.Y (nx8678), .A (
          L1_2_L2_3_G2_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8679 (.Y (nx8680), .A (
          L1_2_L2_4_G2_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8681 (.Y (nx8682), .A (
          L1_2_L2_4_G2_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8683 (.Y (nx8684), .A (
          L1_2_L2_4_G2_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8685 (.Y (nx8686), .A (
          L1_3_L2_0_G2_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8687 (.Y (nx8688), .A (
          L1_3_L2_0_G2_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8689 (.Y (nx8690), .A (
          L1_3_L2_0_G2_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8691 (.Y (nx8692), .A (
          L1_3_L2_1_G2_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8693 (.Y (nx8694), .A (
          L1_3_L2_1_G2_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8695 (.Y (nx8696), .A (
          L1_3_L2_1_G2_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8697 (.Y (nx8698), .A (
          L1_3_L2_2_G2_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8699 (.Y (nx8700), .A (
          L1_3_L2_2_G2_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8701 (.Y (nx8702), .A (
          L1_3_L2_2_G2_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8703 (.Y (nx8704), .A (
          L1_3_L2_3_G2_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8705 (.Y (nx8706), .A (
          L1_3_L2_3_G2_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8707 (.Y (nx8708), .A (
          L1_3_L2_3_G2_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8709 (.Y (nx8710), .A (
          L1_3_L2_4_G3_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8711 (.Y (nx8712), .A (
          L1_3_L2_4_G3_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8713 (.Y (nx8714), .A (
          L1_3_L2_4_G3_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8715 (.Y (nx8716), .A (
          L1_4_L2_0_G3_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8717 (.Y (nx8718), .A (
          L1_4_L2_0_G3_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8719 (.Y (nx8720), .A (
          L1_4_L2_0_G3_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8721 (.Y (nx8722), .A (
          L1_4_L2_1_G3_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8723 (.Y (nx8724), .A (
          L1_4_L2_1_G3_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8725 (.Y (nx8726), .A (
          L1_4_L2_1_G3_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8727 (.Y (nx8728), .A (
          L1_4_L2_2_G4_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8729 (.Y (nx8730), .A (
          L1_4_L2_2_G4_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8731 (.Y (nx8732), .A (
          L1_4_L2_2_G4_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8733 (.Y (nx8734), .A (
          L1_4_L2_3_G5_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8735 (.Y (nx8736), .A (
          L1_4_L2_3_G5_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8737 (.Y (nx8738), .A (
          L1_4_L2_3_G5_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8739 (.Y (nx8740), .A (
          L1_4_L2_4_G5_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8741 (.Y (nx8742), .A (
          L1_4_L2_4_G5_MINI_ALU_WindowCellShiftedLeft_16)) ;
    inv02 ix8743 (.Y (nx8744), .A (
          L1_4_L2_4_G5_MINI_ALU_WindowCellShiftedLeft_16)) ;
endmodule

