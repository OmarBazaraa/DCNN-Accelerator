//
// Verilog description for cell main, 
// Wed May  9 07:36:13 2018
//
// LeonardoSpectrum Level 3, 2017a.2 
//


module main ( CLK, RST, Start, FilterSize, Stride, Instr, Done ) ;

    input CLK ;
    input RST ;
    input Start ;
    input FilterSize ;
    input Stride ;
    input Instr ;
    output Done ;

    wire FirstCycle, MemWR, MemAddr_17, MemAddr_16, MemAddr_15, MemAddr_14, 
         MemAddr_13, MemAddr_12, MemAddr_11, MemAddr_10, MemAddr_9, MemAddr_8, 
         MemAddr_7, MemAddr_6, MemAddr_5, MemAddr_4, MemAddr_3, MemAddr_2, 
         MemAddr_1, MemAddr_0, MemDin_7, MemDin_6, MemDin_5, MemDin_4, MemDin_3, 
         MemDin_2, MemDin_1, MemDin_0, MemDout_39, MemDout_38, MemDout_37, 
         MemDout_36, MemDout_35, MemDout_34, MemDout_33, MemDout_32, MemDout_31, 
         MemDout_30, MemDout_29, MemDout_28, MemDout_27, MemDout_26, MemDout_25, 
         MemDout_24, MemDout_23, MemDout_22, MemDout_21, MemDout_20, MemDout_19, 
         MemDout_18, MemDout_17, MemDout_16, MemDout_15, MemDout_14, MemDout_13, 
         MemDout_12, MemDout_11, MemDout_10, MemDout_9, MemDout_8, MemDout_7, 
         MemDout_6, MemDout_5, MemDout_4, MemDout_3, MemDout_2, MemDout_1, 
         MemDout_0, CacheRST, CacheFilterWR, CacheWindowWR, CacheFilter_0__0__7, 
         CacheFilter_0__0__6, CacheFilter_0__0__5, CacheFilter_0__0__4, 
         CacheFilter_0__0__3, CacheFilter_0__0__2, CacheFilter_0__0__1, 
         CacheFilter_0__0__0, CacheFilter_0__1__7, CacheFilter_0__1__6, 
         CacheFilter_0__1__5, CacheFilter_0__1__4, CacheFilter_0__1__3, 
         CacheFilter_0__1__2, CacheFilter_0__1__1, CacheFilter_0__1__0, 
         CacheFilter_0__2__7, CacheFilter_0__2__6, CacheFilter_0__2__5, 
         CacheFilter_0__2__4, CacheFilter_0__2__3, CacheFilter_0__2__2, 
         CacheFilter_0__2__1, CacheFilter_0__2__0, CacheFilter_0__3__7, 
         CacheFilter_0__3__6, CacheFilter_0__3__5, CacheFilter_0__3__4, 
         CacheFilter_0__3__3, CacheFilter_0__3__2, CacheFilter_0__3__1, 
         CacheFilter_0__3__0, CacheFilter_0__4__7, CacheFilter_0__4__6, 
         CacheFilter_0__4__5, CacheFilter_0__4__4, CacheFilter_0__4__3, 
         CacheFilter_0__4__2, CacheFilter_0__4__1, CacheFilter_0__4__0, 
         CacheFilter_1__0__7, CacheFilter_1__0__6, CacheFilter_1__0__5, 
         CacheFilter_1__0__4, CacheFilter_1__0__3, CacheFilter_1__0__2, 
         CacheFilter_1__0__1, CacheFilter_1__0__0, CacheFilter_1__1__7, 
         CacheFilter_1__1__6, CacheFilter_1__1__5, CacheFilter_1__1__4, 
         CacheFilter_1__1__3, CacheFilter_1__1__2, CacheFilter_1__1__1, 
         CacheFilter_1__1__0, CacheFilter_1__2__7, CacheFilter_1__2__6, 
         CacheFilter_1__2__5, CacheFilter_1__2__4, CacheFilter_1__2__3, 
         CacheFilter_1__2__2, CacheFilter_1__2__1, CacheFilter_1__2__0, 
         CacheFilter_1__3__7, CacheFilter_1__3__6, CacheFilter_1__3__5, 
         CacheFilter_1__3__4, CacheFilter_1__3__3, CacheFilter_1__3__2, 
         CacheFilter_1__3__1, CacheFilter_1__3__0, CacheFilter_1__4__7, 
         CacheFilter_1__4__6, CacheFilter_1__4__5, CacheFilter_1__4__4, 
         CacheFilter_1__4__3, CacheFilter_1__4__2, CacheFilter_1__4__1, 
         CacheFilter_1__4__0, CacheFilter_2__0__7, CacheFilter_2__0__6, 
         CacheFilter_2__0__5, CacheFilter_2__0__4, CacheFilter_2__0__3, 
         CacheFilter_2__0__2, CacheFilter_2__0__1, CacheFilter_2__0__0, 
         CacheFilter_2__1__7, CacheFilter_2__1__6, CacheFilter_2__1__5, 
         CacheFilter_2__1__4, CacheFilter_2__1__3, CacheFilter_2__1__2, 
         CacheFilter_2__1__1, CacheFilter_2__1__0, CacheFilter_2__2__7, 
         CacheFilter_2__2__6, CacheFilter_2__2__5, CacheFilter_2__2__4, 
         CacheFilter_2__2__3, CacheFilter_2__2__2, CacheFilter_2__2__1, 
         CacheFilter_2__2__0, CacheFilter_2__3__7, CacheFilter_2__3__6, 
         CacheFilter_2__3__5, CacheFilter_2__3__4, CacheFilter_2__3__3, 
         CacheFilter_2__3__2, CacheFilter_2__3__1, CacheFilter_2__3__0, 
         CacheFilter_2__4__7, CacheFilter_2__4__6, CacheFilter_2__4__5, 
         CacheFilter_2__4__4, CacheFilter_2__4__3, CacheFilter_2__4__2, 
         CacheFilter_2__4__1, CacheFilter_2__4__0, CacheFilter_3__0__7, 
         CacheFilter_3__0__6, CacheFilter_3__0__5, CacheFilter_3__0__4, 
         CacheFilter_3__0__3, CacheFilter_3__0__2, CacheFilter_3__0__1, 
         CacheFilter_3__0__0, CacheFilter_3__1__7, CacheFilter_3__1__6, 
         CacheFilter_3__1__5, CacheFilter_3__1__4, CacheFilter_3__1__3, 
         CacheFilter_3__1__2, CacheFilter_3__1__1, CacheFilter_3__1__0, 
         CacheFilter_3__2__7, CacheFilter_3__2__6, CacheFilter_3__2__5, 
         CacheFilter_3__2__4, CacheFilter_3__2__3, CacheFilter_3__2__2, 
         CacheFilter_3__2__1, CacheFilter_3__2__0, CacheFilter_3__3__7, 
         CacheFilter_3__3__6, CacheFilter_3__3__5, CacheFilter_3__3__4, 
         CacheFilter_3__3__3, CacheFilter_3__3__2, CacheFilter_3__3__1, 
         CacheFilter_3__3__0, CacheFilter_3__4__7, CacheFilter_3__4__6, 
         CacheFilter_3__4__5, CacheFilter_3__4__4, CacheFilter_3__4__3, 
         CacheFilter_3__4__2, CacheFilter_3__4__1, CacheFilter_3__4__0, 
         CacheFilter_4__0__7, CacheFilter_4__0__6, CacheFilter_4__0__5, 
         CacheFilter_4__0__4, CacheFilter_4__0__3, CacheFilter_4__0__2, 
         CacheFilter_4__0__1, CacheFilter_4__0__0, CacheFilter_4__1__7, 
         CacheFilter_4__1__6, CacheFilter_4__1__5, CacheFilter_4__1__4, 
         CacheFilter_4__1__3, CacheFilter_4__1__2, CacheFilter_4__1__1, 
         CacheFilter_4__1__0, CacheFilter_4__2__7, CacheFilter_4__2__6, 
         CacheFilter_4__2__5, CacheFilter_4__2__4, CacheFilter_4__2__3, 
         CacheFilter_4__2__2, CacheFilter_4__2__1, CacheFilter_4__2__0, 
         CacheFilter_4__3__7, CacheFilter_4__3__6, CacheFilter_4__3__5, 
         CacheFilter_4__3__4, CacheFilter_4__3__3, CacheFilter_4__3__2, 
         CacheFilter_4__3__1, CacheFilter_4__3__0, CacheFilter_4__4__7, 
         CacheFilter_4__4__6, CacheFilter_4__4__5, CacheFilter_4__4__4, 
         CacheFilter_4__4__3, CacheFilter_4__4__2, CacheFilter_4__4__1, 
         CacheFilter_4__4__0, CacheWindow_0__0__7, CacheWindow_0__0__6, 
         CacheWindow_0__0__5, CacheWindow_0__0__4, CacheWindow_0__0__3, 
         CacheWindow_0__0__2, CacheWindow_0__0__1, CacheWindow_0__0__0, 
         CacheWindow_0__1__7, CacheWindow_0__1__6, CacheWindow_0__1__5, 
         CacheWindow_0__1__4, CacheWindow_0__1__3, CacheWindow_0__1__2, 
         CacheWindow_0__1__1, CacheWindow_0__1__0, CacheWindow_0__2__7, 
         CacheWindow_0__2__6, CacheWindow_0__2__5, CacheWindow_0__2__4, 
         CacheWindow_0__2__3, CacheWindow_0__2__2, CacheWindow_0__2__1, 
         CacheWindow_0__2__0, CacheWindow_0__3__7, CacheWindow_0__3__6, 
         CacheWindow_0__3__5, CacheWindow_0__3__4, CacheWindow_0__3__3, 
         CacheWindow_0__3__2, CacheWindow_0__3__1, CacheWindow_0__3__0, 
         CacheWindow_0__4__7, CacheWindow_0__4__6, CacheWindow_0__4__5, 
         CacheWindow_0__4__4, CacheWindow_0__4__3, CacheWindow_0__4__2, 
         CacheWindow_0__4__1, CacheWindow_0__4__0, CacheWindow_1__0__7, 
         CacheWindow_1__0__6, CacheWindow_1__0__5, CacheWindow_1__0__4, 
         CacheWindow_1__0__3, CacheWindow_1__0__2, CacheWindow_1__0__1, 
         CacheWindow_1__0__0, CacheWindow_1__1__7, CacheWindow_1__1__6, 
         CacheWindow_1__1__5, CacheWindow_1__1__4, CacheWindow_1__1__3, 
         CacheWindow_1__1__2, CacheWindow_1__1__1, CacheWindow_1__1__0, 
         CacheWindow_1__2__7, CacheWindow_1__2__6, CacheWindow_1__2__5, 
         CacheWindow_1__2__4, CacheWindow_1__2__3, CacheWindow_1__2__2, 
         CacheWindow_1__2__1, CacheWindow_1__2__0, CacheWindow_1__3__7, 
         CacheWindow_1__3__6, CacheWindow_1__3__5, CacheWindow_1__3__4, 
         CacheWindow_1__3__3, CacheWindow_1__3__2, CacheWindow_1__3__1, 
         CacheWindow_1__3__0, CacheWindow_1__4__7, CacheWindow_1__4__6, 
         CacheWindow_1__4__5, CacheWindow_1__4__4, CacheWindow_1__4__3, 
         CacheWindow_1__4__2, CacheWindow_1__4__1, CacheWindow_1__4__0, 
         CacheWindow_2__0__7, CacheWindow_2__0__6, CacheWindow_2__0__5, 
         CacheWindow_2__0__4, CacheWindow_2__0__3, CacheWindow_2__0__2, 
         CacheWindow_2__0__1, CacheWindow_2__0__0, CacheWindow_2__1__7, 
         CacheWindow_2__1__6, CacheWindow_2__1__5, CacheWindow_2__1__4, 
         CacheWindow_2__1__3, CacheWindow_2__1__2, CacheWindow_2__1__1, 
         CacheWindow_2__1__0, CacheWindow_2__2__7, CacheWindow_2__2__6, 
         CacheWindow_2__2__5, CacheWindow_2__2__4, CacheWindow_2__2__3, 
         CacheWindow_2__2__2, CacheWindow_2__2__1, CacheWindow_2__2__0, 
         CacheWindow_2__3__7, CacheWindow_2__3__6, CacheWindow_2__3__5, 
         CacheWindow_2__3__4, CacheWindow_2__3__3, CacheWindow_2__3__2, 
         CacheWindow_2__3__1, CacheWindow_2__3__0, CacheWindow_2__4__7, 
         CacheWindow_2__4__6, CacheWindow_2__4__5, CacheWindow_2__4__4, 
         CacheWindow_2__4__3, CacheWindow_2__4__2, CacheWindow_2__4__1, 
         CacheWindow_2__4__0, CacheWindow_3__0__7, CacheWindow_3__0__6, 
         CacheWindow_3__0__5, CacheWindow_3__0__4, CacheWindow_3__0__3, 
         CacheWindow_3__0__2, CacheWindow_3__0__1, CacheWindow_3__0__0, 
         CacheWindow_3__1__7, CacheWindow_3__1__6, CacheWindow_3__1__5, 
         CacheWindow_3__1__4, CacheWindow_3__1__3, CacheWindow_3__1__2, 
         CacheWindow_3__1__1, CacheWindow_3__1__0, CacheWindow_3__2__7, 
         CacheWindow_3__2__6, CacheWindow_3__2__5, CacheWindow_3__2__4, 
         CacheWindow_3__2__3, CacheWindow_3__2__2, CacheWindow_3__2__1, 
         CacheWindow_3__2__0, CacheWindow_3__3__7, CacheWindow_3__3__6, 
         CacheWindow_3__3__5, CacheWindow_3__3__4, CacheWindow_3__3__3, 
         CacheWindow_3__3__2, CacheWindow_3__3__1, CacheWindow_3__3__0, 
         CacheWindow_3__4__7, CacheWindow_3__4__6, CacheWindow_3__4__5, 
         CacheWindow_3__4__4, CacheWindow_3__4__3, CacheWindow_3__4__2, 
         CacheWindow_3__4__1, CacheWindow_3__4__0, CacheWindow_4__0__7, 
         CacheWindow_4__0__6, CacheWindow_4__0__5, CacheWindow_4__0__4, 
         CacheWindow_4__0__3, CacheWindow_4__0__2, CacheWindow_4__0__1, 
         CacheWindow_4__0__0, CacheWindow_4__1__7, CacheWindow_4__1__6, 
         CacheWindow_4__1__5, CacheWindow_4__1__4, CacheWindow_4__1__3, 
         CacheWindow_4__1__2, CacheWindow_4__1__1, CacheWindow_4__1__0, 
         CacheWindow_4__2__7, CacheWindow_4__2__6, CacheWindow_4__2__5, 
         CacheWindow_4__2__4, CacheWindow_4__2__3, CacheWindow_4__2__2, 
         CacheWindow_4__2__1, CacheWindow_4__2__0, CacheWindow_4__3__7, 
         CacheWindow_4__3__6, CacheWindow_4__3__5, CacheWindow_4__3__4, 
         CacheWindow_4__3__3, CacheWindow_4__3__2, CacheWindow_4__3__1, 
         CacheWindow_4__3__0, CacheWindow_4__4__7, CacheWindow_4__4__6, 
         CacheWindow_4__4__5, CacheWindow_4__4__4, CacheWindow_4__4__3, 
         CacheWindow_4__4__2, CacheWindow_4__4__1, CacheWindow_4__4__0, 
         AccStartCalc, AccFinishCalc, AccResult_7, AccResult_6, AccResult_5, 
         AccResult_4, AccResult_3, AccResult_2, AccResult_1, AccResult_0, GND0;
    wire [0:0] \$dummy ;




    controller CONTROLLER (.CLK (CLK), .RST (RST), .Start (Start), .FilterSize (
               FilterSize), .Stride (Stride), .Instr (Instr), .CalcFinished (
               AccFinishCalc), .Calc (AccStartCalc), .MemRD (\$dummy [0]), .MemWR (
               MemWR), .MemAddr ({MemAddr_17,MemAddr_16,MemAddr_15,MemAddr_14,
               MemAddr_13,MemAddr_12,MemAddr_11,MemAddr_10,MemAddr_9,MemAddr_8,
               MemAddr_7,MemAddr_6,MemAddr_5,MemAddr_4,MemAddr_3,MemAddr_2,
               MemAddr_1,MemAddr_0}), .CacheFilterWR (CacheFilterWR), .CacheWindowWR (
               CacheWindowWR), .FirstCycle (FirstCycle), .Done (Done)) ;
    accelerator ACCELERATOR (.CLK (CLK), .RST (RST), .Start (AccStartCalc), .FilterSize (
                FilterSize), .Instr (Instr), .FilterDin_0__0__7 (
                CacheFilter_0__0__7), .FilterDin_0__0__6 (CacheFilter_0__0__6), 
                .FilterDin_0__0__5 (CacheFilter_0__0__5), .FilterDin_0__0__4 (
                CacheFilter_0__0__4), .FilterDin_0__0__3 (CacheFilter_0__0__3), 
                .FilterDin_0__0__2 (CacheFilter_0__0__2), .FilterDin_0__0__1 (
                CacheFilter_0__0__1), .FilterDin_0__0__0 (CacheFilter_0__0__0), 
                .FilterDin_0__1__7 (CacheFilter_0__1__7), .FilterDin_0__1__6 (
                CacheFilter_0__1__6), .FilterDin_0__1__5 (CacheFilter_0__1__5), 
                .FilterDin_0__1__4 (CacheFilter_0__1__4), .FilterDin_0__1__3 (
                CacheFilter_0__1__3), .FilterDin_0__1__2 (CacheFilter_0__1__2), 
                .FilterDin_0__1__1 (CacheFilter_0__1__1), .FilterDin_0__1__0 (
                CacheFilter_0__1__0), .FilterDin_0__2__7 (CacheFilter_0__2__7), 
                .FilterDin_0__2__6 (CacheFilter_0__2__6), .FilterDin_0__2__5 (
                CacheFilter_0__2__5), .FilterDin_0__2__4 (CacheFilter_0__2__4), 
                .FilterDin_0__2__3 (CacheFilter_0__2__3), .FilterDin_0__2__2 (
                CacheFilter_0__2__2), .FilterDin_0__2__1 (CacheFilter_0__2__1), 
                .FilterDin_0__2__0 (CacheFilter_0__2__0), .FilterDin_0__3__7 (
                CacheFilter_0__3__7), .FilterDin_0__3__6 (CacheFilter_0__3__6), 
                .FilterDin_0__3__5 (CacheFilter_0__3__5), .FilterDin_0__3__4 (
                CacheFilter_0__3__4), .FilterDin_0__3__3 (CacheFilter_0__3__3), 
                .FilterDin_0__3__2 (CacheFilter_0__3__2), .FilterDin_0__3__1 (
                CacheFilter_0__3__1), .FilterDin_0__3__0 (CacheFilter_0__3__0), 
                .FilterDin_0__4__7 (CacheFilter_0__4__7), .FilterDin_0__4__6 (
                CacheFilter_0__4__6), .FilterDin_0__4__5 (CacheFilter_0__4__5), 
                .FilterDin_0__4__4 (CacheFilter_0__4__4), .FilterDin_0__4__3 (
                CacheFilter_0__4__3), .FilterDin_0__4__2 (CacheFilter_0__4__2), 
                .FilterDin_0__4__1 (CacheFilter_0__4__1), .FilterDin_0__4__0 (
                CacheFilter_0__4__0), .FilterDin_1__0__7 (CacheFilter_1__0__7), 
                .FilterDin_1__0__6 (CacheFilter_1__0__6), .FilterDin_1__0__5 (
                CacheFilter_1__0__5), .FilterDin_1__0__4 (CacheFilter_1__0__4), 
                .FilterDin_1__0__3 (CacheFilter_1__0__3), .FilterDin_1__0__2 (
                CacheFilter_1__0__2), .FilterDin_1__0__1 (CacheFilter_1__0__1), 
                .FilterDin_1__0__0 (CacheFilter_1__0__0), .FilterDin_1__1__7 (
                CacheFilter_1__1__7), .FilterDin_1__1__6 (CacheFilter_1__1__6), 
                .FilterDin_1__1__5 (CacheFilter_1__1__5), .FilterDin_1__1__4 (
                CacheFilter_1__1__4), .FilterDin_1__1__3 (CacheFilter_1__1__3), 
                .FilterDin_1__1__2 (CacheFilter_1__1__2), .FilterDin_1__1__1 (
                CacheFilter_1__1__1), .FilterDin_1__1__0 (CacheFilter_1__1__0), 
                .FilterDin_1__2__7 (CacheFilter_1__2__7), .FilterDin_1__2__6 (
                CacheFilter_1__2__6), .FilterDin_1__2__5 (CacheFilter_1__2__5), 
                .FilterDin_1__2__4 (CacheFilter_1__2__4), .FilterDin_1__2__3 (
                CacheFilter_1__2__3), .FilterDin_1__2__2 (CacheFilter_1__2__2), 
                .FilterDin_1__2__1 (CacheFilter_1__2__1), .FilterDin_1__2__0 (
                CacheFilter_1__2__0), .FilterDin_1__3__7 (CacheFilter_1__3__7), 
                .FilterDin_1__3__6 (CacheFilter_1__3__6), .FilterDin_1__3__5 (
                CacheFilter_1__3__5), .FilterDin_1__3__4 (CacheFilter_1__3__4), 
                .FilterDin_1__3__3 (CacheFilter_1__3__3), .FilterDin_1__3__2 (
                CacheFilter_1__3__2), .FilterDin_1__3__1 (CacheFilter_1__3__1), 
                .FilterDin_1__3__0 (CacheFilter_1__3__0), .FilterDin_1__4__7 (
                CacheFilter_1__4__7), .FilterDin_1__4__6 (CacheFilter_1__4__6), 
                .FilterDin_1__4__5 (CacheFilter_1__4__5), .FilterDin_1__4__4 (
                CacheFilter_1__4__4), .FilterDin_1__4__3 (CacheFilter_1__4__3), 
                .FilterDin_1__4__2 (CacheFilter_1__4__2), .FilterDin_1__4__1 (
                CacheFilter_1__4__1), .FilterDin_1__4__0 (CacheFilter_1__4__0), 
                .FilterDin_2__0__7 (CacheFilter_2__0__7), .FilterDin_2__0__6 (
                CacheFilter_2__0__6), .FilterDin_2__0__5 (CacheFilter_2__0__5), 
                .FilterDin_2__0__4 (CacheFilter_2__0__4), .FilterDin_2__0__3 (
                CacheFilter_2__0__3), .FilterDin_2__0__2 (CacheFilter_2__0__2), 
                .FilterDin_2__0__1 (CacheFilter_2__0__1), .FilterDin_2__0__0 (
                CacheFilter_2__0__0), .FilterDin_2__1__7 (CacheFilter_2__1__7), 
                .FilterDin_2__1__6 (CacheFilter_2__1__6), .FilterDin_2__1__5 (
                CacheFilter_2__1__5), .FilterDin_2__1__4 (CacheFilter_2__1__4), 
                .FilterDin_2__1__3 (CacheFilter_2__1__3), .FilterDin_2__1__2 (
                CacheFilter_2__1__2), .FilterDin_2__1__1 (CacheFilter_2__1__1), 
                .FilterDin_2__1__0 (CacheFilter_2__1__0), .FilterDin_2__2__7 (
                CacheFilter_2__2__7), .FilterDin_2__2__6 (CacheFilter_2__2__6), 
                .FilterDin_2__2__5 (CacheFilter_2__2__5), .FilterDin_2__2__4 (
                CacheFilter_2__2__4), .FilterDin_2__2__3 (CacheFilter_2__2__3), 
                .FilterDin_2__2__2 (CacheFilter_2__2__2), .FilterDin_2__2__1 (
                CacheFilter_2__2__1), .FilterDin_2__2__0 (CacheFilter_2__2__0), 
                .FilterDin_2__3__7 (CacheFilter_2__3__7), .FilterDin_2__3__6 (
                CacheFilter_2__3__6), .FilterDin_2__3__5 (CacheFilter_2__3__5), 
                .FilterDin_2__3__4 (CacheFilter_2__3__4), .FilterDin_2__3__3 (
                CacheFilter_2__3__3), .FilterDin_2__3__2 (CacheFilter_2__3__2), 
                .FilterDin_2__3__1 (CacheFilter_2__3__1), .FilterDin_2__3__0 (
                CacheFilter_2__3__0), .FilterDin_2__4__7 (CacheFilter_2__4__7), 
                .FilterDin_2__4__6 (CacheFilter_2__4__6), .FilterDin_2__4__5 (
                CacheFilter_2__4__5), .FilterDin_2__4__4 (CacheFilter_2__4__4), 
                .FilterDin_2__4__3 (CacheFilter_2__4__3), .FilterDin_2__4__2 (
                CacheFilter_2__4__2), .FilterDin_2__4__1 (CacheFilter_2__4__1), 
                .FilterDin_2__4__0 (CacheFilter_2__4__0), .FilterDin_3__0__7 (
                CacheFilter_3__0__7), .FilterDin_3__0__6 (CacheFilter_3__0__6), 
                .FilterDin_3__0__5 (CacheFilter_3__0__5), .FilterDin_3__0__4 (
                CacheFilter_3__0__4), .FilterDin_3__0__3 (CacheFilter_3__0__3), 
                .FilterDin_3__0__2 (CacheFilter_3__0__2), .FilterDin_3__0__1 (
                CacheFilter_3__0__1), .FilterDin_3__0__0 (CacheFilter_3__0__0), 
                .FilterDin_3__1__7 (CacheFilter_3__1__7), .FilterDin_3__1__6 (
                CacheFilter_3__1__6), .FilterDin_3__1__5 (CacheFilter_3__1__5), 
                .FilterDin_3__1__4 (CacheFilter_3__1__4), .FilterDin_3__1__3 (
                CacheFilter_3__1__3), .FilterDin_3__1__2 (CacheFilter_3__1__2), 
                .FilterDin_3__1__1 (CacheFilter_3__1__1), .FilterDin_3__1__0 (
                CacheFilter_3__1__0), .FilterDin_3__2__7 (CacheFilter_3__2__7), 
                .FilterDin_3__2__6 (CacheFilter_3__2__6), .FilterDin_3__2__5 (
                CacheFilter_3__2__5), .FilterDin_3__2__4 (CacheFilter_3__2__4), 
                .FilterDin_3__2__3 (CacheFilter_3__2__3), .FilterDin_3__2__2 (
                CacheFilter_3__2__2), .FilterDin_3__2__1 (CacheFilter_3__2__1), 
                .FilterDin_3__2__0 (CacheFilter_3__2__0), .FilterDin_3__3__7 (
                CacheFilter_3__3__7), .FilterDin_3__3__6 (CacheFilter_3__3__6), 
                .FilterDin_3__3__5 (CacheFilter_3__3__5), .FilterDin_3__3__4 (
                CacheFilter_3__3__4), .FilterDin_3__3__3 (CacheFilter_3__3__3), 
                .FilterDin_3__3__2 (CacheFilter_3__3__2), .FilterDin_3__3__1 (
                CacheFilter_3__3__1), .FilterDin_3__3__0 (CacheFilter_3__3__0), 
                .FilterDin_3__4__7 (CacheFilter_3__4__7), .FilterDin_3__4__6 (
                CacheFilter_3__4__6), .FilterDin_3__4__5 (CacheFilter_3__4__5), 
                .FilterDin_3__4__4 (CacheFilter_3__4__4), .FilterDin_3__4__3 (
                CacheFilter_3__4__3), .FilterDin_3__4__2 (CacheFilter_3__4__2), 
                .FilterDin_3__4__1 (CacheFilter_3__4__1), .FilterDin_3__4__0 (
                CacheFilter_3__4__0), .FilterDin_4__0__7 (CacheFilter_4__0__7), 
                .FilterDin_4__0__6 (CacheFilter_4__0__6), .FilterDin_4__0__5 (
                CacheFilter_4__0__5), .FilterDin_4__0__4 (CacheFilter_4__0__4), 
                .FilterDin_4__0__3 (CacheFilter_4__0__3), .FilterDin_4__0__2 (
                CacheFilter_4__0__2), .FilterDin_4__0__1 (CacheFilter_4__0__1), 
                .FilterDin_4__0__0 (CacheFilter_4__0__0), .FilterDin_4__1__7 (
                CacheFilter_4__1__7), .FilterDin_4__1__6 (CacheFilter_4__1__6), 
                .FilterDin_4__1__5 (CacheFilter_4__1__5), .FilterDin_4__1__4 (
                CacheFilter_4__1__4), .FilterDin_4__1__3 (CacheFilter_4__1__3), 
                .FilterDin_4__1__2 (CacheFilter_4__1__2), .FilterDin_4__1__1 (
                CacheFilter_4__1__1), .FilterDin_4__1__0 (CacheFilter_4__1__0), 
                .FilterDin_4__2__7 (CacheFilter_4__2__7), .FilterDin_4__2__6 (
                CacheFilter_4__2__6), .FilterDin_4__2__5 (CacheFilter_4__2__5), 
                .FilterDin_4__2__4 (CacheFilter_4__2__4), .FilterDin_4__2__3 (
                CacheFilter_4__2__3), .FilterDin_4__2__2 (CacheFilter_4__2__2), 
                .FilterDin_4__2__1 (CacheFilter_4__2__1), .FilterDin_4__2__0 (
                CacheFilter_4__2__0), .FilterDin_4__3__7 (CacheFilter_4__3__7), 
                .FilterDin_4__3__6 (CacheFilter_4__3__6), .FilterDin_4__3__5 (
                CacheFilter_4__3__5), .FilterDin_4__3__4 (CacheFilter_4__3__4), 
                .FilterDin_4__3__3 (CacheFilter_4__3__3), .FilterDin_4__3__2 (
                CacheFilter_4__3__2), .FilterDin_4__3__1 (CacheFilter_4__3__1), 
                .FilterDin_4__3__0 (CacheFilter_4__3__0), .FilterDin_4__4__7 (
                CacheFilter_4__4__7), .FilterDin_4__4__6 (CacheFilter_4__4__6), 
                .FilterDin_4__4__5 (CacheFilter_4__4__5), .FilterDin_4__4__4 (
                CacheFilter_4__4__4), .FilterDin_4__4__3 (CacheFilter_4__4__3), 
                .FilterDin_4__4__2 (CacheFilter_4__4__2), .FilterDin_4__4__1 (
                CacheFilter_4__4__1), .FilterDin_4__4__0 (CacheFilter_4__4__0), 
                .WindowDin_0__0__7 (CacheWindow_0__0__7), .WindowDin_0__0__6 (
                CacheWindow_0__0__6), .WindowDin_0__0__5 (CacheWindow_0__0__5), 
                .WindowDin_0__0__4 (CacheWindow_0__0__4), .WindowDin_0__0__3 (
                CacheWindow_0__0__3), .WindowDin_0__0__2 (CacheWindow_0__0__2), 
                .WindowDin_0__0__1 (CacheWindow_0__0__1), .WindowDin_0__0__0 (
                CacheWindow_0__0__0), .WindowDin_0__1__7 (CacheWindow_0__1__7), 
                .WindowDin_0__1__6 (CacheWindow_0__1__6), .WindowDin_0__1__5 (
                CacheWindow_0__1__5), .WindowDin_0__1__4 (CacheWindow_0__1__4), 
                .WindowDin_0__1__3 (CacheWindow_0__1__3), .WindowDin_0__1__2 (
                CacheWindow_0__1__2), .WindowDin_0__1__1 (CacheWindow_0__1__1), 
                .WindowDin_0__1__0 (CacheWindow_0__1__0), .WindowDin_0__2__7 (
                CacheWindow_0__2__7), .WindowDin_0__2__6 (CacheWindow_0__2__6), 
                .WindowDin_0__2__5 (CacheWindow_0__2__5), .WindowDin_0__2__4 (
                CacheWindow_0__2__4), .WindowDin_0__2__3 (CacheWindow_0__2__3), 
                .WindowDin_0__2__2 (CacheWindow_0__2__2), .WindowDin_0__2__1 (
                CacheWindow_0__2__1), .WindowDin_0__2__0 (CacheWindow_0__2__0), 
                .WindowDin_0__3__7 (CacheWindow_0__3__7), .WindowDin_0__3__6 (
                CacheWindow_0__3__6), .WindowDin_0__3__5 (CacheWindow_0__3__5), 
                .WindowDin_0__3__4 (CacheWindow_0__3__4), .WindowDin_0__3__3 (
                CacheWindow_0__3__3), .WindowDin_0__3__2 (CacheWindow_0__3__2), 
                .WindowDin_0__3__1 (CacheWindow_0__3__1), .WindowDin_0__3__0 (
                CacheWindow_0__3__0), .WindowDin_0__4__7 (CacheWindow_0__4__7), 
                .WindowDin_0__4__6 (CacheWindow_0__4__6), .WindowDin_0__4__5 (
                CacheWindow_0__4__5), .WindowDin_0__4__4 (CacheWindow_0__4__4), 
                .WindowDin_0__4__3 (CacheWindow_0__4__3), .WindowDin_0__4__2 (
                CacheWindow_0__4__2), .WindowDin_0__4__1 (CacheWindow_0__4__1), 
                .WindowDin_0__4__0 (CacheWindow_0__4__0), .WindowDin_1__0__7 (
                CacheWindow_1__0__7), .WindowDin_1__0__6 (CacheWindow_1__0__6), 
                .WindowDin_1__0__5 (CacheWindow_1__0__5), .WindowDin_1__0__4 (
                CacheWindow_1__0__4), .WindowDin_1__0__3 (CacheWindow_1__0__3), 
                .WindowDin_1__0__2 (CacheWindow_1__0__2), .WindowDin_1__0__1 (
                CacheWindow_1__0__1), .WindowDin_1__0__0 (CacheWindow_1__0__0), 
                .WindowDin_1__1__7 (CacheWindow_1__1__7), .WindowDin_1__1__6 (
                CacheWindow_1__1__6), .WindowDin_1__1__5 (CacheWindow_1__1__5), 
                .WindowDin_1__1__4 (CacheWindow_1__1__4), .WindowDin_1__1__3 (
                CacheWindow_1__1__3), .WindowDin_1__1__2 (CacheWindow_1__1__2), 
                .WindowDin_1__1__1 (CacheWindow_1__1__1), .WindowDin_1__1__0 (
                CacheWindow_1__1__0), .WindowDin_1__2__7 (CacheWindow_1__2__7), 
                .WindowDin_1__2__6 (CacheWindow_1__2__6), .WindowDin_1__2__5 (
                CacheWindow_1__2__5), .WindowDin_1__2__4 (CacheWindow_1__2__4), 
                .WindowDin_1__2__3 (CacheWindow_1__2__3), .WindowDin_1__2__2 (
                CacheWindow_1__2__2), .WindowDin_1__2__1 (CacheWindow_1__2__1), 
                .WindowDin_1__2__0 (CacheWindow_1__2__0), .WindowDin_1__3__7 (
                CacheWindow_1__3__7), .WindowDin_1__3__6 (CacheWindow_1__3__6), 
                .WindowDin_1__3__5 (CacheWindow_1__3__5), .WindowDin_1__3__4 (
                CacheWindow_1__3__4), .WindowDin_1__3__3 (CacheWindow_1__3__3), 
                .WindowDin_1__3__2 (CacheWindow_1__3__2), .WindowDin_1__3__1 (
                CacheWindow_1__3__1), .WindowDin_1__3__0 (CacheWindow_1__3__0), 
                .WindowDin_1__4__7 (CacheWindow_1__4__7), .WindowDin_1__4__6 (
                CacheWindow_1__4__6), .WindowDin_1__4__5 (CacheWindow_1__4__5), 
                .WindowDin_1__4__4 (CacheWindow_1__4__4), .WindowDin_1__4__3 (
                CacheWindow_1__4__3), .WindowDin_1__4__2 (CacheWindow_1__4__2), 
                .WindowDin_1__4__1 (CacheWindow_1__4__1), .WindowDin_1__4__0 (
                CacheWindow_1__4__0), .WindowDin_2__0__7 (CacheWindow_2__0__7), 
                .WindowDin_2__0__6 (CacheWindow_2__0__6), .WindowDin_2__0__5 (
                CacheWindow_2__0__5), .WindowDin_2__0__4 (CacheWindow_2__0__4), 
                .WindowDin_2__0__3 (CacheWindow_2__0__3), .WindowDin_2__0__2 (
                CacheWindow_2__0__2), .WindowDin_2__0__1 (CacheWindow_2__0__1), 
                .WindowDin_2__0__0 (CacheWindow_2__0__0), .WindowDin_2__1__7 (
                CacheWindow_2__1__7), .WindowDin_2__1__6 (CacheWindow_2__1__6), 
                .WindowDin_2__1__5 (CacheWindow_2__1__5), .WindowDin_2__1__4 (
                CacheWindow_2__1__4), .WindowDin_2__1__3 (CacheWindow_2__1__3), 
                .WindowDin_2__1__2 (CacheWindow_2__1__2), .WindowDin_2__1__1 (
                CacheWindow_2__1__1), .WindowDin_2__1__0 (CacheWindow_2__1__0), 
                .WindowDin_2__2__7 (CacheWindow_2__2__7), .WindowDin_2__2__6 (
                CacheWindow_2__2__6), .WindowDin_2__2__5 (CacheWindow_2__2__5), 
                .WindowDin_2__2__4 (CacheWindow_2__2__4), .WindowDin_2__2__3 (
                CacheWindow_2__2__3), .WindowDin_2__2__2 (CacheWindow_2__2__2), 
                .WindowDin_2__2__1 (CacheWindow_2__2__1), .WindowDin_2__2__0 (
                CacheWindow_2__2__0), .WindowDin_2__3__7 (CacheWindow_2__3__7), 
                .WindowDin_2__3__6 (CacheWindow_2__3__6), .WindowDin_2__3__5 (
                CacheWindow_2__3__5), .WindowDin_2__3__4 (CacheWindow_2__3__4), 
                .WindowDin_2__3__3 (CacheWindow_2__3__3), .WindowDin_2__3__2 (
                CacheWindow_2__3__2), .WindowDin_2__3__1 (CacheWindow_2__3__1), 
                .WindowDin_2__3__0 (CacheWindow_2__3__0), .WindowDin_2__4__7 (
                CacheWindow_2__4__7), .WindowDin_2__4__6 (CacheWindow_2__4__6), 
                .WindowDin_2__4__5 (CacheWindow_2__4__5), .WindowDin_2__4__4 (
                CacheWindow_2__4__4), .WindowDin_2__4__3 (CacheWindow_2__4__3), 
                .WindowDin_2__4__2 (CacheWindow_2__4__2), .WindowDin_2__4__1 (
                CacheWindow_2__4__1), .WindowDin_2__4__0 (CacheWindow_2__4__0), 
                .WindowDin_3__0__7 (CacheWindow_3__0__7), .WindowDin_3__0__6 (
                CacheWindow_3__0__6), .WindowDin_3__0__5 (CacheWindow_3__0__5), 
                .WindowDin_3__0__4 (CacheWindow_3__0__4), .WindowDin_3__0__3 (
                CacheWindow_3__0__3), .WindowDin_3__0__2 (CacheWindow_3__0__2), 
                .WindowDin_3__0__1 (CacheWindow_3__0__1), .WindowDin_3__0__0 (
                CacheWindow_3__0__0), .WindowDin_3__1__7 (CacheWindow_3__1__7), 
                .WindowDin_3__1__6 (CacheWindow_3__1__6), .WindowDin_3__1__5 (
                CacheWindow_3__1__5), .WindowDin_3__1__4 (CacheWindow_3__1__4), 
                .WindowDin_3__1__3 (CacheWindow_3__1__3), .WindowDin_3__1__2 (
                CacheWindow_3__1__2), .WindowDin_3__1__1 (CacheWindow_3__1__1), 
                .WindowDin_3__1__0 (CacheWindow_3__1__0), .WindowDin_3__2__7 (
                CacheWindow_3__2__7), .WindowDin_3__2__6 (CacheWindow_3__2__6), 
                .WindowDin_3__2__5 (CacheWindow_3__2__5), .WindowDin_3__2__4 (
                CacheWindow_3__2__4), .WindowDin_3__2__3 (CacheWindow_3__2__3), 
                .WindowDin_3__2__2 (CacheWindow_3__2__2), .WindowDin_3__2__1 (
                CacheWindow_3__2__1), .WindowDin_3__2__0 (CacheWindow_3__2__0), 
                .WindowDin_3__3__7 (CacheWindow_3__3__7), .WindowDin_3__3__6 (
                CacheWindow_3__3__6), .WindowDin_3__3__5 (CacheWindow_3__3__5), 
                .WindowDin_3__3__4 (CacheWindow_3__3__4), .WindowDin_3__3__3 (
                CacheWindow_3__3__3), .WindowDin_3__3__2 (CacheWindow_3__3__2), 
                .WindowDin_3__3__1 (CacheWindow_3__3__1), .WindowDin_3__3__0 (
                CacheWindow_3__3__0), .WindowDin_3__4__7 (CacheWindow_3__4__7), 
                .WindowDin_3__4__6 (CacheWindow_3__4__6), .WindowDin_3__4__5 (
                CacheWindow_3__4__5), .WindowDin_3__4__4 (CacheWindow_3__4__4), 
                .WindowDin_3__4__3 (CacheWindow_3__4__3), .WindowDin_3__4__2 (
                CacheWindow_3__4__2), .WindowDin_3__4__1 (CacheWindow_3__4__1), 
                .WindowDin_3__4__0 (CacheWindow_3__4__0), .WindowDin_4__0__7 (
                CacheWindow_4__0__7), .WindowDin_4__0__6 (CacheWindow_4__0__6), 
                .WindowDin_4__0__5 (CacheWindow_4__0__5), .WindowDin_4__0__4 (
                CacheWindow_4__0__4), .WindowDin_4__0__3 (CacheWindow_4__0__3), 
                .WindowDin_4__0__2 (CacheWindow_4__0__2), .WindowDin_4__0__1 (
                CacheWindow_4__0__1), .WindowDin_4__0__0 (CacheWindow_4__0__0), 
                .WindowDin_4__1__7 (CacheWindow_4__1__7), .WindowDin_4__1__6 (
                CacheWindow_4__1__6), .WindowDin_4__1__5 (CacheWindow_4__1__5), 
                .WindowDin_4__1__4 (CacheWindow_4__1__4), .WindowDin_4__1__3 (
                CacheWindow_4__1__3), .WindowDin_4__1__2 (CacheWindow_4__1__2), 
                .WindowDin_4__1__1 (CacheWindow_4__1__1), .WindowDin_4__1__0 (
                CacheWindow_4__1__0), .WindowDin_4__2__7 (CacheWindow_4__2__7), 
                .WindowDin_4__2__6 (CacheWindow_4__2__6), .WindowDin_4__2__5 (
                CacheWindow_4__2__5), .WindowDin_4__2__4 (CacheWindow_4__2__4), 
                .WindowDin_4__2__3 (CacheWindow_4__2__3), .WindowDin_4__2__2 (
                CacheWindow_4__2__2), .WindowDin_4__2__1 (CacheWindow_4__2__1), 
                .WindowDin_4__2__0 (CacheWindow_4__2__0), .WindowDin_4__3__7 (
                CacheWindow_4__3__7), .WindowDin_4__3__6 (CacheWindow_4__3__6), 
                .WindowDin_4__3__5 (CacheWindow_4__3__5), .WindowDin_4__3__4 (
                CacheWindow_4__3__4), .WindowDin_4__3__3 (CacheWindow_4__3__3), 
                .WindowDin_4__3__2 (CacheWindow_4__3__2), .WindowDin_4__3__1 (
                CacheWindow_4__3__1), .WindowDin_4__3__0 (CacheWindow_4__3__0), 
                .WindowDin_4__4__7 (CacheWindow_4__4__7), .WindowDin_4__4__6 (
                CacheWindow_4__4__6), .WindowDin_4__4__5 (CacheWindow_4__4__5), 
                .WindowDin_4__4__4 (CacheWindow_4__4__4), .WindowDin_4__4__3 (
                CacheWindow_4__4__3), .WindowDin_4__4__2 (CacheWindow_4__4__2), 
                .WindowDin_4__4__1 (CacheWindow_4__4__1), .WindowDin_4__4__0 (
                CacheWindow_4__4__0), .Done (AccFinishCalc), .Result ({
                AccResult_7,AccResult_6,AccResult_5,AccResult_4,AccResult_3,
                AccResult_2,AccResult_1,AccResult_0})) ;
    RAM_8_18 RAM (.CLK (CLK), .WR (MemWR), .Address ({MemAddr_17,MemAddr_16,
             MemAddr_15,MemAddr_14,MemAddr_13,MemAddr_12,MemAddr_11,MemAddr_10,
             MemAddr_9,MemAddr_8,MemAddr_7,MemAddr_6,MemAddr_5,MemAddr_4,
             MemAddr_3,MemAddr_2,MemAddr_1,MemAddr_0}), .Din ({MemDin_7,MemDin_6
             ,MemDin_5,MemDin_4,MemDin_3,MemDin_2,MemDin_1,MemDin_0}), .Dout ({
             MemDout_39,MemDout_38,MemDout_37,MemDout_36,MemDout_35,MemDout_34,
             MemDout_33,MemDout_32,MemDout_31,MemDout_30,MemDout_29,MemDout_28,
             MemDout_27,MemDout_26,MemDout_25,MemDout_24,MemDout_23,MemDout_22,
             MemDout_21,MemDout_20,MemDout_19,MemDout_18,MemDout_17,MemDout_16,
             MemDout_15,MemDout_14,MemDout_13,MemDout_12,MemDout_11,MemDout_10,
             MemDout_9,MemDout_8,MemDout_7,MemDout_6,MemDout_5,MemDout_4,
             MemDout_3,MemDout_2,MemDout_1,MemDout_0})) ;
    or (CacheRST, RST, FirstCycle) ;
    cache CACHE (.CLK (CLK), .RST (CacheRST), .FilterSize (FilterSize), .FilterWR (
          CacheFilterWR), .WindowWR (CacheWindowWR), .Din ({MemDout_39,
          MemDout_38,MemDout_37,MemDout_36,MemDout_35,MemDout_34,MemDout_33,
          MemDout_32,MemDout_31,MemDout_30,MemDout_29,MemDout_28,MemDout_27,
          MemDout_26,MemDout_25,MemDout_24,MemDout_23,MemDout_22,MemDout_21,
          MemDout_20,MemDout_19,MemDout_18,MemDout_17,MemDout_16,MemDout_15,
          MemDout_14,MemDout_13,MemDout_12,MemDout_11,MemDout_10,MemDout_9,
          MemDout_8,MemDout_7,MemDout_6,MemDout_5,MemDout_4,MemDout_3,MemDout_2,
          MemDout_1,MemDout_0}), .FilterDout_0__0__7 (CacheFilter_0__0__7), .FilterDout_0__0__6 (
          CacheFilter_0__0__6), .FilterDout_0__0__5 (CacheFilter_0__0__5), .FilterDout_0__0__4 (
          CacheFilter_0__0__4), .FilterDout_0__0__3 (CacheFilter_0__0__3), .FilterDout_0__0__2 (
          CacheFilter_0__0__2), .FilterDout_0__0__1 (CacheFilter_0__0__1), .FilterDout_0__0__0 (
          CacheFilter_0__0__0), .FilterDout_0__1__7 (CacheFilter_0__1__7), .FilterDout_0__1__6 (
          CacheFilter_0__1__6), .FilterDout_0__1__5 (CacheFilter_0__1__5), .FilterDout_0__1__4 (
          CacheFilter_0__1__4), .FilterDout_0__1__3 (CacheFilter_0__1__3), .FilterDout_0__1__2 (
          CacheFilter_0__1__2), .FilterDout_0__1__1 (CacheFilter_0__1__1), .FilterDout_0__1__0 (
          CacheFilter_0__1__0), .FilterDout_0__2__7 (CacheFilter_0__2__7), .FilterDout_0__2__6 (
          CacheFilter_0__2__6), .FilterDout_0__2__5 (CacheFilter_0__2__5), .FilterDout_0__2__4 (
          CacheFilter_0__2__4), .FilterDout_0__2__3 (CacheFilter_0__2__3), .FilterDout_0__2__2 (
          CacheFilter_0__2__2), .FilterDout_0__2__1 (CacheFilter_0__2__1), .FilterDout_0__2__0 (
          CacheFilter_0__2__0), .FilterDout_0__3__7 (CacheFilter_0__3__7), .FilterDout_0__3__6 (
          CacheFilter_0__3__6), .FilterDout_0__3__5 (CacheFilter_0__3__5), .FilterDout_0__3__4 (
          CacheFilter_0__3__4), .FilterDout_0__3__3 (CacheFilter_0__3__3), .FilterDout_0__3__2 (
          CacheFilter_0__3__2), .FilterDout_0__3__1 (CacheFilter_0__3__1), .FilterDout_0__3__0 (
          CacheFilter_0__3__0), .FilterDout_0__4__7 (CacheFilter_0__4__7), .FilterDout_0__4__6 (
          CacheFilter_0__4__6), .FilterDout_0__4__5 (CacheFilter_0__4__5), .FilterDout_0__4__4 (
          CacheFilter_0__4__4), .FilterDout_0__4__3 (CacheFilter_0__4__3), .FilterDout_0__4__2 (
          CacheFilter_0__4__2), .FilterDout_0__4__1 (CacheFilter_0__4__1), .FilterDout_0__4__0 (
          CacheFilter_0__4__0), .FilterDout_1__0__7 (CacheFilter_1__0__7), .FilterDout_1__0__6 (
          CacheFilter_1__0__6), .FilterDout_1__0__5 (CacheFilter_1__0__5), .FilterDout_1__0__4 (
          CacheFilter_1__0__4), .FilterDout_1__0__3 (CacheFilter_1__0__3), .FilterDout_1__0__2 (
          CacheFilter_1__0__2), .FilterDout_1__0__1 (CacheFilter_1__0__1), .FilterDout_1__0__0 (
          CacheFilter_1__0__0), .FilterDout_1__1__7 (CacheFilter_1__1__7), .FilterDout_1__1__6 (
          CacheFilter_1__1__6), .FilterDout_1__1__5 (CacheFilter_1__1__5), .FilterDout_1__1__4 (
          CacheFilter_1__1__4), .FilterDout_1__1__3 (CacheFilter_1__1__3), .FilterDout_1__1__2 (
          CacheFilter_1__1__2), .FilterDout_1__1__1 (CacheFilter_1__1__1), .FilterDout_1__1__0 (
          CacheFilter_1__1__0), .FilterDout_1__2__7 (CacheFilter_1__2__7), .FilterDout_1__2__6 (
          CacheFilter_1__2__6), .FilterDout_1__2__5 (CacheFilter_1__2__5), .FilterDout_1__2__4 (
          CacheFilter_1__2__4), .FilterDout_1__2__3 (CacheFilter_1__2__3), .FilterDout_1__2__2 (
          CacheFilter_1__2__2), .FilterDout_1__2__1 (CacheFilter_1__2__1), .FilterDout_1__2__0 (
          CacheFilter_1__2__0), .FilterDout_1__3__7 (CacheFilter_1__3__7), .FilterDout_1__3__6 (
          CacheFilter_1__3__6), .FilterDout_1__3__5 (CacheFilter_1__3__5), .FilterDout_1__3__4 (
          CacheFilter_1__3__4), .FilterDout_1__3__3 (CacheFilter_1__3__3), .FilterDout_1__3__2 (
          CacheFilter_1__3__2), .FilterDout_1__3__1 (CacheFilter_1__3__1), .FilterDout_1__3__0 (
          CacheFilter_1__3__0), .FilterDout_1__4__7 (CacheFilter_1__4__7), .FilterDout_1__4__6 (
          CacheFilter_1__4__6), .FilterDout_1__4__5 (CacheFilter_1__4__5), .FilterDout_1__4__4 (
          CacheFilter_1__4__4), .FilterDout_1__4__3 (CacheFilter_1__4__3), .FilterDout_1__4__2 (
          CacheFilter_1__4__2), .FilterDout_1__4__1 (CacheFilter_1__4__1), .FilterDout_1__4__0 (
          CacheFilter_1__4__0), .FilterDout_2__0__7 (CacheFilter_2__0__7), .FilterDout_2__0__6 (
          CacheFilter_2__0__6), .FilterDout_2__0__5 (CacheFilter_2__0__5), .FilterDout_2__0__4 (
          CacheFilter_2__0__4), .FilterDout_2__0__3 (CacheFilter_2__0__3), .FilterDout_2__0__2 (
          CacheFilter_2__0__2), .FilterDout_2__0__1 (CacheFilter_2__0__1), .FilterDout_2__0__0 (
          CacheFilter_2__0__0), .FilterDout_2__1__7 (CacheFilter_2__1__7), .FilterDout_2__1__6 (
          CacheFilter_2__1__6), .FilterDout_2__1__5 (CacheFilter_2__1__5), .FilterDout_2__1__4 (
          CacheFilter_2__1__4), .FilterDout_2__1__3 (CacheFilter_2__1__3), .FilterDout_2__1__2 (
          CacheFilter_2__1__2), .FilterDout_2__1__1 (CacheFilter_2__1__1), .FilterDout_2__1__0 (
          CacheFilter_2__1__0), .FilterDout_2__2__7 (CacheFilter_2__2__7), .FilterDout_2__2__6 (
          CacheFilter_2__2__6), .FilterDout_2__2__5 (CacheFilter_2__2__5), .FilterDout_2__2__4 (
          CacheFilter_2__2__4), .FilterDout_2__2__3 (CacheFilter_2__2__3), .FilterDout_2__2__2 (
          CacheFilter_2__2__2), .FilterDout_2__2__1 (CacheFilter_2__2__1), .FilterDout_2__2__0 (
          CacheFilter_2__2__0), .FilterDout_2__3__7 (CacheFilter_2__3__7), .FilterDout_2__3__6 (
          CacheFilter_2__3__6), .FilterDout_2__3__5 (CacheFilter_2__3__5), .FilterDout_2__3__4 (
          CacheFilter_2__3__4), .FilterDout_2__3__3 (CacheFilter_2__3__3), .FilterDout_2__3__2 (
          CacheFilter_2__3__2), .FilterDout_2__3__1 (CacheFilter_2__3__1), .FilterDout_2__3__0 (
          CacheFilter_2__3__0), .FilterDout_2__4__7 (CacheFilter_2__4__7), .FilterDout_2__4__6 (
          CacheFilter_2__4__6), .FilterDout_2__4__5 (CacheFilter_2__4__5), .FilterDout_2__4__4 (
          CacheFilter_2__4__4), .FilterDout_2__4__3 (CacheFilter_2__4__3), .FilterDout_2__4__2 (
          CacheFilter_2__4__2), .FilterDout_2__4__1 (CacheFilter_2__4__1), .FilterDout_2__4__0 (
          CacheFilter_2__4__0), .FilterDout_3__0__7 (CacheFilter_3__0__7), .FilterDout_3__0__6 (
          CacheFilter_3__0__6), .FilterDout_3__0__5 (CacheFilter_3__0__5), .FilterDout_3__0__4 (
          CacheFilter_3__0__4), .FilterDout_3__0__3 (CacheFilter_3__0__3), .FilterDout_3__0__2 (
          CacheFilter_3__0__2), .FilterDout_3__0__1 (CacheFilter_3__0__1), .FilterDout_3__0__0 (
          CacheFilter_3__0__0), .FilterDout_3__1__7 (CacheFilter_3__1__7), .FilterDout_3__1__6 (
          CacheFilter_3__1__6), .FilterDout_3__1__5 (CacheFilter_3__1__5), .FilterDout_3__1__4 (
          CacheFilter_3__1__4), .FilterDout_3__1__3 (CacheFilter_3__1__3), .FilterDout_3__1__2 (
          CacheFilter_3__1__2), .FilterDout_3__1__1 (CacheFilter_3__1__1), .FilterDout_3__1__0 (
          CacheFilter_3__1__0), .FilterDout_3__2__7 (CacheFilter_3__2__7), .FilterDout_3__2__6 (
          CacheFilter_3__2__6), .FilterDout_3__2__5 (CacheFilter_3__2__5), .FilterDout_3__2__4 (
          CacheFilter_3__2__4), .FilterDout_3__2__3 (CacheFilter_3__2__3), .FilterDout_3__2__2 (
          CacheFilter_3__2__2), .FilterDout_3__2__1 (CacheFilter_3__2__1), .FilterDout_3__2__0 (
          CacheFilter_3__2__0), .FilterDout_3__3__7 (CacheFilter_3__3__7), .FilterDout_3__3__6 (
          CacheFilter_3__3__6), .FilterDout_3__3__5 (CacheFilter_3__3__5), .FilterDout_3__3__4 (
          CacheFilter_3__3__4), .FilterDout_3__3__3 (CacheFilter_3__3__3), .FilterDout_3__3__2 (
          CacheFilter_3__3__2), .FilterDout_3__3__1 (CacheFilter_3__3__1), .FilterDout_3__3__0 (
          CacheFilter_3__3__0), .FilterDout_3__4__7 (CacheFilter_3__4__7), .FilterDout_3__4__6 (
          CacheFilter_3__4__6), .FilterDout_3__4__5 (CacheFilter_3__4__5), .FilterDout_3__4__4 (
          CacheFilter_3__4__4), .FilterDout_3__4__3 (CacheFilter_3__4__3), .FilterDout_3__4__2 (
          CacheFilter_3__4__2), .FilterDout_3__4__1 (CacheFilter_3__4__1), .FilterDout_3__4__0 (
          CacheFilter_3__4__0), .FilterDout_4__0__7 (CacheFilter_4__0__7), .FilterDout_4__0__6 (
          CacheFilter_4__0__6), .FilterDout_4__0__5 (CacheFilter_4__0__5), .FilterDout_4__0__4 (
          CacheFilter_4__0__4), .FilterDout_4__0__3 (CacheFilter_4__0__3), .FilterDout_4__0__2 (
          CacheFilter_4__0__2), .FilterDout_4__0__1 (CacheFilter_4__0__1), .FilterDout_4__0__0 (
          CacheFilter_4__0__0), .FilterDout_4__1__7 (CacheFilter_4__1__7), .FilterDout_4__1__6 (
          CacheFilter_4__1__6), .FilterDout_4__1__5 (CacheFilter_4__1__5), .FilterDout_4__1__4 (
          CacheFilter_4__1__4), .FilterDout_4__1__3 (CacheFilter_4__1__3), .FilterDout_4__1__2 (
          CacheFilter_4__1__2), .FilterDout_4__1__1 (CacheFilter_4__1__1), .FilterDout_4__1__0 (
          CacheFilter_4__1__0), .FilterDout_4__2__7 (CacheFilter_4__2__7), .FilterDout_4__2__6 (
          CacheFilter_4__2__6), .FilterDout_4__2__5 (CacheFilter_4__2__5), .FilterDout_4__2__4 (
          CacheFilter_4__2__4), .FilterDout_4__2__3 (CacheFilter_4__2__3), .FilterDout_4__2__2 (
          CacheFilter_4__2__2), .FilterDout_4__2__1 (CacheFilter_4__2__1), .FilterDout_4__2__0 (
          CacheFilter_4__2__0), .FilterDout_4__3__7 (CacheFilter_4__3__7), .FilterDout_4__3__6 (
          CacheFilter_4__3__6), .FilterDout_4__3__5 (CacheFilter_4__3__5), .FilterDout_4__3__4 (
          CacheFilter_4__3__4), .FilterDout_4__3__3 (CacheFilter_4__3__3), .FilterDout_4__3__2 (
          CacheFilter_4__3__2), .FilterDout_4__3__1 (CacheFilter_4__3__1), .FilterDout_4__3__0 (
          CacheFilter_4__3__0), .FilterDout_4__4__7 (CacheFilter_4__4__7), .FilterDout_4__4__6 (
          CacheFilter_4__4__6), .FilterDout_4__4__5 (CacheFilter_4__4__5), .FilterDout_4__4__4 (
          CacheFilter_4__4__4), .FilterDout_4__4__3 (CacheFilter_4__4__3), .FilterDout_4__4__2 (
          CacheFilter_4__4__2), .FilterDout_4__4__1 (CacheFilter_4__4__1), .FilterDout_4__4__0 (
          CacheFilter_4__4__0), .WindowDout_0__0__7 (CacheWindow_0__0__7), .WindowDout_0__0__6 (
          CacheWindow_0__0__6), .WindowDout_0__0__5 (CacheWindow_0__0__5), .WindowDout_0__0__4 (
          CacheWindow_0__0__4), .WindowDout_0__0__3 (CacheWindow_0__0__3), .WindowDout_0__0__2 (
          CacheWindow_0__0__2), .WindowDout_0__0__1 (CacheWindow_0__0__1), .WindowDout_0__0__0 (
          CacheWindow_0__0__0), .WindowDout_0__1__7 (CacheWindow_0__1__7), .WindowDout_0__1__6 (
          CacheWindow_0__1__6), .WindowDout_0__1__5 (CacheWindow_0__1__5), .WindowDout_0__1__4 (
          CacheWindow_0__1__4), .WindowDout_0__1__3 (CacheWindow_0__1__3), .WindowDout_0__1__2 (
          CacheWindow_0__1__2), .WindowDout_0__1__1 (CacheWindow_0__1__1), .WindowDout_0__1__0 (
          CacheWindow_0__1__0), .WindowDout_0__2__7 (CacheWindow_0__2__7), .WindowDout_0__2__6 (
          CacheWindow_0__2__6), .WindowDout_0__2__5 (CacheWindow_0__2__5), .WindowDout_0__2__4 (
          CacheWindow_0__2__4), .WindowDout_0__2__3 (CacheWindow_0__2__3), .WindowDout_0__2__2 (
          CacheWindow_0__2__2), .WindowDout_0__2__1 (CacheWindow_0__2__1), .WindowDout_0__2__0 (
          CacheWindow_0__2__0), .WindowDout_0__3__7 (CacheWindow_0__3__7), .WindowDout_0__3__6 (
          CacheWindow_0__3__6), .WindowDout_0__3__5 (CacheWindow_0__3__5), .WindowDout_0__3__4 (
          CacheWindow_0__3__4), .WindowDout_0__3__3 (CacheWindow_0__3__3), .WindowDout_0__3__2 (
          CacheWindow_0__3__2), .WindowDout_0__3__1 (CacheWindow_0__3__1), .WindowDout_0__3__0 (
          CacheWindow_0__3__0), .WindowDout_0__4__7 (CacheWindow_0__4__7), .WindowDout_0__4__6 (
          CacheWindow_0__4__6), .WindowDout_0__4__5 (CacheWindow_0__4__5), .WindowDout_0__4__4 (
          CacheWindow_0__4__4), .WindowDout_0__4__3 (CacheWindow_0__4__3), .WindowDout_0__4__2 (
          CacheWindow_0__4__2), .WindowDout_0__4__1 (CacheWindow_0__4__1), .WindowDout_0__4__0 (
          CacheWindow_0__4__0), .WindowDout_1__0__7 (CacheWindow_1__0__7), .WindowDout_1__0__6 (
          CacheWindow_1__0__6), .WindowDout_1__0__5 (CacheWindow_1__0__5), .WindowDout_1__0__4 (
          CacheWindow_1__0__4), .WindowDout_1__0__3 (CacheWindow_1__0__3), .WindowDout_1__0__2 (
          CacheWindow_1__0__2), .WindowDout_1__0__1 (CacheWindow_1__0__1), .WindowDout_1__0__0 (
          CacheWindow_1__0__0), .WindowDout_1__1__7 (CacheWindow_1__1__7), .WindowDout_1__1__6 (
          CacheWindow_1__1__6), .WindowDout_1__1__5 (CacheWindow_1__1__5), .WindowDout_1__1__4 (
          CacheWindow_1__1__4), .WindowDout_1__1__3 (CacheWindow_1__1__3), .WindowDout_1__1__2 (
          CacheWindow_1__1__2), .WindowDout_1__1__1 (CacheWindow_1__1__1), .WindowDout_1__1__0 (
          CacheWindow_1__1__0), .WindowDout_1__2__7 (CacheWindow_1__2__7), .WindowDout_1__2__6 (
          CacheWindow_1__2__6), .WindowDout_1__2__5 (CacheWindow_1__2__5), .WindowDout_1__2__4 (
          CacheWindow_1__2__4), .WindowDout_1__2__3 (CacheWindow_1__2__3), .WindowDout_1__2__2 (
          CacheWindow_1__2__2), .WindowDout_1__2__1 (CacheWindow_1__2__1), .WindowDout_1__2__0 (
          CacheWindow_1__2__0), .WindowDout_1__3__7 (CacheWindow_1__3__7), .WindowDout_1__3__6 (
          CacheWindow_1__3__6), .WindowDout_1__3__5 (CacheWindow_1__3__5), .WindowDout_1__3__4 (
          CacheWindow_1__3__4), .WindowDout_1__3__3 (CacheWindow_1__3__3), .WindowDout_1__3__2 (
          CacheWindow_1__3__2), .WindowDout_1__3__1 (CacheWindow_1__3__1), .WindowDout_1__3__0 (
          CacheWindow_1__3__0), .WindowDout_1__4__7 (CacheWindow_1__4__7), .WindowDout_1__4__6 (
          CacheWindow_1__4__6), .WindowDout_1__4__5 (CacheWindow_1__4__5), .WindowDout_1__4__4 (
          CacheWindow_1__4__4), .WindowDout_1__4__3 (CacheWindow_1__4__3), .WindowDout_1__4__2 (
          CacheWindow_1__4__2), .WindowDout_1__4__1 (CacheWindow_1__4__1), .WindowDout_1__4__0 (
          CacheWindow_1__4__0), .WindowDout_2__0__7 (CacheWindow_2__0__7), .WindowDout_2__0__6 (
          CacheWindow_2__0__6), .WindowDout_2__0__5 (CacheWindow_2__0__5), .WindowDout_2__0__4 (
          CacheWindow_2__0__4), .WindowDout_2__0__3 (CacheWindow_2__0__3), .WindowDout_2__0__2 (
          CacheWindow_2__0__2), .WindowDout_2__0__1 (CacheWindow_2__0__1), .WindowDout_2__0__0 (
          CacheWindow_2__0__0), .WindowDout_2__1__7 (CacheWindow_2__1__7), .WindowDout_2__1__6 (
          CacheWindow_2__1__6), .WindowDout_2__1__5 (CacheWindow_2__1__5), .WindowDout_2__1__4 (
          CacheWindow_2__1__4), .WindowDout_2__1__3 (CacheWindow_2__1__3), .WindowDout_2__1__2 (
          CacheWindow_2__1__2), .WindowDout_2__1__1 (CacheWindow_2__1__1), .WindowDout_2__1__0 (
          CacheWindow_2__1__0), .WindowDout_2__2__7 (CacheWindow_2__2__7), .WindowDout_2__2__6 (
          CacheWindow_2__2__6), .WindowDout_2__2__5 (CacheWindow_2__2__5), .WindowDout_2__2__4 (
          CacheWindow_2__2__4), .WindowDout_2__2__3 (CacheWindow_2__2__3), .WindowDout_2__2__2 (
          CacheWindow_2__2__2), .WindowDout_2__2__1 (CacheWindow_2__2__1), .WindowDout_2__2__0 (
          CacheWindow_2__2__0), .WindowDout_2__3__7 (CacheWindow_2__3__7), .WindowDout_2__3__6 (
          CacheWindow_2__3__6), .WindowDout_2__3__5 (CacheWindow_2__3__5), .WindowDout_2__3__4 (
          CacheWindow_2__3__4), .WindowDout_2__3__3 (CacheWindow_2__3__3), .WindowDout_2__3__2 (
          CacheWindow_2__3__2), .WindowDout_2__3__1 (CacheWindow_2__3__1), .WindowDout_2__3__0 (
          CacheWindow_2__3__0), .WindowDout_2__4__7 (CacheWindow_2__4__7), .WindowDout_2__4__6 (
          CacheWindow_2__4__6), .WindowDout_2__4__5 (CacheWindow_2__4__5), .WindowDout_2__4__4 (
          CacheWindow_2__4__4), .WindowDout_2__4__3 (CacheWindow_2__4__3), .WindowDout_2__4__2 (
          CacheWindow_2__4__2), .WindowDout_2__4__1 (CacheWindow_2__4__1), .WindowDout_2__4__0 (
          CacheWindow_2__4__0), .WindowDout_3__0__7 (CacheWindow_3__0__7), .WindowDout_3__0__6 (
          CacheWindow_3__0__6), .WindowDout_3__0__5 (CacheWindow_3__0__5), .WindowDout_3__0__4 (
          CacheWindow_3__0__4), .WindowDout_3__0__3 (CacheWindow_3__0__3), .WindowDout_3__0__2 (
          CacheWindow_3__0__2), .WindowDout_3__0__1 (CacheWindow_3__0__1), .WindowDout_3__0__0 (
          CacheWindow_3__0__0), .WindowDout_3__1__7 (CacheWindow_3__1__7), .WindowDout_3__1__6 (
          CacheWindow_3__1__6), .WindowDout_3__1__5 (CacheWindow_3__1__5), .WindowDout_3__1__4 (
          CacheWindow_3__1__4), .WindowDout_3__1__3 (CacheWindow_3__1__3), .WindowDout_3__1__2 (
          CacheWindow_3__1__2), .WindowDout_3__1__1 (CacheWindow_3__1__1), .WindowDout_3__1__0 (
          CacheWindow_3__1__0), .WindowDout_3__2__7 (CacheWindow_3__2__7), .WindowDout_3__2__6 (
          CacheWindow_3__2__6), .WindowDout_3__2__5 (CacheWindow_3__2__5), .WindowDout_3__2__4 (
          CacheWindow_3__2__4), .WindowDout_3__2__3 (CacheWindow_3__2__3), .WindowDout_3__2__2 (
          CacheWindow_3__2__2), .WindowDout_3__2__1 (CacheWindow_3__2__1), .WindowDout_3__2__0 (
          CacheWindow_3__2__0), .WindowDout_3__3__7 (CacheWindow_3__3__7), .WindowDout_3__3__6 (
          CacheWindow_3__3__6), .WindowDout_3__3__5 (CacheWindow_3__3__5), .WindowDout_3__3__4 (
          CacheWindow_3__3__4), .WindowDout_3__3__3 (CacheWindow_3__3__3), .WindowDout_3__3__2 (
          CacheWindow_3__3__2), .WindowDout_3__3__1 (CacheWindow_3__3__1), .WindowDout_3__3__0 (
          CacheWindow_3__3__0), .WindowDout_3__4__7 (CacheWindow_3__4__7), .WindowDout_3__4__6 (
          CacheWindow_3__4__6), .WindowDout_3__4__5 (CacheWindow_3__4__5), .WindowDout_3__4__4 (
          CacheWindow_3__4__4), .WindowDout_3__4__3 (CacheWindow_3__4__3), .WindowDout_3__4__2 (
          CacheWindow_3__4__2), .WindowDout_3__4__1 (CacheWindow_3__4__1), .WindowDout_3__4__0 (
          CacheWindow_3__4__0), .WindowDout_4__0__7 (CacheWindow_4__0__7), .WindowDout_4__0__6 (
          CacheWindow_4__0__6), .WindowDout_4__0__5 (CacheWindow_4__0__5), .WindowDout_4__0__4 (
          CacheWindow_4__0__4), .WindowDout_4__0__3 (CacheWindow_4__0__3), .WindowDout_4__0__2 (
          CacheWindow_4__0__2), .WindowDout_4__0__1 (CacheWindow_4__0__1), .WindowDout_4__0__0 (
          CacheWindow_4__0__0), .WindowDout_4__1__7 (CacheWindow_4__1__7), .WindowDout_4__1__6 (
          CacheWindow_4__1__6), .WindowDout_4__1__5 (CacheWindow_4__1__5), .WindowDout_4__1__4 (
          CacheWindow_4__1__4), .WindowDout_4__1__3 (CacheWindow_4__1__3), .WindowDout_4__1__2 (
          CacheWindow_4__1__2), .WindowDout_4__1__1 (CacheWindow_4__1__1), .WindowDout_4__1__0 (
          CacheWindow_4__1__0), .WindowDout_4__2__7 (CacheWindow_4__2__7), .WindowDout_4__2__6 (
          CacheWindow_4__2__6), .WindowDout_4__2__5 (CacheWindow_4__2__5), .WindowDout_4__2__4 (
          CacheWindow_4__2__4), .WindowDout_4__2__3 (CacheWindow_4__2__3), .WindowDout_4__2__2 (
          CacheWindow_4__2__2), .WindowDout_4__2__1 (CacheWindow_4__2__1), .WindowDout_4__2__0 (
          CacheWindow_4__2__0), .WindowDout_4__3__7 (CacheWindow_4__3__7), .WindowDout_4__3__6 (
          CacheWindow_4__3__6), .WindowDout_4__3__5 (CacheWindow_4__3__5), .WindowDout_4__3__4 (
          CacheWindow_4__3__4), .WindowDout_4__3__3 (CacheWindow_4__3__3), .WindowDout_4__3__2 (
          CacheWindow_4__3__2), .WindowDout_4__3__1 (CacheWindow_4__3__1), .WindowDout_4__3__0 (
          CacheWindow_4__3__0), .WindowDout_4__4__7 (CacheWindow_4__4__7), .WindowDout_4__4__6 (
          CacheWindow_4__4__6), .WindowDout_4__4__5 (CacheWindow_4__4__5), .WindowDout_4__4__4 (
          CacheWindow_4__4__4), .WindowDout_4__4__3 (CacheWindow_4__4__3), .WindowDout_4__4__2 (
          CacheWindow_4__4__2), .WindowDout_4__4__1 (CacheWindow_4__4__1), .WindowDout_4__4__0 (
          CacheWindow_4__4__0), .ResultWR (GND0), .ResultDin ({AccResult_7,
          AccResult_6,AccResult_5,AccResult_4,AccResult_3,AccResult_2,
          AccResult_1,AccResult_0}), .ResultDout ({MemDin_7,MemDin_6,MemDin_5,
          MemDin_4,MemDin_3,MemDin_2,MemDin_1,MemDin_0})) ;
    assign GND0 = 0 ;
endmodule


module cache ( CLK, RST, FilterSize, FilterWR, WindowWR, Din, FilterDout_0__0__7, 
               FilterDout_0__0__6, FilterDout_0__0__5, FilterDout_0__0__4, 
               FilterDout_0__0__3, FilterDout_0__0__2, FilterDout_0__0__1, 
               FilterDout_0__0__0, FilterDout_0__1__7, FilterDout_0__1__6, 
               FilterDout_0__1__5, FilterDout_0__1__4, FilterDout_0__1__3, 
               FilterDout_0__1__2, FilterDout_0__1__1, FilterDout_0__1__0, 
               FilterDout_0__2__7, FilterDout_0__2__6, FilterDout_0__2__5, 
               FilterDout_0__2__4, FilterDout_0__2__3, FilterDout_0__2__2, 
               FilterDout_0__2__1, FilterDout_0__2__0, FilterDout_0__3__7, 
               FilterDout_0__3__6, FilterDout_0__3__5, FilterDout_0__3__4, 
               FilterDout_0__3__3, FilterDout_0__3__2, FilterDout_0__3__1, 
               FilterDout_0__3__0, FilterDout_0__4__7, FilterDout_0__4__6, 
               FilterDout_0__4__5, FilterDout_0__4__4, FilterDout_0__4__3, 
               FilterDout_0__4__2, FilterDout_0__4__1, FilterDout_0__4__0, 
               FilterDout_1__0__7, FilterDout_1__0__6, FilterDout_1__0__5, 
               FilterDout_1__0__4, FilterDout_1__0__3, FilterDout_1__0__2, 
               FilterDout_1__0__1, FilterDout_1__0__0, FilterDout_1__1__7, 
               FilterDout_1__1__6, FilterDout_1__1__5, FilterDout_1__1__4, 
               FilterDout_1__1__3, FilterDout_1__1__2, FilterDout_1__1__1, 
               FilterDout_1__1__0, FilterDout_1__2__7, FilterDout_1__2__6, 
               FilterDout_1__2__5, FilterDout_1__2__4, FilterDout_1__2__3, 
               FilterDout_1__2__2, FilterDout_1__2__1, FilterDout_1__2__0, 
               FilterDout_1__3__7, FilterDout_1__3__6, FilterDout_1__3__5, 
               FilterDout_1__3__4, FilterDout_1__3__3, FilterDout_1__3__2, 
               FilterDout_1__3__1, FilterDout_1__3__0, FilterDout_1__4__7, 
               FilterDout_1__4__6, FilterDout_1__4__5, FilterDout_1__4__4, 
               FilterDout_1__4__3, FilterDout_1__4__2, FilterDout_1__4__1, 
               FilterDout_1__4__0, FilterDout_2__0__7, FilterDout_2__0__6, 
               FilterDout_2__0__5, FilterDout_2__0__4, FilterDout_2__0__3, 
               FilterDout_2__0__2, FilterDout_2__0__1, FilterDout_2__0__0, 
               FilterDout_2__1__7, FilterDout_2__1__6, FilterDout_2__1__5, 
               FilterDout_2__1__4, FilterDout_2__1__3, FilterDout_2__1__2, 
               FilterDout_2__1__1, FilterDout_2__1__0, FilterDout_2__2__7, 
               FilterDout_2__2__6, FilterDout_2__2__5, FilterDout_2__2__4, 
               FilterDout_2__2__3, FilterDout_2__2__2, FilterDout_2__2__1, 
               FilterDout_2__2__0, FilterDout_2__3__7, FilterDout_2__3__6, 
               FilterDout_2__3__5, FilterDout_2__3__4, FilterDout_2__3__3, 
               FilterDout_2__3__2, FilterDout_2__3__1, FilterDout_2__3__0, 
               FilterDout_2__4__7, FilterDout_2__4__6, FilterDout_2__4__5, 
               FilterDout_2__4__4, FilterDout_2__4__3, FilterDout_2__4__2, 
               FilterDout_2__4__1, FilterDout_2__4__0, FilterDout_3__0__7, 
               FilterDout_3__0__6, FilterDout_3__0__5, FilterDout_3__0__4, 
               FilterDout_3__0__3, FilterDout_3__0__2, FilterDout_3__0__1, 
               FilterDout_3__0__0, FilterDout_3__1__7, FilterDout_3__1__6, 
               FilterDout_3__1__5, FilterDout_3__1__4, FilterDout_3__1__3, 
               FilterDout_3__1__2, FilterDout_3__1__1, FilterDout_3__1__0, 
               FilterDout_3__2__7, FilterDout_3__2__6, FilterDout_3__2__5, 
               FilterDout_3__2__4, FilterDout_3__2__3, FilterDout_3__2__2, 
               FilterDout_3__2__1, FilterDout_3__2__0, FilterDout_3__3__7, 
               FilterDout_3__3__6, FilterDout_3__3__5, FilterDout_3__3__4, 
               FilterDout_3__3__3, FilterDout_3__3__2, FilterDout_3__3__1, 
               FilterDout_3__3__0, FilterDout_3__4__7, FilterDout_3__4__6, 
               FilterDout_3__4__5, FilterDout_3__4__4, FilterDout_3__4__3, 
               FilterDout_3__4__2, FilterDout_3__4__1, FilterDout_3__4__0, 
               FilterDout_4__0__7, FilterDout_4__0__6, FilterDout_4__0__5, 
               FilterDout_4__0__4, FilterDout_4__0__3, FilterDout_4__0__2, 
               FilterDout_4__0__1, FilterDout_4__0__0, FilterDout_4__1__7, 
               FilterDout_4__1__6, FilterDout_4__1__5, FilterDout_4__1__4, 
               FilterDout_4__1__3, FilterDout_4__1__2, FilterDout_4__1__1, 
               FilterDout_4__1__0, FilterDout_4__2__7, FilterDout_4__2__6, 
               FilterDout_4__2__5, FilterDout_4__2__4, FilterDout_4__2__3, 
               FilterDout_4__2__2, FilterDout_4__2__1, FilterDout_4__2__0, 
               FilterDout_4__3__7, FilterDout_4__3__6, FilterDout_4__3__5, 
               FilterDout_4__3__4, FilterDout_4__3__3, FilterDout_4__3__2, 
               FilterDout_4__3__1, FilterDout_4__3__0, FilterDout_4__4__7, 
               FilterDout_4__4__6, FilterDout_4__4__5, FilterDout_4__4__4, 
               FilterDout_4__4__3, FilterDout_4__4__2, FilterDout_4__4__1, 
               FilterDout_4__4__0, WindowDout_0__0__7, WindowDout_0__0__6, 
               WindowDout_0__0__5, WindowDout_0__0__4, WindowDout_0__0__3, 
               WindowDout_0__0__2, WindowDout_0__0__1, WindowDout_0__0__0, 
               WindowDout_0__1__7, WindowDout_0__1__6, WindowDout_0__1__5, 
               WindowDout_0__1__4, WindowDout_0__1__3, WindowDout_0__1__2, 
               WindowDout_0__1__1, WindowDout_0__1__0, WindowDout_0__2__7, 
               WindowDout_0__2__6, WindowDout_0__2__5, WindowDout_0__2__4, 
               WindowDout_0__2__3, WindowDout_0__2__2, WindowDout_0__2__1, 
               WindowDout_0__2__0, WindowDout_0__3__7, WindowDout_0__3__6, 
               WindowDout_0__3__5, WindowDout_0__3__4, WindowDout_0__3__3, 
               WindowDout_0__3__2, WindowDout_0__3__1, WindowDout_0__3__0, 
               WindowDout_0__4__7, WindowDout_0__4__6, WindowDout_0__4__5, 
               WindowDout_0__4__4, WindowDout_0__4__3, WindowDout_0__4__2, 
               WindowDout_0__4__1, WindowDout_0__4__0, WindowDout_1__0__7, 
               WindowDout_1__0__6, WindowDout_1__0__5, WindowDout_1__0__4, 
               WindowDout_1__0__3, WindowDout_1__0__2, WindowDout_1__0__1, 
               WindowDout_1__0__0, WindowDout_1__1__7, WindowDout_1__1__6, 
               WindowDout_1__1__5, WindowDout_1__1__4, WindowDout_1__1__3, 
               WindowDout_1__1__2, WindowDout_1__1__1, WindowDout_1__1__0, 
               WindowDout_1__2__7, WindowDout_1__2__6, WindowDout_1__2__5, 
               WindowDout_1__2__4, WindowDout_1__2__3, WindowDout_1__2__2, 
               WindowDout_1__2__1, WindowDout_1__2__0, WindowDout_1__3__7, 
               WindowDout_1__3__6, WindowDout_1__3__5, WindowDout_1__3__4, 
               WindowDout_1__3__3, WindowDout_1__3__2, WindowDout_1__3__1, 
               WindowDout_1__3__0, WindowDout_1__4__7, WindowDout_1__4__6, 
               WindowDout_1__4__5, WindowDout_1__4__4, WindowDout_1__4__3, 
               WindowDout_1__4__2, WindowDout_1__4__1, WindowDout_1__4__0, 
               WindowDout_2__0__7, WindowDout_2__0__6, WindowDout_2__0__5, 
               WindowDout_2__0__4, WindowDout_2__0__3, WindowDout_2__0__2, 
               WindowDout_2__0__1, WindowDout_2__0__0, WindowDout_2__1__7, 
               WindowDout_2__1__6, WindowDout_2__1__5, WindowDout_2__1__4, 
               WindowDout_2__1__3, WindowDout_2__1__2, WindowDout_2__1__1, 
               WindowDout_2__1__0, WindowDout_2__2__7, WindowDout_2__2__6, 
               WindowDout_2__2__5, WindowDout_2__2__4, WindowDout_2__2__3, 
               WindowDout_2__2__2, WindowDout_2__2__1, WindowDout_2__2__0, 
               WindowDout_2__3__7, WindowDout_2__3__6, WindowDout_2__3__5, 
               WindowDout_2__3__4, WindowDout_2__3__3, WindowDout_2__3__2, 
               WindowDout_2__3__1, WindowDout_2__3__0, WindowDout_2__4__7, 
               WindowDout_2__4__6, WindowDout_2__4__5, WindowDout_2__4__4, 
               WindowDout_2__4__3, WindowDout_2__4__2, WindowDout_2__4__1, 
               WindowDout_2__4__0, WindowDout_3__0__7, WindowDout_3__0__6, 
               WindowDout_3__0__5, WindowDout_3__0__4, WindowDout_3__0__3, 
               WindowDout_3__0__2, WindowDout_3__0__1, WindowDout_3__0__0, 
               WindowDout_3__1__7, WindowDout_3__1__6, WindowDout_3__1__5, 
               WindowDout_3__1__4, WindowDout_3__1__3, WindowDout_3__1__2, 
               WindowDout_3__1__1, WindowDout_3__1__0, WindowDout_3__2__7, 
               WindowDout_3__2__6, WindowDout_3__2__5, WindowDout_3__2__4, 
               WindowDout_3__2__3, WindowDout_3__2__2, WindowDout_3__2__1, 
               WindowDout_3__2__0, WindowDout_3__3__7, WindowDout_3__3__6, 
               WindowDout_3__3__5, WindowDout_3__3__4, WindowDout_3__3__3, 
               WindowDout_3__3__2, WindowDout_3__3__1, WindowDout_3__3__0, 
               WindowDout_3__4__7, WindowDout_3__4__6, WindowDout_3__4__5, 
               WindowDout_3__4__4, WindowDout_3__4__3, WindowDout_3__4__2, 
               WindowDout_3__4__1, WindowDout_3__4__0, WindowDout_4__0__7, 
               WindowDout_4__0__6, WindowDout_4__0__5, WindowDout_4__0__4, 
               WindowDout_4__0__3, WindowDout_4__0__2, WindowDout_4__0__1, 
               WindowDout_4__0__0, WindowDout_4__1__7, WindowDout_4__1__6, 
               WindowDout_4__1__5, WindowDout_4__1__4, WindowDout_4__1__3, 
               WindowDout_4__1__2, WindowDout_4__1__1, WindowDout_4__1__0, 
               WindowDout_4__2__7, WindowDout_4__2__6, WindowDout_4__2__5, 
               WindowDout_4__2__4, WindowDout_4__2__3, WindowDout_4__2__2, 
               WindowDout_4__2__1, WindowDout_4__2__0, WindowDout_4__3__7, 
               WindowDout_4__3__6, WindowDout_4__3__5, WindowDout_4__3__4, 
               WindowDout_4__3__3, WindowDout_4__3__2, WindowDout_4__3__1, 
               WindowDout_4__3__0, WindowDout_4__4__7, WindowDout_4__4__6, 
               WindowDout_4__4__5, WindowDout_4__4__4, WindowDout_4__4__3, 
               WindowDout_4__4__2, WindowDout_4__4__1, WindowDout_4__4__0, 
               ResultWR, ResultDin, ResultDout ) ;

    input CLK ;
    input RST ;
    input FilterSize ;
    input FilterWR ;
    input WindowWR ;
    input [39:0]Din ;
    output FilterDout_0__0__7 ;
    output FilterDout_0__0__6 ;
    output FilterDout_0__0__5 ;
    output FilterDout_0__0__4 ;
    output FilterDout_0__0__3 ;
    output FilterDout_0__0__2 ;
    output FilterDout_0__0__1 ;
    output FilterDout_0__0__0 ;
    output FilterDout_0__1__7 ;
    output FilterDout_0__1__6 ;
    output FilterDout_0__1__5 ;
    output FilterDout_0__1__4 ;
    output FilterDout_0__1__3 ;
    output FilterDout_0__1__2 ;
    output FilterDout_0__1__1 ;
    output FilterDout_0__1__0 ;
    output FilterDout_0__2__7 ;
    output FilterDout_0__2__6 ;
    output FilterDout_0__2__5 ;
    output FilterDout_0__2__4 ;
    output FilterDout_0__2__3 ;
    output FilterDout_0__2__2 ;
    output FilterDout_0__2__1 ;
    output FilterDout_0__2__0 ;
    output FilterDout_0__3__7 ;
    output FilterDout_0__3__6 ;
    output FilterDout_0__3__5 ;
    output FilterDout_0__3__4 ;
    output FilterDout_0__3__3 ;
    output FilterDout_0__3__2 ;
    output FilterDout_0__3__1 ;
    output FilterDout_0__3__0 ;
    output FilterDout_0__4__7 ;
    output FilterDout_0__4__6 ;
    output FilterDout_0__4__5 ;
    output FilterDout_0__4__4 ;
    output FilterDout_0__4__3 ;
    output FilterDout_0__4__2 ;
    output FilterDout_0__4__1 ;
    output FilterDout_0__4__0 ;
    output FilterDout_1__0__7 ;
    output FilterDout_1__0__6 ;
    output FilterDout_1__0__5 ;
    output FilterDout_1__0__4 ;
    output FilterDout_1__0__3 ;
    output FilterDout_1__0__2 ;
    output FilterDout_1__0__1 ;
    output FilterDout_1__0__0 ;
    output FilterDout_1__1__7 ;
    output FilterDout_1__1__6 ;
    output FilterDout_1__1__5 ;
    output FilterDout_1__1__4 ;
    output FilterDout_1__1__3 ;
    output FilterDout_1__1__2 ;
    output FilterDout_1__1__1 ;
    output FilterDout_1__1__0 ;
    output FilterDout_1__2__7 ;
    output FilterDout_1__2__6 ;
    output FilterDout_1__2__5 ;
    output FilterDout_1__2__4 ;
    output FilterDout_1__2__3 ;
    output FilterDout_1__2__2 ;
    output FilterDout_1__2__1 ;
    output FilterDout_1__2__0 ;
    output FilterDout_1__3__7 ;
    output FilterDout_1__3__6 ;
    output FilterDout_1__3__5 ;
    output FilterDout_1__3__4 ;
    output FilterDout_1__3__3 ;
    output FilterDout_1__3__2 ;
    output FilterDout_1__3__1 ;
    output FilterDout_1__3__0 ;
    output FilterDout_1__4__7 ;
    output FilterDout_1__4__6 ;
    output FilterDout_1__4__5 ;
    output FilterDout_1__4__4 ;
    output FilterDout_1__4__3 ;
    output FilterDout_1__4__2 ;
    output FilterDout_1__4__1 ;
    output FilterDout_1__4__0 ;
    output FilterDout_2__0__7 ;
    output FilterDout_2__0__6 ;
    output FilterDout_2__0__5 ;
    output FilterDout_2__0__4 ;
    output FilterDout_2__0__3 ;
    output FilterDout_2__0__2 ;
    output FilterDout_2__0__1 ;
    output FilterDout_2__0__0 ;
    output FilterDout_2__1__7 ;
    output FilterDout_2__1__6 ;
    output FilterDout_2__1__5 ;
    output FilterDout_2__1__4 ;
    output FilterDout_2__1__3 ;
    output FilterDout_2__1__2 ;
    output FilterDout_2__1__1 ;
    output FilterDout_2__1__0 ;
    output FilterDout_2__2__7 ;
    output FilterDout_2__2__6 ;
    output FilterDout_2__2__5 ;
    output FilterDout_2__2__4 ;
    output FilterDout_2__2__3 ;
    output FilterDout_2__2__2 ;
    output FilterDout_2__2__1 ;
    output FilterDout_2__2__0 ;
    output FilterDout_2__3__7 ;
    output FilterDout_2__3__6 ;
    output FilterDout_2__3__5 ;
    output FilterDout_2__3__4 ;
    output FilterDout_2__3__3 ;
    output FilterDout_2__3__2 ;
    output FilterDout_2__3__1 ;
    output FilterDout_2__3__0 ;
    output FilterDout_2__4__7 ;
    output FilterDout_2__4__6 ;
    output FilterDout_2__4__5 ;
    output FilterDout_2__4__4 ;
    output FilterDout_2__4__3 ;
    output FilterDout_2__4__2 ;
    output FilterDout_2__4__1 ;
    output FilterDout_2__4__0 ;
    output FilterDout_3__0__7 ;
    output FilterDout_3__0__6 ;
    output FilterDout_3__0__5 ;
    output FilterDout_3__0__4 ;
    output FilterDout_3__0__3 ;
    output FilterDout_3__0__2 ;
    output FilterDout_3__0__1 ;
    output FilterDout_3__0__0 ;
    output FilterDout_3__1__7 ;
    output FilterDout_3__1__6 ;
    output FilterDout_3__1__5 ;
    output FilterDout_3__1__4 ;
    output FilterDout_3__1__3 ;
    output FilterDout_3__1__2 ;
    output FilterDout_3__1__1 ;
    output FilterDout_3__1__0 ;
    output FilterDout_3__2__7 ;
    output FilterDout_3__2__6 ;
    output FilterDout_3__2__5 ;
    output FilterDout_3__2__4 ;
    output FilterDout_3__2__3 ;
    output FilterDout_3__2__2 ;
    output FilterDout_3__2__1 ;
    output FilterDout_3__2__0 ;
    output FilterDout_3__3__7 ;
    output FilterDout_3__3__6 ;
    output FilterDout_3__3__5 ;
    output FilterDout_3__3__4 ;
    output FilterDout_3__3__3 ;
    output FilterDout_3__3__2 ;
    output FilterDout_3__3__1 ;
    output FilterDout_3__3__0 ;
    output FilterDout_3__4__7 ;
    output FilterDout_3__4__6 ;
    output FilterDout_3__4__5 ;
    output FilterDout_3__4__4 ;
    output FilterDout_3__4__3 ;
    output FilterDout_3__4__2 ;
    output FilterDout_3__4__1 ;
    output FilterDout_3__4__0 ;
    output FilterDout_4__0__7 ;
    output FilterDout_4__0__6 ;
    output FilterDout_4__0__5 ;
    output FilterDout_4__0__4 ;
    output FilterDout_4__0__3 ;
    output FilterDout_4__0__2 ;
    output FilterDout_4__0__1 ;
    output FilterDout_4__0__0 ;
    output FilterDout_4__1__7 ;
    output FilterDout_4__1__6 ;
    output FilterDout_4__1__5 ;
    output FilterDout_4__1__4 ;
    output FilterDout_4__1__3 ;
    output FilterDout_4__1__2 ;
    output FilterDout_4__1__1 ;
    output FilterDout_4__1__0 ;
    output FilterDout_4__2__7 ;
    output FilterDout_4__2__6 ;
    output FilterDout_4__2__5 ;
    output FilterDout_4__2__4 ;
    output FilterDout_4__2__3 ;
    output FilterDout_4__2__2 ;
    output FilterDout_4__2__1 ;
    output FilterDout_4__2__0 ;
    output FilterDout_4__3__7 ;
    output FilterDout_4__3__6 ;
    output FilterDout_4__3__5 ;
    output FilterDout_4__3__4 ;
    output FilterDout_4__3__3 ;
    output FilterDout_4__3__2 ;
    output FilterDout_4__3__1 ;
    output FilterDout_4__3__0 ;
    output FilterDout_4__4__7 ;
    output FilterDout_4__4__6 ;
    output FilterDout_4__4__5 ;
    output FilterDout_4__4__4 ;
    output FilterDout_4__4__3 ;
    output FilterDout_4__4__2 ;
    output FilterDout_4__4__1 ;
    output FilterDout_4__4__0 ;
    output WindowDout_0__0__7 ;
    output WindowDout_0__0__6 ;
    output WindowDout_0__0__5 ;
    output WindowDout_0__0__4 ;
    output WindowDout_0__0__3 ;
    output WindowDout_0__0__2 ;
    output WindowDout_0__0__1 ;
    output WindowDout_0__0__0 ;
    output WindowDout_0__1__7 ;
    output WindowDout_0__1__6 ;
    output WindowDout_0__1__5 ;
    output WindowDout_0__1__4 ;
    output WindowDout_0__1__3 ;
    output WindowDout_0__1__2 ;
    output WindowDout_0__1__1 ;
    output WindowDout_0__1__0 ;
    output WindowDout_0__2__7 ;
    output WindowDout_0__2__6 ;
    output WindowDout_0__2__5 ;
    output WindowDout_0__2__4 ;
    output WindowDout_0__2__3 ;
    output WindowDout_0__2__2 ;
    output WindowDout_0__2__1 ;
    output WindowDout_0__2__0 ;
    output WindowDout_0__3__7 ;
    output WindowDout_0__3__6 ;
    output WindowDout_0__3__5 ;
    output WindowDout_0__3__4 ;
    output WindowDout_0__3__3 ;
    output WindowDout_0__3__2 ;
    output WindowDout_0__3__1 ;
    output WindowDout_0__3__0 ;
    output WindowDout_0__4__7 ;
    output WindowDout_0__4__6 ;
    output WindowDout_0__4__5 ;
    output WindowDout_0__4__4 ;
    output WindowDout_0__4__3 ;
    output WindowDout_0__4__2 ;
    output WindowDout_0__4__1 ;
    output WindowDout_0__4__0 ;
    output WindowDout_1__0__7 ;
    output WindowDout_1__0__6 ;
    output WindowDout_1__0__5 ;
    output WindowDout_1__0__4 ;
    output WindowDout_1__0__3 ;
    output WindowDout_1__0__2 ;
    output WindowDout_1__0__1 ;
    output WindowDout_1__0__0 ;
    output WindowDout_1__1__7 ;
    output WindowDout_1__1__6 ;
    output WindowDout_1__1__5 ;
    output WindowDout_1__1__4 ;
    output WindowDout_1__1__3 ;
    output WindowDout_1__1__2 ;
    output WindowDout_1__1__1 ;
    output WindowDout_1__1__0 ;
    output WindowDout_1__2__7 ;
    output WindowDout_1__2__6 ;
    output WindowDout_1__2__5 ;
    output WindowDout_1__2__4 ;
    output WindowDout_1__2__3 ;
    output WindowDout_1__2__2 ;
    output WindowDout_1__2__1 ;
    output WindowDout_1__2__0 ;
    output WindowDout_1__3__7 ;
    output WindowDout_1__3__6 ;
    output WindowDout_1__3__5 ;
    output WindowDout_1__3__4 ;
    output WindowDout_1__3__3 ;
    output WindowDout_1__3__2 ;
    output WindowDout_1__3__1 ;
    output WindowDout_1__3__0 ;
    output WindowDout_1__4__7 ;
    output WindowDout_1__4__6 ;
    output WindowDout_1__4__5 ;
    output WindowDout_1__4__4 ;
    output WindowDout_1__4__3 ;
    output WindowDout_1__4__2 ;
    output WindowDout_1__4__1 ;
    output WindowDout_1__4__0 ;
    output WindowDout_2__0__7 ;
    output WindowDout_2__0__6 ;
    output WindowDout_2__0__5 ;
    output WindowDout_2__0__4 ;
    output WindowDout_2__0__3 ;
    output WindowDout_2__0__2 ;
    output WindowDout_2__0__1 ;
    output WindowDout_2__0__0 ;
    output WindowDout_2__1__7 ;
    output WindowDout_2__1__6 ;
    output WindowDout_2__1__5 ;
    output WindowDout_2__1__4 ;
    output WindowDout_2__1__3 ;
    output WindowDout_2__1__2 ;
    output WindowDout_2__1__1 ;
    output WindowDout_2__1__0 ;
    output WindowDout_2__2__7 ;
    output WindowDout_2__2__6 ;
    output WindowDout_2__2__5 ;
    output WindowDout_2__2__4 ;
    output WindowDout_2__2__3 ;
    output WindowDout_2__2__2 ;
    output WindowDout_2__2__1 ;
    output WindowDout_2__2__0 ;
    output WindowDout_2__3__7 ;
    output WindowDout_2__3__6 ;
    output WindowDout_2__3__5 ;
    output WindowDout_2__3__4 ;
    output WindowDout_2__3__3 ;
    output WindowDout_2__3__2 ;
    output WindowDout_2__3__1 ;
    output WindowDout_2__3__0 ;
    output WindowDout_2__4__7 ;
    output WindowDout_2__4__6 ;
    output WindowDout_2__4__5 ;
    output WindowDout_2__4__4 ;
    output WindowDout_2__4__3 ;
    output WindowDout_2__4__2 ;
    output WindowDout_2__4__1 ;
    output WindowDout_2__4__0 ;
    output WindowDout_3__0__7 ;
    output WindowDout_3__0__6 ;
    output WindowDout_3__0__5 ;
    output WindowDout_3__0__4 ;
    output WindowDout_3__0__3 ;
    output WindowDout_3__0__2 ;
    output WindowDout_3__0__1 ;
    output WindowDout_3__0__0 ;
    output WindowDout_3__1__7 ;
    output WindowDout_3__1__6 ;
    output WindowDout_3__1__5 ;
    output WindowDout_3__1__4 ;
    output WindowDout_3__1__3 ;
    output WindowDout_3__1__2 ;
    output WindowDout_3__1__1 ;
    output WindowDout_3__1__0 ;
    output WindowDout_3__2__7 ;
    output WindowDout_3__2__6 ;
    output WindowDout_3__2__5 ;
    output WindowDout_3__2__4 ;
    output WindowDout_3__2__3 ;
    output WindowDout_3__2__2 ;
    output WindowDout_3__2__1 ;
    output WindowDout_3__2__0 ;
    output WindowDout_3__3__7 ;
    output WindowDout_3__3__6 ;
    output WindowDout_3__3__5 ;
    output WindowDout_3__3__4 ;
    output WindowDout_3__3__3 ;
    output WindowDout_3__3__2 ;
    output WindowDout_3__3__1 ;
    output WindowDout_3__3__0 ;
    output WindowDout_3__4__7 ;
    output WindowDout_3__4__6 ;
    output WindowDout_3__4__5 ;
    output WindowDout_3__4__4 ;
    output WindowDout_3__4__3 ;
    output WindowDout_3__4__2 ;
    output WindowDout_3__4__1 ;
    output WindowDout_3__4__0 ;
    output WindowDout_4__0__7 ;
    output WindowDout_4__0__6 ;
    output WindowDout_4__0__5 ;
    output WindowDout_4__0__4 ;
    output WindowDout_4__0__3 ;
    output WindowDout_4__0__2 ;
    output WindowDout_4__0__1 ;
    output WindowDout_4__0__0 ;
    output WindowDout_4__1__7 ;
    output WindowDout_4__1__6 ;
    output WindowDout_4__1__5 ;
    output WindowDout_4__1__4 ;
    output WindowDout_4__1__3 ;
    output WindowDout_4__1__2 ;
    output WindowDout_4__1__1 ;
    output WindowDout_4__1__0 ;
    output WindowDout_4__2__7 ;
    output WindowDout_4__2__6 ;
    output WindowDout_4__2__5 ;
    output WindowDout_4__2__4 ;
    output WindowDout_4__2__3 ;
    output WindowDout_4__2__2 ;
    output WindowDout_4__2__1 ;
    output WindowDout_4__2__0 ;
    output WindowDout_4__3__7 ;
    output WindowDout_4__3__6 ;
    output WindowDout_4__3__5 ;
    output WindowDout_4__3__4 ;
    output WindowDout_4__3__3 ;
    output WindowDout_4__3__2 ;
    output WindowDout_4__3__1 ;
    output WindowDout_4__3__0 ;
    output WindowDout_4__4__7 ;
    output WindowDout_4__4__6 ;
    output WindowDout_4__4__5 ;
    output WindowDout_4__4__4 ;
    output WindowDout_4__4__3 ;
    output WindowDout_4__4__2 ;
    output WindowDout_4__4__1 ;
    output WindowDout_4__4__0 ;
    input ResultWR ;
    input [7:0]ResultDin ;
    output [7:0]ResultDout ;

    wire nx82, nx86, nx96, nx106, nx116, nx126, nx136, nx146, nx156, nx166, 
         nx218, nx228, nx238, nx248, nx258, nx268, nx278, nx288, nx1897, nx1907, 
         nx1917, nx1927, nx1937, nx1947, nx1957, nx1967, nx1981, nx1991, nx2001, 
         nx2011, nx2021, nx2031, nx2041, nx2051, nx2061, nx2071, nx2081, nx2091, 
         nx2101, nx2111, nx2121, nx2131, nx2141, nx2151, nx2161, nx2171, nx2181, 
         nx2191, nx2201, nx2211, nx2221, nx2231, nx2241, nx2251, nx2261, nx2271, 
         nx2281, nx2291, nx2301, nx2311, nx2321, nx2331, nx2341, nx2351, nx2361, 
         nx2371, nx2381, nx2391, nx2401, nx2411, nx2421, nx2431, nx2441, nx2451, 
         nx2461, nx2471, nx2481, nx2491, nx2501, nx2511, nx2521, nx2531, nx2541, 
         nx2551, nx2561, nx2571, nx2581, nx2591, nx2601, nx2611, nx2621, nx2631, 
         nx2641, nx2651, nx2661, nx2671, nx2681, nx2691, nx2701, nx2711, nx2721, 
         nx2731, nx2741, nx2751, nx2761, nx2771, nx2781, nx2791, nx2801, nx2811, 
         nx2821, nx2831, nx2841, nx2851, nx2861, nx2871, nx2881, nx2891, nx2901, 
         nx2911, nx2921, nx2931, nx2941, nx2951, nx2961, nx2971, nx2981, nx2991, 
         nx3001, nx3011, nx3021, nx3031, nx3041, nx3051, nx3061, nx3071, nx3081, 
         nx3091, nx3101, nx3111, nx3121, nx3131, nx3141, nx3151, nx3161, nx3171, 
         nx3181, nx3191, nx3201, nx3211, nx3221, nx3231, nx3241, nx3251, nx3261, 
         nx3271, nx3281, nx3291, nx3301, nx3311, nx3321, nx3331, nx3341, nx3351, 
         nx3361, nx3371, nx3381, nx3391, nx3401, nx3411, nx3421, nx3431, nx3441, 
         nx3451, nx3461, nx3471, nx3481, nx3491, nx3501, nx3511, nx3521, nx3531, 
         nx3541, nx3551, nx3561, nx3571, nx3581, nx3591, nx3601, nx3611, nx3621, 
         nx3631, nx3641, nx3651, nx3661, nx3671, nx3681, nx3691, nx3701, nx3711, 
         nx3721, nx3731, nx3741, nx3751, nx3761, nx3771, nx3781, nx3791, nx3801, 
         nx3811, nx3821, nx3831, nx3841, nx3851, nx3861, nx3871, nx3881, nx3891, 
         nx3901, nx3911, nx3921, nx3931, nx3941, nx3951, nx3961, nx3971, nx3981, 
         nx3991, nx4001, nx4011, nx4021, nx4031, nx4041, nx4051, nx4061, nx4071, 
         nx4081, nx4091, nx4101, nx4111, nx4121, nx4131, nx4141, nx4151, nx4161, 
         nx4171, nx4181, nx4191, nx4201, nx4211, nx4221, nx4231, nx4241, nx4251, 
         nx4261, nx4271, nx4281, nx4291, nx4301, nx4311, nx4321, nx4331, nx4341, 
         nx4351, nx4361, nx4371, nx4381, nx4391, nx4401, nx4411, nx4421, nx4431, 
         nx4441, nx4451, nx4461, nx4471, nx4481, nx4491, nx4501, nx4511, nx4521, 
         nx4531, nx4541, nx4551, nx4561, nx4571, nx4581, nx4591, nx4601, nx4611, 
         nx4621, nx4631, nx4641, nx4651, nx4661, nx4671, nx4681, nx4691, nx4701, 
         nx4711, nx4721, nx4731, nx4741, nx4751, nx4761, nx4771, nx4781, nx4791, 
         nx4801, nx4811, nx4821, nx4831, nx4841, nx4851, nx4861, nx4871, nx4881, 
         nx4891, nx4901, nx4911, nx4921, nx4931, nx4941, nx4951, nx4961, nx4971, 
         nx4981, nx4991, nx5001, nx5011, nx5021, nx5031, nx5041, nx5051, nx5061, 
         nx5071, nx5081, nx5091, nx5101, nx5111, nx5121, nx5131, nx5141, nx5151, 
         nx5161, nx5171, nx5181, nx5191, nx5201, nx5211, nx5221, nx5231, nx5241, 
         nx5251, nx5261, nx5271, nx5281, nx5291, nx5301, nx5311, nx5321, nx5331, 
         nx5341, nx5351, nx5361, nx5371, nx5381, nx5391, nx5401, nx5411, nx5421, 
         nx5431, nx5441, nx5451, nx5461, nx5471, nx5481, nx5491, nx5501, nx5511, 
         nx5521, nx5531, nx5541, nx5551, nx5561, nx5571, nx5581, nx5591, nx5601, 
         nx5611, nx5621, nx5631, nx5641, nx5651, nx5661, nx5671, nx5681, nx5691, 
         nx5701, nx5711, nx5721, nx5731, nx5741, nx5751, nx5761, nx5771, nx5781, 
         nx5791, nx5801, nx5811, nx5821, nx5831, nx5841, nx5851, nx5861, nx5871, 
         nx5881, nx5891, nx5901, nx5911, nx5921, nx5931, nx5941, nx5951, nx5961, 
         nx5971, nx6008, nx6075, nx6149, nx6152, nx6156, nx6158, nx6162, nx6164, 
         nx6168, nx6170, nx6174, nx6176, nx6180, nx6182, nx6186, nx6188, nx6192, 
         nx6194, nx6198, nx6200, nx6204, nx6206, nx6210, nx6212, nx6216, nx6218, 
         nx6222, nx6224, nx6228, nx6230, nx6234, nx6236, nx6240, nx6242, nx6318, 
         nx6320, nx6324, nx6326, nx6330, nx6332, nx6336, nx6338, nx6342, nx6344, 
         nx6348, nx6350, nx6354, nx6356, nx6360, nx6362, nx6366, nx6368, nx6372, 
         nx6374, nx6378, nx6380, nx6384, nx6386, nx6390, nx6392, nx6396, nx6398, 
         nx6402, nx6404, nx6408, nx6410, nx6486, nx6488, nx6492, nx6494, nx6498, 
         nx6500, nx6504, nx6506, nx6510, nx6512, nx6516, nx6518, nx6522, nx6524, 
         nx6528, nx6530, nx6534, nx6536, nx6540, nx6542, nx6546, nx6548, nx6552, 
         nx6554, nx6558, nx6560, nx6564, nx6566, nx6570, nx6572, nx6576, nx6578, 
         nx6582, nx6584, nx6588, nx6590, nx6594, nx6596, nx6600, nx6602, nx6606, 
         nx6608, nx6612, nx6614, nx6618, nx6620, nx6624, nx6626, nx6630, nx6632, 
         nx6636, nx6638, nx6642, nx6644, nx6648, nx6650, nx6654, nx6656, nx6660, 
         nx6662, nx6666, nx6668, nx6672, nx6674, nx6678, nx6680, nx6684, nx6686, 
         nx6690, nx6692, nx6696, nx6698, nx6702, nx6704, nx6708, nx6710, nx6714, 
         nx6716, nx6720, nx6722, nx6726, nx6728, nx6732, nx6734, nx6738, nx6740, 
         nx6744, nx6746, nx6750, nx6752, nx6756, nx6758, nx6762, nx6764, nx6768, 
         nx6770, nx6774, nx6776, nx6780, nx6782, nx6786, nx6788, nx6792, nx6794, 
         nx6798, nx6800, nx6804, nx6806, nx6810, nx6812, nx6816, nx6818, nx6822, 
         nx6824, nx6828, nx6830, nx6834, nx6836, nx6840, nx6842, nx6846, nx6848, 
         nx6852, nx6854, nx6858, nx6860, nx6864, nx6866, nx6870, nx6872, nx6876, 
         nx6878, nx6882, nx6884, nx6888, nx6890, nx6894, nx6896, nx6900, nx6902, 
         nx6906, nx6908, nx6912, nx6914, nx6918, nx6920, nx6924, nx6926, nx6930, 
         nx6932, nx6936, nx6938, nx6942, nx6944, nx6948, nx6950, nx6954, nx6956, 
         nx6960, nx6962, nx6966, nx7016, nx7090, nx7093, nx7097, nx7099, nx7103, 
         nx7105, nx7109, nx7111, nx7115, nx7117, nx7121, nx7123, nx7127, nx7129, 
         nx7133, nx7135, nx7139, nx7141, nx7145, nx7147, nx7151, nx7153, nx7157, 
         nx7159, nx7163, nx7165, nx7169, nx7171, nx7175, nx7177, nx7181, nx7183, 
         nx7259, nx7261, nx7265, nx7267, nx7271, nx7273, nx7277, nx7279, nx7283, 
         nx7285, nx7289, nx7291, nx7295, nx7297, nx7301, nx7303, nx7307, nx7309, 
         nx7313, nx7315, nx7319, nx7321, nx7325, nx7327, nx7331, nx7333, nx7337, 
         nx7339, nx7343, nx7345, nx7349, nx7351, nx7427, nx7429, nx7433, nx7435, 
         nx7439, nx7441, nx7445, nx7447, nx7451, nx7453, nx7457, nx7459, nx7463, 
         nx7465, nx7469, nx7471, nx7475, nx7477, nx7481, nx7483, nx7487, nx7489, 
         nx7493, nx7495, nx7499, nx7501, nx7505, nx7507, nx7511, nx7513, nx7517, 
         nx7519, nx7523, nx7525, nx7529, nx7531, nx7535, nx7537, nx7541, nx7543, 
         nx7547, nx7549, nx7553, nx7555, nx7559, nx7561, nx7565, nx7567, nx7571, 
         nx7573, nx7577, nx7579, nx7583, nx7585, nx7589, nx7591, nx7595, nx7597, 
         nx7601, nx7603, nx7607, nx7609, nx7613, nx7615, nx7619, nx7621, nx7625, 
         nx7627, nx7631, nx7633, nx7637, nx7639, nx7643, nx7645, nx7649, nx7651, 
         nx7655, nx7657, nx7661, nx7663, nx7667, nx7669, nx7673, nx7675, nx7679, 
         nx7681, nx7685, nx7687, nx7691, nx7693, nx7697, nx7699, nx7703, nx7705, 
         nx7709, nx7711, nx7715, nx7717, nx7721, nx7723, nx7727, nx7729, nx7733, 
         nx7735, nx7739, nx7741, nx7745, nx7747, nx7751, nx7753, nx7757, nx7759, 
         nx7763, nx7765, nx7769, nx7771, nx7775, nx7777, nx7781, nx7783, nx7787, 
         nx7789, nx7793, nx7795, nx7799, nx7801, nx7805, nx7807, nx7811, nx7813, 
         nx7817, nx7819, nx7823, nx7825, nx7829, nx7831, nx7835, nx7837, nx7841, 
         nx7843, nx7847, nx7849, nx7853, nx7855, nx7859, nx7861, nx7865, nx7867, 
         nx7871, nx7873, nx7877, nx7879, nx7883, nx7885, nx7889, nx7891, nx7895, 
         nx7897, nx7901, nx7903, nx7910, nx7912, nx7914, nx7916, nx7918, nx7920, 
         nx7922, nx7924, nx7926, nx7928, nx7930, nx7932, nx7934, nx7936, nx7938, 
         nx7940, nx7942, nx7944, nx7946, nx7948, nx7950, nx7952, nx7954, nx7956, 
         nx7958, nx7960, nx7962, nx7964, nx7966, nx7968, nx7970, nx7972, nx7974, 
         nx7976, nx7978, nx7980, nx7982, nx7984, nx7986, nx7988, nx7990, nx7992, 
         nx7994, nx7996, nx7998, nx8000, nx8002, nx8004, nx8006, nx8008, nx8010, 
         nx8012, nx8014, nx8016, nx8018, nx8020, nx8022, nx8024, nx8026, nx8028, 
         nx8030, nx8032, nx8034, nx8036, nx8042, nx8044, nx8046, nx8048, nx8050, 
         nx8052, nx8054, nx8056, nx8058, nx8060, nx8062, nx8064, nx8066, nx8068, 
         nx8070, nx8074, nx8076, nx8078, nx8080, nx8086, nx8088, nx8090, nx8092, 
         nx8104, nx8106, nx8108, nx8110, nx8112, nx8114, nx8116, nx8118, nx8120, 
         nx8122, nx8126, nx8128, nx8130, nx8132, nx8134, nx8138, nx8140, nx8142, 
         nx8144, nx8160, nx8162, nx8164, nx8166, nx8168, nx8170, nx8172, nx8174, 
         nx8176, nx8178, nx8180, nx8186, nx8188, nx8190, nx8192, nx8194, nx8198, 
         nx8200, nx8202, nx8204, nx8206, nx8208, nx8210, nx8212, nx8214, nx8216, 
         nx8218, nx8220, nx8222, nx8224, nx8226, nx8236, nx8238, nx8240, nx8242, 
         nx8244, nx8246, nx8248, nx8250, nx8252, nx8254, nx8256, nx8258, nx8260, 
         nx8262, nx8264, nx8266, nx8268, nx8270, nx8272, nx8274, nx8276, nx8278, 
         nx8280, nx8282, nx8284, nx8286, nx8288, nx8290, nx8292, nx8294, nx8300, 
         nx8302;
    wire [183:0] \$dummy ;




    dff RESULT_REG_reg_Dout_0 (.Q (ResultDout[0]), .QB (\$dummy [0]), .D (nx1897
        ), .CLK (CLK)) ;
    nor02ii ix1898 (.Y (nx1897), .A0 (RST), .A1 (ResultDout[0])) ;
    dff RESULT_REG_reg_Dout_1 (.Q (ResultDout[1]), .QB (\$dummy [1]), .D (nx1907
        ), .CLK (CLK)) ;
    nor02ii ix1908 (.Y (nx1907), .A0 (RST), .A1 (ResultDout[1])) ;
    dff RESULT_REG_reg_Dout_2 (.Q (ResultDout[2]), .QB (\$dummy [2]), .D (nx1917
        ), .CLK (CLK)) ;
    nor02ii ix1918 (.Y (nx1917), .A0 (RST), .A1 (ResultDout[2])) ;
    dff RESULT_REG_reg_Dout_3 (.Q (ResultDout[3]), .QB (\$dummy [3]), .D (nx1927
        ), .CLK (CLK)) ;
    nor02ii ix1928 (.Y (nx1927), .A0 (RST), .A1 (ResultDout[3])) ;
    dff RESULT_REG_reg_Dout_4 (.Q (ResultDout[4]), .QB (\$dummy [4]), .D (nx1937
        ), .CLK (CLK)) ;
    nor02ii ix1938 (.Y (nx1937), .A0 (RST), .A1 (ResultDout[4])) ;
    dff RESULT_REG_reg_Dout_5 (.Q (ResultDout[5]), .QB (\$dummy [5]), .D (nx1947
        ), .CLK (CLK)) ;
    nor02ii ix1948 (.Y (nx1947), .A0 (RST), .A1 (ResultDout[5])) ;
    dff RESULT_REG_reg_Dout_6 (.Q (ResultDout[6]), .QB (\$dummy [6]), .D (nx1957
        ), .CLK (CLK)) ;
    nor02ii ix1958 (.Y (nx1957), .A0 (RST), .A1 (ResultDout[6])) ;
    dff RESULT_REG_reg_Dout_7 (.Q (ResultDout[7]), .QB (\$dummy [7]), .D (nx1967
        ), .CLK (CLK)) ;
    nor02ii ix1968 (.Y (nx1967), .A0 (RST), .A1 (ResultDout[7])) ;
    dff L0_4_L1_4_Wij_reg_Dout_0 (.Q (WindowDout_4__4__0), .QB (\$dummy [8]), .D (
        nx1981), .CLK (CLK)) ;
    nor02ii ix87 (.Y (nx86), .A0 (RST), .A1 (Din[32])) ;
    aoi21 ix6009 (.Y (nx6008), .A0 (WindowWR), .A1 (FilterSize), .B0 (RST)) ;
    dff L0_4_L1_4_Wij_reg_Dout_1 (.Q (WindowDout_4__4__1), .QB (\$dummy [9]), .D (
        nx1991), .CLK (CLK)) ;
    nor02ii ix97 (.Y (nx96), .A0 (RST), .A1 (Din[33])) ;
    dff L0_4_L1_4_Wij_reg_Dout_2 (.Q (WindowDout_4__4__2), .QB (\$dummy [10]), .D (
        nx2001), .CLK (CLK)) ;
    nor02ii ix107 (.Y (nx106), .A0 (RST), .A1 (Din[34])) ;
    dff L0_4_L1_4_Wij_reg_Dout_3 (.Q (WindowDout_4__4__3), .QB (\$dummy [11]), .D (
        nx2011), .CLK (CLK)) ;
    nor02ii ix117 (.Y (nx116), .A0 (RST), .A1 (Din[35])) ;
    dff L0_4_L1_4_Wij_reg_Dout_4 (.Q (WindowDout_4__4__4), .QB (\$dummy [12]), .D (
        nx2021), .CLK (CLK)) ;
    nor02ii ix127 (.Y (nx126), .A0 (RST), .A1 (Din[36])) ;
    dff L0_4_L1_4_Wij_reg_Dout_5 (.Q (WindowDout_4__4__5), .QB (\$dummy [13]), .D (
        nx2031), .CLK (CLK)) ;
    nor02ii ix137 (.Y (nx136), .A0 (RST), .A1 (Din[37])) ;
    dff L0_4_L1_4_Wij_reg_Dout_6 (.Q (WindowDout_4__4__6), .QB (\$dummy [14]), .D (
        nx2041), .CLK (CLK)) ;
    nor02ii ix147 (.Y (nx146), .A0 (RST), .A1 (Din[38])) ;
    dff L0_4_L1_4_Wij_reg_Dout_7 (.Q (WindowDout_4__4__7), .QB (\$dummy [15]), .D (
        nx2051), .CLK (CLK)) ;
    nor02ii ix157 (.Y (nx156), .A0 (RST), .A1 (Din[39])) ;
    dff L0_4_L1_3_Wij_reg_Dout_0 (.Q (WindowDout_4__3__0), .QB (\$dummy [16]), .D (
        nx2141), .CLK (CLK)) ;
    nor02ii ix219 (.Y (nx218), .A0 (RST), .A1 (Din[24])) ;
    dff L0_4_L1_3_Wij_reg_Dout_1 (.Q (WindowDout_4__3__1), .QB (\$dummy [17]), .D (
        nx2151), .CLK (CLK)) ;
    nor02ii ix229 (.Y (nx228), .A0 (RST), .A1 (Din[25])) ;
    dff L0_4_L1_3_Wij_reg_Dout_2 (.Q (WindowDout_4__3__2), .QB (\$dummy [18]), .D (
        nx2161), .CLK (CLK)) ;
    nor02ii ix239 (.Y (nx238), .A0 (RST), .A1 (Din[26])) ;
    dff L0_4_L1_3_Wij_reg_Dout_3 (.Q (WindowDout_4__3__3), .QB (\$dummy [19]), .D (
        nx2171), .CLK (CLK)) ;
    nor02ii ix249 (.Y (nx248), .A0 (RST), .A1 (Din[27])) ;
    dff L0_4_L1_3_Wij_reg_Dout_4 (.Q (WindowDout_4__3__4), .QB (\$dummy [20]), .D (
        nx2181), .CLK (CLK)) ;
    nor02ii ix259 (.Y (nx258), .A0 (RST), .A1 (Din[28])) ;
    dff L0_4_L1_3_Wij_reg_Dout_5 (.Q (WindowDout_4__3__5), .QB (\$dummy [21]), .D (
        nx2191), .CLK (CLK)) ;
    nor02ii ix269 (.Y (nx268), .A0 (RST), .A1 (Din[29])) ;
    dff L0_4_L1_3_Wij_reg_Dout_6 (.Q (WindowDout_4__3__6), .QB (\$dummy [22]), .D (
        nx2201), .CLK (CLK)) ;
    nor02ii ix279 (.Y (nx278), .A0 (RST), .A1 (Din[30])) ;
    dff L0_4_L1_3_Wij_reg_Dout_7 (.Q (WindowDout_4__3__7), .QB (\$dummy [23]), .D (
        nx2211), .CLK (CLK)) ;
    nor02ii ix289 (.Y (nx288), .A0 (RST), .A1 (Din[31])) ;
    dff L0_4_L1_2_Wij_reg_Dout_0 (.Q (WindowDout_4__2__0), .QB (\$dummy [24]), .D (
        nx2301), .CLK (CLK)) ;
    ao32 ix2302 (.Y (nx2301), .A0 (Din[16]), .A1 (nx8052), .A2 (WindowWR), .B0 (
         WindowDout_4__2__0), .B1 (nx8160)) ;
    nor02_2x ix6076 (.Y (nx6075), .A0 (WindowWR), .A1 (RST)) ;
    dff L0_4_L1_2_Wij_reg_Dout_1 (.Q (WindowDout_4__2__1), .QB (\$dummy [25]), .D (
        nx2311), .CLK (CLK)) ;
    ao32 ix2312 (.Y (nx2311), .A0 (Din[17]), .A1 (nx8052), .A2 (WindowWR), .B0 (
         WindowDout_4__2__1), .B1 (nx8160)) ;
    dff L0_4_L1_2_Wij_reg_Dout_2 (.Q (WindowDout_4__2__2), .QB (\$dummy [26]), .D (
        nx2321), .CLK (CLK)) ;
    ao32 ix2322 (.Y (nx2321), .A0 (Din[18]), .A1 (nx8052), .A2 (WindowWR), .B0 (
         WindowDout_4__2__2), .B1 (nx8160)) ;
    dff L0_4_L1_2_Wij_reg_Dout_3 (.Q (WindowDout_4__2__3), .QB (\$dummy [27]), .D (
        nx2331), .CLK (CLK)) ;
    ao32 ix2332 (.Y (nx2331), .A0 (Din[19]), .A1 (nx8052), .A2 (WindowWR), .B0 (
         WindowDout_4__2__3), .B1 (nx8160)) ;
    dff L0_4_L1_2_Wij_reg_Dout_4 (.Q (WindowDout_4__2__4), .QB (\$dummy [28]), .D (
        nx2341), .CLK (CLK)) ;
    ao32 ix2342 (.Y (nx2341), .A0 (Din[20]), .A1 (nx8052), .A2 (WindowWR), .B0 (
         WindowDout_4__2__4), .B1 (nx8160)) ;
    dff L0_4_L1_2_Wij_reg_Dout_5 (.Q (WindowDout_4__2__5), .QB (\$dummy [29]), .D (
        nx2351), .CLK (CLK)) ;
    ao32 ix2352 (.Y (nx2351), .A0 (Din[21]), .A1 (nx8052), .A2 (WindowWR), .B0 (
         WindowDout_4__2__5), .B1 (nx8160)) ;
    dff L0_4_L1_2_Wij_reg_Dout_6 (.Q (WindowDout_4__2__6), .QB (\$dummy [30]), .D (
        nx2361), .CLK (CLK)) ;
    ao32 ix2362 (.Y (nx2361), .A0 (Din[22]), .A1 (nx8052), .A2 (WindowWR), .B0 (
         WindowDout_4__2__6), .B1 (nx8160)) ;
    dff L0_4_L1_2_Wij_reg_Dout_7 (.Q (WindowDout_4__2__7), .QB (\$dummy [31]), .D (
        nx2371), .CLK (CLK)) ;
    ao32 ix2372 (.Y (nx2371), .A0 (Din[23]), .A1 (nx8054), .A2 (WindowWR), .B0 (
         WindowDout_4__2__7), .B1 (nx8162)) ;
    dff L0_4_L1_1_Wij_reg_Dout_0 (.Q (WindowDout_4__1__0), .QB (\$dummy [32]), .D (
        nx2461), .CLK (CLK)) ;
    ao32 ix2462 (.Y (nx2461), .A0 (Din[8]), .A1 (nx8054), .A2 (WindowWR), .B0 (
         WindowDout_4__1__0), .B1 (nx8162)) ;
    dff L0_4_L1_1_Wij_reg_Dout_1 (.Q (WindowDout_4__1__1), .QB (\$dummy [33]), .D (
        nx2471), .CLK (CLK)) ;
    ao32 ix2472 (.Y (nx2471), .A0 (Din[9]), .A1 (nx8054), .A2 (WindowWR), .B0 (
         WindowDout_4__1__1), .B1 (nx8162)) ;
    dff L0_4_L1_1_Wij_reg_Dout_2 (.Q (WindowDout_4__1__2), .QB (\$dummy [34]), .D (
        nx2481), .CLK (CLK)) ;
    ao32 ix2482 (.Y (nx2481), .A0 (Din[10]), .A1 (nx8054), .A2 (WindowWR), .B0 (
         WindowDout_4__1__2), .B1 (nx8162)) ;
    dff L0_4_L1_1_Wij_reg_Dout_3 (.Q (WindowDout_4__1__3), .QB (\$dummy [35]), .D (
        nx2491), .CLK (CLK)) ;
    ao32 ix2492 (.Y (nx2491), .A0 (Din[11]), .A1 (nx8054), .A2 (WindowWR), .B0 (
         WindowDout_4__1__3), .B1 (nx8162)) ;
    dff L0_4_L1_1_Wij_reg_Dout_4 (.Q (WindowDout_4__1__4), .QB (\$dummy [36]), .D (
        nx2501), .CLK (CLK)) ;
    ao32 ix2502 (.Y (nx2501), .A0 (Din[12]), .A1 (nx8054), .A2 (WindowWR), .B0 (
         WindowDout_4__1__4), .B1 (nx8162)) ;
    dff L0_4_L1_1_Wij_reg_Dout_5 (.Q (WindowDout_4__1__5), .QB (\$dummy [37]), .D (
        nx2511), .CLK (CLK)) ;
    ao32 ix2512 (.Y (nx2511), .A0 (Din[13]), .A1 (nx8054), .A2 (WindowWR), .B0 (
         WindowDout_4__1__5), .B1 (nx8162)) ;
    dff L0_4_L1_1_Wij_reg_Dout_6 (.Q (WindowDout_4__1__6), .QB (\$dummy [38]), .D (
        nx2521), .CLK (CLK)) ;
    ao32 ix2522 (.Y (nx2521), .A0 (Din[14]), .A1 (nx8056), .A2 (WindowWR), .B0 (
         WindowDout_4__1__6), .B1 (nx8164)) ;
    dff L0_4_L1_1_Wij_reg_Dout_7 (.Q (WindowDout_4__1__7), .QB (\$dummy [39]), .D (
        nx2531), .CLK (CLK)) ;
    ao32 ix2532 (.Y (nx2531), .A0 (Din[15]), .A1 (nx8056), .A2 (WindowWR), .B0 (
         WindowDout_4__1__7), .B1 (nx8164)) ;
    dff L0_4_L1_0_Wij_reg_Dout_0 (.Q (WindowDout_4__0__0), .QB (\$dummy [40]), .D (
        nx2621), .CLK (CLK)) ;
    ao32 ix2622 (.Y (nx2621), .A0 (Din[0]), .A1 (nx8056), .A2 (WindowWR), .B0 (
         WindowDout_4__0__0), .B1 (nx8164)) ;
    dff L0_4_L1_0_Wij_reg_Dout_1 (.Q (WindowDout_4__0__1), .QB (\$dummy [41]), .D (
        nx2631), .CLK (CLK)) ;
    ao32 ix2632 (.Y (nx2631), .A0 (Din[1]), .A1 (nx8056), .A2 (WindowWR), .B0 (
         WindowDout_4__0__1), .B1 (nx8164)) ;
    dff L0_4_L1_0_Wij_reg_Dout_2 (.Q (WindowDout_4__0__2), .QB (\$dummy [42]), .D (
        nx2641), .CLK (CLK)) ;
    ao32 ix2642 (.Y (nx2641), .A0 (Din[2]), .A1 (nx8056), .A2 (WindowWR), .B0 (
         WindowDout_4__0__2), .B1 (nx8164)) ;
    dff L0_4_L1_0_Wij_reg_Dout_3 (.Q (WindowDout_4__0__3), .QB (\$dummy [43]), .D (
        nx2651), .CLK (CLK)) ;
    ao32 ix2652 (.Y (nx2651), .A0 (Din[3]), .A1 (nx8056), .A2 (WindowWR), .B0 (
         WindowDout_4__0__3), .B1 (nx8164)) ;
    dff L0_4_L1_0_Wij_reg_Dout_4 (.Q (WindowDout_4__0__4), .QB (\$dummy [44]), .D (
        nx2661), .CLK (CLK)) ;
    ao32 ix2662 (.Y (nx2661), .A0 (Din[4]), .A1 (nx8056), .A2 (WindowWR), .B0 (
         WindowDout_4__0__4), .B1 (nx8164)) ;
    dff L0_4_L1_0_Wij_reg_Dout_5 (.Q (WindowDout_4__0__5), .QB (\$dummy [45]), .D (
        nx2671), .CLK (CLK)) ;
    ao32 ix2672 (.Y (nx2671), .A0 (Din[5]), .A1 (nx8058), .A2 (WindowWR), .B0 (
         WindowDout_4__0__5), .B1 (nx8166)) ;
    dff L0_4_L1_0_Wij_reg_Dout_6 (.Q (WindowDout_4__0__6), .QB (\$dummy [46]), .D (
        nx2681), .CLK (CLK)) ;
    ao32 ix2682 (.Y (nx2681), .A0 (Din[6]), .A1 (nx8058), .A2 (WindowWR), .B0 (
         WindowDout_4__0__6), .B1 (nx8166)) ;
    dff L0_4_L1_0_Wij_reg_Dout_7 (.Q (WindowDout_4__0__7), .QB (\$dummy [47]), .D (
        nx2691), .CLK (CLK)) ;
    ao32 ix2692 (.Y (nx2691), .A0 (Din[7]), .A1 (nx8058), .A2 (WindowWR), .B0 (
         WindowDout_4__0__7), .B1 (nx8166)) ;
    oai21 ix2782 (.Y (nx2781), .A0 (nx6149), .A1 (nx7910), .B0 (nx6152)) ;
    dff L0_3_L1_4_Wij_reg_Dout_0 (.Q (WindowDout_3__4__0), .QB (nx6149), .D (
        nx2781), .CLK (CLK)) ;
    nand03 ix6153 (.Y (nx6152), .A0 (nx8058), .A1 (WindowDout_4__4__0), .A2 (
           nx7910)) ;
    oai21 ix2792 (.Y (nx2791), .A0 (nx6156), .A1 (nx7910), .B0 (nx6158)) ;
    dff L0_3_L1_4_Wij_reg_Dout_1 (.Q (WindowDout_3__4__1), .QB (nx6156), .D (
        nx2791), .CLK (CLK)) ;
    nand03 ix6159 (.Y (nx6158), .A0 (nx8058), .A1 (WindowDout_4__4__1), .A2 (
           nx7910)) ;
    oai21 ix2802 (.Y (nx2801), .A0 (nx6162), .A1 (nx7910), .B0 (nx6164)) ;
    dff L0_3_L1_4_Wij_reg_Dout_2 (.Q (WindowDout_3__4__2), .QB (nx6162), .D (
        nx2801), .CLK (CLK)) ;
    nand03 ix6165 (.Y (nx6164), .A0 (nx8058), .A1 (WindowDout_4__4__2), .A2 (
           nx7910)) ;
    oai21 ix2812 (.Y (nx2811), .A0 (nx6168), .A1 (nx7910), .B0 (nx6170)) ;
    dff L0_3_L1_4_Wij_reg_Dout_3 (.Q (WindowDout_3__4__3), .QB (nx6168), .D (
        nx2811), .CLK (CLK)) ;
    nand03 ix6171 (.Y (nx6170), .A0 (nx8058), .A1 (WindowDout_4__4__3), .A2 (
           nx7912)) ;
    oai21 ix2822 (.Y (nx2821), .A0 (nx6174), .A1 (nx7912), .B0 (nx6176)) ;
    dff L0_3_L1_4_Wij_reg_Dout_4 (.Q (WindowDout_3__4__4), .QB (nx6174), .D (
        nx2821), .CLK (CLK)) ;
    nand03 ix6177 (.Y (nx6176), .A0 (nx8060), .A1 (WindowDout_4__4__4), .A2 (
           nx7912)) ;
    oai21 ix2832 (.Y (nx2831), .A0 (nx6180), .A1 (nx7912), .B0 (nx6182)) ;
    dff L0_3_L1_4_Wij_reg_Dout_5 (.Q (WindowDout_3__4__5), .QB (nx6180), .D (
        nx2831), .CLK (CLK)) ;
    nand03 ix6183 (.Y (nx6182), .A0 (nx8060), .A1 (WindowDout_4__4__5), .A2 (
           nx7912)) ;
    oai21 ix2842 (.Y (nx2841), .A0 (nx6186), .A1 (nx7912), .B0 (nx6188)) ;
    dff L0_3_L1_4_Wij_reg_Dout_6 (.Q (WindowDout_3__4__6), .QB (nx6186), .D (
        nx2841), .CLK (CLK)) ;
    nand03 ix6189 (.Y (nx6188), .A0 (nx8060), .A1 (WindowDout_4__4__6), .A2 (
           nx7912)) ;
    oai21 ix2852 (.Y (nx2851), .A0 (nx6192), .A1 (nx7914), .B0 (nx6194)) ;
    dff L0_3_L1_4_Wij_reg_Dout_7 (.Q (WindowDout_3__4__7), .QB (nx6192), .D (
        nx2851), .CLK (CLK)) ;
    nand03 ix6195 (.Y (nx6194), .A0 (nx8060), .A1 (WindowDout_4__4__7), .A2 (
           nx7914)) ;
    oai21 ix2942 (.Y (nx2941), .A0 (nx6198), .A1 (nx7914), .B0 (nx6200)) ;
    dff L0_3_L1_3_Wij_reg_Dout_0 (.Q (WindowDout_3__3__0), .QB (nx6198), .D (
        nx2941), .CLK (CLK)) ;
    nand03 ix6201 (.Y (nx6200), .A0 (nx8060), .A1 (WindowDout_4__3__0), .A2 (
           nx7914)) ;
    oai21 ix2952 (.Y (nx2951), .A0 (nx6204), .A1 (nx7914), .B0 (nx6206)) ;
    dff L0_3_L1_3_Wij_reg_Dout_1 (.Q (WindowDout_3__3__1), .QB (nx6204), .D (
        nx2951), .CLK (CLK)) ;
    nand03 ix6207 (.Y (nx6206), .A0 (nx8060), .A1 (WindowDout_4__3__1), .A2 (
           nx7914)) ;
    oai21 ix2962 (.Y (nx2961), .A0 (nx6210), .A1 (nx7914), .B0 (nx6212)) ;
    dff L0_3_L1_3_Wij_reg_Dout_2 (.Q (WindowDout_3__3__2), .QB (nx6210), .D (
        nx2961), .CLK (CLK)) ;
    nand03 ix6213 (.Y (nx6212), .A0 (nx8060), .A1 (WindowDout_4__3__2), .A2 (
           nx7916)) ;
    oai21 ix2972 (.Y (nx2971), .A0 (nx6216), .A1 (nx7916), .B0 (nx6218)) ;
    dff L0_3_L1_3_Wij_reg_Dout_3 (.Q (WindowDout_3__3__3), .QB (nx6216), .D (
        nx2971), .CLK (CLK)) ;
    nand03 ix6219 (.Y (nx6218), .A0 (nx8062), .A1 (WindowDout_4__3__3), .A2 (
           nx7916)) ;
    oai21 ix2982 (.Y (nx2981), .A0 (nx6222), .A1 (nx7916), .B0 (nx6224)) ;
    dff L0_3_L1_3_Wij_reg_Dout_4 (.Q (WindowDout_3__3__4), .QB (nx6222), .D (
        nx2981), .CLK (CLK)) ;
    nand03 ix6225 (.Y (nx6224), .A0 (nx8062), .A1 (WindowDout_4__3__4), .A2 (
           nx7916)) ;
    oai21 ix2992 (.Y (nx2991), .A0 (nx6228), .A1 (nx7916), .B0 (nx6230)) ;
    dff L0_3_L1_3_Wij_reg_Dout_5 (.Q (WindowDout_3__3__5), .QB (nx6228), .D (
        nx2991), .CLK (CLK)) ;
    nand03 ix6231 (.Y (nx6230), .A0 (nx8062), .A1 (WindowDout_4__3__5), .A2 (
           nx7916)) ;
    oai21 ix3002 (.Y (nx3001), .A0 (nx6234), .A1 (nx7918), .B0 (nx6236)) ;
    dff L0_3_L1_3_Wij_reg_Dout_6 (.Q (WindowDout_3__3__6), .QB (nx6234), .D (
        nx3001), .CLK (CLK)) ;
    nand03 ix6237 (.Y (nx6236), .A0 (nx8062), .A1 (WindowDout_4__3__6), .A2 (
           nx7918)) ;
    oai21 ix3012 (.Y (nx3011), .A0 (nx6240), .A1 (nx7918), .B0 (nx6242)) ;
    dff L0_3_L1_3_Wij_reg_Dout_7 (.Q (WindowDout_3__3__7), .QB (nx6240), .D (
        nx3011), .CLK (CLK)) ;
    nand03 ix6243 (.Y (nx6242), .A0 (nx8062), .A1 (WindowDout_4__3__7), .A2 (
           nx7918)) ;
    dff L0_3_L1_2_Wij_reg_Dout_0 (.Q (WindowDout_3__2__0), .QB (\$dummy [48]), .D (
        nx3101), .CLK (CLK)) ;
    ao32 ix3102 (.Y (nx3101), .A0 (nx8062), .A1 (WindowDout_4__2__0), .A2 (
         WindowWR), .B0 (WindowDout_3__2__0), .B1 (nx8166)) ;
    dff L0_3_L1_2_Wij_reg_Dout_1 (.Q (WindowDout_3__2__1), .QB (\$dummy [49]), .D (
        nx3111), .CLK (CLK)) ;
    ao32 ix3112 (.Y (nx3111), .A0 (nx8062), .A1 (WindowDout_4__2__1), .A2 (
         WindowWR), .B0 (WindowDout_3__2__1), .B1 (nx8166)) ;
    dff L0_3_L1_2_Wij_reg_Dout_2 (.Q (WindowDout_3__2__2), .QB (\$dummy [50]), .D (
        nx3121), .CLK (CLK)) ;
    ao32 ix3122 (.Y (nx3121), .A0 (nx8064), .A1 (WindowDout_4__2__2), .A2 (
         WindowWR), .B0 (WindowDout_3__2__2), .B1 (nx8166)) ;
    dff L0_3_L1_2_Wij_reg_Dout_3 (.Q (WindowDout_3__2__3), .QB (\$dummy [51]), .D (
        nx3131), .CLK (CLK)) ;
    ao32 ix3132 (.Y (nx3131), .A0 (nx8064), .A1 (WindowDout_4__2__3), .A2 (
         WindowWR), .B0 (WindowDout_3__2__3), .B1 (nx8166)) ;
    dff L0_3_L1_2_Wij_reg_Dout_4 (.Q (WindowDout_3__2__4), .QB (\$dummy [52]), .D (
        nx3141), .CLK (CLK)) ;
    ao32 ix3142 (.Y (nx3141), .A0 (nx8064), .A1 (WindowDout_4__2__4), .A2 (
         WindowWR), .B0 (WindowDout_3__2__4), .B1 (nx8168)) ;
    dff L0_3_L1_2_Wij_reg_Dout_5 (.Q (WindowDout_3__2__5), .QB (\$dummy [53]), .D (
        nx3151), .CLK (CLK)) ;
    ao32 ix3152 (.Y (nx3151), .A0 (nx8064), .A1 (WindowDout_4__2__5), .A2 (
         WindowWR), .B0 (WindowDout_3__2__5), .B1 (nx8168)) ;
    dff L0_3_L1_2_Wij_reg_Dout_6 (.Q (WindowDout_3__2__6), .QB (\$dummy [54]), .D (
        nx3161), .CLK (CLK)) ;
    ao32 ix3162 (.Y (nx3161), .A0 (nx8064), .A1 (WindowDout_4__2__6), .A2 (
         WindowWR), .B0 (WindowDout_3__2__6), .B1 (nx8168)) ;
    dff L0_3_L1_2_Wij_reg_Dout_7 (.Q (WindowDout_3__2__7), .QB (\$dummy [55]), .D (
        nx3171), .CLK (CLK)) ;
    ao32 ix3172 (.Y (nx3171), .A0 (nx8064), .A1 (WindowDout_4__2__7), .A2 (
         WindowWR), .B0 (WindowDout_3__2__7), .B1 (nx8168)) ;
    dff L0_3_L1_1_Wij_reg_Dout_0 (.Q (WindowDout_3__1__0), .QB (\$dummy [56]), .D (
        nx3261), .CLK (CLK)) ;
    ao32 ix3262 (.Y (nx3261), .A0 (nx8064), .A1 (WindowDout_4__1__0), .A2 (
         WindowWR), .B0 (WindowDout_3__1__0), .B1 (nx8168)) ;
    dff L0_3_L1_1_Wij_reg_Dout_1 (.Q (WindowDout_3__1__1), .QB (\$dummy [57]), .D (
        nx3271), .CLK (CLK)) ;
    ao32 ix3272 (.Y (nx3271), .A0 (nx8066), .A1 (WindowDout_4__1__1), .A2 (
         WindowWR), .B0 (WindowDout_3__1__1), .B1 (nx8168)) ;
    dff L0_3_L1_1_Wij_reg_Dout_2 (.Q (WindowDout_3__1__2), .QB (\$dummy [58]), .D (
        nx3281), .CLK (CLK)) ;
    ao32 ix3282 (.Y (nx3281), .A0 (nx8066), .A1 (WindowDout_4__1__2), .A2 (
         WindowWR), .B0 (WindowDout_3__1__2), .B1 (nx8168)) ;
    dff L0_3_L1_1_Wij_reg_Dout_3 (.Q (WindowDout_3__1__3), .QB (\$dummy [59]), .D (
        nx3291), .CLK (CLK)) ;
    ao32 ix3292 (.Y (nx3291), .A0 (nx8066), .A1 (WindowDout_4__1__3), .A2 (
         WindowWR), .B0 (WindowDout_3__1__3), .B1 (nx8170)) ;
    dff L0_3_L1_1_Wij_reg_Dout_4 (.Q (WindowDout_3__1__4), .QB (\$dummy [60]), .D (
        nx3301), .CLK (CLK)) ;
    ao32 ix3302 (.Y (nx3301), .A0 (nx8066), .A1 (WindowDout_4__1__4), .A2 (
         WindowWR), .B0 (WindowDout_3__1__4), .B1 (nx8170)) ;
    dff L0_3_L1_1_Wij_reg_Dout_5 (.Q (WindowDout_3__1__5), .QB (\$dummy [61]), .D (
        nx3311), .CLK (CLK)) ;
    ao32 ix3312 (.Y (nx3311), .A0 (nx8066), .A1 (WindowDout_4__1__5), .A2 (
         WindowWR), .B0 (WindowDout_3__1__5), .B1 (nx8170)) ;
    dff L0_3_L1_1_Wij_reg_Dout_6 (.Q (WindowDout_3__1__6), .QB (\$dummy [62]), .D (
        nx3321), .CLK (CLK)) ;
    ao32 ix3322 (.Y (nx3321), .A0 (nx8066), .A1 (WindowDout_4__1__6), .A2 (
         WindowWR), .B0 (WindowDout_3__1__6), .B1 (nx8170)) ;
    dff L0_3_L1_1_Wij_reg_Dout_7 (.Q (WindowDout_3__1__7), .QB (\$dummy [63]), .D (
        nx3331), .CLK (CLK)) ;
    ao32 ix3332 (.Y (nx3331), .A0 (nx8066), .A1 (WindowDout_4__1__7), .A2 (
         WindowWR), .B0 (WindowDout_3__1__7), .B1 (nx8170)) ;
    dff L0_3_L1_0_Wij_reg_Dout_0 (.Q (WindowDout_3__0__0), .QB (\$dummy [64]), .D (
        nx3421), .CLK (CLK)) ;
    ao32 ix3422 (.Y (nx3421), .A0 (nx8068), .A1 (WindowDout_4__0__0), .A2 (
         WindowWR), .B0 (WindowDout_3__0__0), .B1 (nx8170)) ;
    dff L0_3_L1_0_Wij_reg_Dout_1 (.Q (WindowDout_3__0__1), .QB (\$dummy [65]), .D (
        nx3431), .CLK (CLK)) ;
    ao32 ix3432 (.Y (nx3431), .A0 (nx8068), .A1 (WindowDout_4__0__1), .A2 (
         WindowWR), .B0 (WindowDout_3__0__1), .B1 (nx8170)) ;
    dff L0_3_L1_0_Wij_reg_Dout_2 (.Q (WindowDout_3__0__2), .QB (\$dummy [66]), .D (
        nx3441), .CLK (CLK)) ;
    ao32 ix3442 (.Y (nx3441), .A0 (nx8068), .A1 (WindowDout_4__0__2), .A2 (
         WindowWR), .B0 (WindowDout_3__0__2), .B1 (nx8172)) ;
    dff L0_3_L1_0_Wij_reg_Dout_3 (.Q (WindowDout_3__0__3), .QB (\$dummy [67]), .D (
        nx3451), .CLK (CLK)) ;
    ao32 ix3452 (.Y (nx3451), .A0 (nx8068), .A1 (WindowDout_4__0__3), .A2 (
         WindowWR), .B0 (WindowDout_3__0__3), .B1 (nx8172)) ;
    dff L0_3_L1_0_Wij_reg_Dout_4 (.Q (WindowDout_3__0__4), .QB (\$dummy [68]), .D (
        nx3461), .CLK (CLK)) ;
    ao32 ix3462 (.Y (nx3461), .A0 (nx8068), .A1 (WindowDout_4__0__4), .A2 (
         WindowWR), .B0 (WindowDout_3__0__4), .B1 (nx8172)) ;
    dff L0_3_L1_0_Wij_reg_Dout_5 (.Q (WindowDout_3__0__5), .QB (\$dummy [69]), .D (
        nx3471), .CLK (CLK)) ;
    ao32 ix3472 (.Y (nx3471), .A0 (nx8068), .A1 (WindowDout_4__0__5), .A2 (
         WindowWR), .B0 (WindowDout_3__0__5), .B1 (nx8172)) ;
    dff L0_3_L1_0_Wij_reg_Dout_6 (.Q (WindowDout_3__0__6), .QB (\$dummy [70]), .D (
        nx3481), .CLK (CLK)) ;
    ao32 ix3482 (.Y (nx3481), .A0 (nx8068), .A1 (WindowDout_4__0__6), .A2 (
         WindowWR), .B0 (WindowDout_3__0__6), .B1 (nx8172)) ;
    dff L0_3_L1_0_Wij_reg_Dout_7 (.Q (WindowDout_3__0__7), .QB (\$dummy [71]), .D (
        nx3491), .CLK (CLK)) ;
    ao32 ix3492 (.Y (nx3491), .A0 (nx8070), .A1 (WindowDout_4__0__7), .A2 (
         WindowWR), .B0 (WindowDout_3__0__7), .B1 (nx8172)) ;
    oai21 ix3582 (.Y (nx3581), .A0 (nx6318), .A1 (nx7918), .B0 (nx6320)) ;
    dff L0_2_L1_4_Wij_reg_Dout_0 (.Q (WindowDout_2__4__0), .QB (nx6318), .D (
        nx3581), .CLK (CLK)) ;
    oai21 ix3592 (.Y (nx3591), .A0 (nx6324), .A1 (nx7918), .B0 (nx6326)) ;
    dff L0_2_L1_4_Wij_reg_Dout_1 (.Q (WindowDout_2__4__1), .QB (nx6324), .D (
        nx3591), .CLK (CLK)) ;
    oai21 ix3602 (.Y (nx3601), .A0 (nx6330), .A1 (nx7920), .B0 (nx6332)) ;
    dff L0_2_L1_4_Wij_reg_Dout_2 (.Q (WindowDout_2__4__2), .QB (nx6330), .D (
        nx3601), .CLK (CLK)) ;
    oai21 ix3612 (.Y (nx3611), .A0 (nx6336), .A1 (nx7920), .B0 (nx6338)) ;
    dff L0_2_L1_4_Wij_reg_Dout_3 (.Q (WindowDout_2__4__3), .QB (nx6336), .D (
        nx3611), .CLK (CLK)) ;
    oai21 ix3622 (.Y (nx3621), .A0 (nx6342), .A1 (nx7920), .B0 (nx6344)) ;
    dff L0_2_L1_4_Wij_reg_Dout_4 (.Q (WindowDout_2__4__4), .QB (nx6342), .D (
        nx3621), .CLK (CLK)) ;
    oai21 ix3632 (.Y (nx3631), .A0 (nx6348), .A1 (nx7922), .B0 (nx6350)) ;
    dff L0_2_L1_4_Wij_reg_Dout_5 (.Q (WindowDout_2__4__5), .QB (nx6348), .D (
        nx3631), .CLK (CLK)) ;
    oai21 ix3642 (.Y (nx3641), .A0 (nx6354), .A1 (nx7922), .B0 (nx6356)) ;
    dff L0_2_L1_4_Wij_reg_Dout_6 (.Q (WindowDout_2__4__6), .QB (nx6354), .D (
        nx3641), .CLK (CLK)) ;
    oai21 ix3652 (.Y (nx3651), .A0 (nx6360), .A1 (nx7922), .B0 (nx6362)) ;
    dff L0_2_L1_4_Wij_reg_Dout_7 (.Q (WindowDout_2__4__7), .QB (nx6360), .D (
        nx3651), .CLK (CLK)) ;
    oai21 ix3742 (.Y (nx3741), .A0 (nx6366), .A1 (nx7922), .B0 (nx6368)) ;
    dff L0_2_L1_3_Wij_reg_Dout_0 (.Q (WindowDout_2__3__0), .QB (nx6366), .D (
        nx3741), .CLK (CLK)) ;
    oai21 ix3752 (.Y (nx3751), .A0 (nx6372), .A1 (nx7924), .B0 (nx6374)) ;
    dff L0_2_L1_3_Wij_reg_Dout_1 (.Q (WindowDout_2__3__1), .QB (nx6372), .D (
        nx3751), .CLK (CLK)) ;
    oai21 ix3762 (.Y (nx3761), .A0 (nx6378), .A1 (nx7924), .B0 (nx6380)) ;
    dff L0_2_L1_3_Wij_reg_Dout_2 (.Q (WindowDout_2__3__2), .QB (nx6378), .D (
        nx3761), .CLK (CLK)) ;
    oai21 ix3772 (.Y (nx3771), .A0 (nx6384), .A1 (nx7924), .B0 (nx6386)) ;
    dff L0_2_L1_3_Wij_reg_Dout_3 (.Q (WindowDout_2__3__3), .QB (nx6384), .D (
        nx3771), .CLK (CLK)) ;
    oai21 ix3782 (.Y (nx3781), .A0 (nx6390), .A1 (nx7926), .B0 (nx6392)) ;
    dff L0_2_L1_3_Wij_reg_Dout_4 (.Q (WindowDout_2__3__4), .QB (nx6390), .D (
        nx3781), .CLK (CLK)) ;
    oai21 ix3792 (.Y (nx3791), .A0 (nx6396), .A1 (nx7926), .B0 (nx6398)) ;
    dff L0_2_L1_3_Wij_reg_Dout_5 (.Q (WindowDout_2__3__5), .QB (nx6396), .D (
        nx3791), .CLK (CLK)) ;
    oai21 ix3802 (.Y (nx3801), .A0 (nx6402), .A1 (nx7926), .B0 (nx6404)) ;
    dff L0_2_L1_3_Wij_reg_Dout_6 (.Q (WindowDout_2__3__6), .QB (nx6402), .D (
        nx3801), .CLK (CLK)) ;
    oai21 ix3812 (.Y (nx3811), .A0 (nx6408), .A1 (nx7926), .B0 (nx6410)) ;
    dff L0_2_L1_3_Wij_reg_Dout_7 (.Q (WindowDout_2__3__7), .QB (nx6408), .D (
        nx3811), .CLK (CLK)) ;
    dff L0_2_L1_2_Wij_reg_Dout_0 (.Q (WindowDout_2__2__0), .QB (\$dummy [72]), .D (
        nx3901), .CLK (CLK)) ;
    ao32 ix3902 (.Y (nx3901), .A0 (nx8074), .A1 (WindowDout_3__2__0), .A2 (
         WindowWR), .B0 (WindowDout_2__2__0), .B1 (nx8172)) ;
    dff L0_2_L1_2_Wij_reg_Dout_1 (.Q (WindowDout_2__2__1), .QB (\$dummy [73]), .D (
        nx3911), .CLK (CLK)) ;
    ao32 ix3912 (.Y (nx3911), .A0 (nx8074), .A1 (WindowDout_3__2__1), .A2 (
         WindowWR), .B0 (WindowDout_2__2__1), .B1 (nx8174)) ;
    dff L0_2_L1_2_Wij_reg_Dout_2 (.Q (WindowDout_2__2__2), .QB (\$dummy [74]), .D (
        nx3921), .CLK (CLK)) ;
    ao32 ix3922 (.Y (nx3921), .A0 (nx8074), .A1 (WindowDout_3__2__2), .A2 (
         WindowWR), .B0 (WindowDout_2__2__2), .B1 (nx8174)) ;
    dff L0_2_L1_2_Wij_reg_Dout_3 (.Q (WindowDout_2__2__3), .QB (\$dummy [75]), .D (
        nx3931), .CLK (CLK)) ;
    ao32 ix3932 (.Y (nx3931), .A0 (nx8074), .A1 (WindowDout_3__2__3), .A2 (
         WindowWR), .B0 (WindowDout_2__2__3), .B1 (nx8174)) ;
    dff L0_2_L1_2_Wij_reg_Dout_4 (.Q (WindowDout_2__2__4), .QB (\$dummy [76]), .D (
        nx3941), .CLK (CLK)) ;
    ao32 ix3942 (.Y (nx3941), .A0 (nx8076), .A1 (WindowDout_3__2__4), .A2 (
         WindowWR), .B0 (WindowDout_2__2__4), .B1 (nx8174)) ;
    dff L0_2_L1_2_Wij_reg_Dout_5 (.Q (WindowDout_2__2__5), .QB (\$dummy [77]), .D (
        nx3951), .CLK (CLK)) ;
    ao32 ix3952 (.Y (nx3951), .A0 (nx8076), .A1 (WindowDout_3__2__5), .A2 (
         WindowWR), .B0 (WindowDout_2__2__5), .B1 (nx8174)) ;
    dff L0_2_L1_2_Wij_reg_Dout_6 (.Q (WindowDout_2__2__6), .QB (\$dummy [78]), .D (
        nx3961), .CLK (CLK)) ;
    ao32 ix3962 (.Y (nx3961), .A0 (nx8076), .A1 (WindowDout_3__2__6), .A2 (
         WindowWR), .B0 (WindowDout_2__2__6), .B1 (nx8174)) ;
    dff L0_2_L1_2_Wij_reg_Dout_7 (.Q (WindowDout_2__2__7), .QB (\$dummy [79]), .D (
        nx3971), .CLK (CLK)) ;
    ao32 ix3972 (.Y (nx3971), .A0 (nx8076), .A1 (WindowDout_3__2__7), .A2 (
         WindowWR), .B0 (WindowDout_2__2__7), .B1 (nx8174)) ;
    dff L0_2_L1_1_Wij_reg_Dout_0 (.Q (WindowDout_2__1__0), .QB (\$dummy [80]), .D (
        nx4061), .CLK (CLK)) ;
    ao32 ix4062 (.Y (nx4061), .A0 (nx8076), .A1 (WindowDout_3__1__0), .A2 (
         WindowWR), .B0 (WindowDout_2__1__0), .B1 (nx8176)) ;
    dff L0_2_L1_1_Wij_reg_Dout_1 (.Q (WindowDout_2__1__1), .QB (\$dummy [81]), .D (
        nx4071), .CLK (CLK)) ;
    ao32 ix4072 (.Y (nx4071), .A0 (nx8076), .A1 (WindowDout_3__1__1), .A2 (
         WindowWR), .B0 (WindowDout_2__1__1), .B1 (nx8176)) ;
    dff L0_2_L1_1_Wij_reg_Dout_2 (.Q (WindowDout_2__1__2), .QB (\$dummy [82]), .D (
        nx4081), .CLK (CLK)) ;
    ao32 ix4082 (.Y (nx4081), .A0 (nx8076), .A1 (WindowDout_3__1__2), .A2 (
         WindowWR), .B0 (WindowDout_2__1__2), .B1 (nx8176)) ;
    dff L0_2_L1_1_Wij_reg_Dout_3 (.Q (WindowDout_2__1__3), .QB (\$dummy [83]), .D (
        nx4091), .CLK (CLK)) ;
    ao32 ix4092 (.Y (nx4091), .A0 (nx8078), .A1 (WindowDout_3__1__3), .A2 (
         WindowWR), .B0 (WindowDout_2__1__3), .B1 (nx8176)) ;
    dff L0_2_L1_1_Wij_reg_Dout_4 (.Q (WindowDout_2__1__4), .QB (\$dummy [84]), .D (
        nx4101), .CLK (CLK)) ;
    ao32 ix4102 (.Y (nx4101), .A0 (nx8078), .A1 (WindowDout_3__1__4), .A2 (
         WindowWR), .B0 (WindowDout_2__1__4), .B1 (nx8176)) ;
    dff L0_2_L1_1_Wij_reg_Dout_5 (.Q (WindowDout_2__1__5), .QB (\$dummy [85]), .D (
        nx4111), .CLK (CLK)) ;
    ao32 ix4112 (.Y (nx4111), .A0 (nx8078), .A1 (WindowDout_3__1__5), .A2 (
         WindowWR), .B0 (WindowDout_2__1__5), .B1 (nx8176)) ;
    dff L0_2_L1_1_Wij_reg_Dout_6 (.Q (WindowDout_2__1__6), .QB (\$dummy [86]), .D (
        nx4121), .CLK (CLK)) ;
    ao32 ix4122 (.Y (nx4121), .A0 (nx8078), .A1 (WindowDout_3__1__6), .A2 (
         WindowWR), .B0 (WindowDout_2__1__6), .B1 (nx8176)) ;
    dff L0_2_L1_1_Wij_reg_Dout_7 (.Q (WindowDout_2__1__7), .QB (\$dummy [87]), .D (
        nx4131), .CLK (CLK)) ;
    ao32 ix4132 (.Y (nx4131), .A0 (nx8078), .A1 (WindowDout_3__1__7), .A2 (
         WindowWR), .B0 (WindowDout_2__1__7), .B1 (nx8178)) ;
    dff L0_2_L1_0_Wij_reg_Dout_0 (.Q (WindowDout_2__0__0), .QB (\$dummy [88]), .D (
        nx4221), .CLK (CLK)) ;
    ao32 ix4222 (.Y (nx4221), .A0 (nx8078), .A1 (WindowDout_3__0__0), .A2 (
         WindowWR), .B0 (WindowDout_2__0__0), .B1 (nx8178)) ;
    dff L0_2_L1_0_Wij_reg_Dout_1 (.Q (WindowDout_2__0__1), .QB (\$dummy [89]), .D (
        nx4231), .CLK (CLK)) ;
    ao32 ix4232 (.Y (nx4231), .A0 (nx8078), .A1 (WindowDout_3__0__1), .A2 (
         WindowWR), .B0 (WindowDout_2__0__1), .B1 (nx8178)) ;
    dff L0_2_L1_0_Wij_reg_Dout_2 (.Q (WindowDout_2__0__2), .QB (\$dummy [90]), .D (
        nx4241), .CLK (CLK)) ;
    ao32 ix4242 (.Y (nx4241), .A0 (nx8080), .A1 (WindowDout_3__0__2), .A2 (
         WindowWR), .B0 (WindowDout_2__0__2), .B1 (nx8178)) ;
    dff L0_2_L1_0_Wij_reg_Dout_3 (.Q (WindowDout_2__0__3), .QB (\$dummy [91]), .D (
        nx4251), .CLK (CLK)) ;
    ao32 ix4252 (.Y (nx4251), .A0 (nx8080), .A1 (WindowDout_3__0__3), .A2 (
         WindowWR), .B0 (WindowDout_2__0__3), .B1 (nx8178)) ;
    dff L0_2_L1_0_Wij_reg_Dout_4 (.Q (WindowDout_2__0__4), .QB (\$dummy [92]), .D (
        nx4261), .CLK (CLK)) ;
    ao32 ix4262 (.Y (nx4261), .A0 (nx8080), .A1 (WindowDout_3__0__4), .A2 (
         WindowWR), .B0 (WindowDout_2__0__4), .B1 (nx8178)) ;
    dff L0_2_L1_0_Wij_reg_Dout_5 (.Q (WindowDout_2__0__5), .QB (\$dummy [93]), .D (
        nx4271), .CLK (CLK)) ;
    ao32 ix4272 (.Y (nx4271), .A0 (nx8080), .A1 (WindowDout_3__0__5), .A2 (
         WindowWR), .B0 (WindowDout_2__0__5), .B1 (nx8178)) ;
    dff L0_2_L1_0_Wij_reg_Dout_6 (.Q (WindowDout_2__0__6), .QB (\$dummy [94]), .D (
        nx4281), .CLK (CLK)) ;
    ao32 ix4282 (.Y (nx4281), .A0 (nx8080), .A1 (WindowDout_3__0__6), .A2 (
         WindowWR), .B0 (WindowDout_2__0__6), .B1 (nx8180)) ;
    dff L0_2_L1_0_Wij_reg_Dout_7 (.Q (WindowDout_2__0__7), .QB (\$dummy [95]), .D (
        nx4291), .CLK (CLK)) ;
    ao32 ix4292 (.Y (nx4291), .A0 (nx8080), .A1 (WindowDout_3__0__7), .A2 (
         WindowWR), .B0 (WindowDout_2__0__7), .B1 (nx8180)) ;
    oai21 ix4382 (.Y (nx4381), .A0 (nx6486), .A1 (nx7928), .B0 (nx6488)) ;
    dff L0_1_L1_4_Wij_reg_Dout_0 (.Q (WindowDout_1__4__0), .QB (nx6486), .D (
        nx4381), .CLK (CLK)) ;
    oai21 ix4392 (.Y (nx4391), .A0 (nx6492), .A1 (nx7928), .B0 (nx6494)) ;
    dff L0_1_L1_4_Wij_reg_Dout_1 (.Q (WindowDout_1__4__1), .QB (nx6492), .D (
        nx4391), .CLK (CLK)) ;
    oai21 ix4402 (.Y (nx4401), .A0 (nx6498), .A1 (nx7928), .B0 (nx6500)) ;
    dff L0_1_L1_4_Wij_reg_Dout_2 (.Q (WindowDout_1__4__2), .QB (nx6498), .D (
        nx4401), .CLK (CLK)) ;
    oai21 ix4412 (.Y (nx4411), .A0 (nx6504), .A1 (nx7930), .B0 (nx6506)) ;
    dff L0_1_L1_4_Wij_reg_Dout_3 (.Q (WindowDout_1__4__3), .QB (nx6504), .D (
        nx4411), .CLK (CLK)) ;
    oai21 ix4422 (.Y (nx4421), .A0 (nx6510), .A1 (nx7930), .B0 (nx6512)) ;
    dff L0_1_L1_4_Wij_reg_Dout_4 (.Q (WindowDout_1__4__4), .QB (nx6510), .D (
        nx4421), .CLK (CLK)) ;
    oai21 ix4432 (.Y (nx4431), .A0 (nx6516), .A1 (nx7930), .B0 (nx6518)) ;
    dff L0_1_L1_4_Wij_reg_Dout_5 (.Q (WindowDout_1__4__5), .QB (nx6516), .D (
        nx4431), .CLK (CLK)) ;
    oai21 ix4442 (.Y (nx4441), .A0 (nx6522), .A1 (nx7930), .B0 (nx6524)) ;
    dff L0_1_L1_4_Wij_reg_Dout_6 (.Q (WindowDout_1__4__6), .QB (nx6522), .D (
        nx4441), .CLK (CLK)) ;
    oai21 ix4452 (.Y (nx4451), .A0 (nx6528), .A1 (nx7932), .B0 (nx6530)) ;
    dff L0_1_L1_4_Wij_reg_Dout_7 (.Q (WindowDout_1__4__7), .QB (nx6528), .D (
        nx4451), .CLK (CLK)) ;
    oai21 ix4702 (.Y (nx4701), .A0 (nx6534), .A1 (nx7932), .B0 (nx6536)) ;
    dff L0_1_L1_3_Wij_reg_Dout_0 (.Q (WindowDout_1__3__0), .QB (nx6534), .D (
        nx4701), .CLK (CLK)) ;
    oai21 ix4712 (.Y (nx4711), .A0 (nx6540), .A1 (nx7932), .B0 (nx6542)) ;
    dff L0_1_L1_3_Wij_reg_Dout_1 (.Q (WindowDout_1__3__1), .QB (nx6540), .D (
        nx4711), .CLK (CLK)) ;
    oai21 ix4722 (.Y (nx4721), .A0 (nx6546), .A1 (nx7934), .B0 (nx6548)) ;
    dff L0_1_L1_3_Wij_reg_Dout_2 (.Q (WindowDout_1__3__2), .QB (nx6546), .D (
        nx4721), .CLK (CLK)) ;
    oai21 ix4732 (.Y (nx4731), .A0 (nx6552), .A1 (nx7934), .B0 (nx6554)) ;
    dff L0_1_L1_3_Wij_reg_Dout_3 (.Q (WindowDout_1__3__3), .QB (nx6552), .D (
        nx4731), .CLK (CLK)) ;
    oai21 ix4742 (.Y (nx4741), .A0 (nx6558), .A1 (nx7934), .B0 (nx6560)) ;
    dff L0_1_L1_3_Wij_reg_Dout_4 (.Q (WindowDout_1__3__4), .QB (nx6558), .D (
        nx4741), .CLK (CLK)) ;
    oai21 ix4752 (.Y (nx4751), .A0 (nx6564), .A1 (nx7934), .B0 (nx6566)) ;
    dff L0_1_L1_3_Wij_reg_Dout_5 (.Q (WindowDout_1__3__5), .QB (nx6564), .D (
        nx4751), .CLK (CLK)) ;
    oai21 ix4762 (.Y (nx4761), .A0 (nx6570), .A1 (nx7936), .B0 (nx6572)) ;
    dff L0_1_L1_3_Wij_reg_Dout_6 (.Q (WindowDout_1__3__6), .QB (nx6570), .D (
        nx4761), .CLK (CLK)) ;
    oai21 ix4772 (.Y (nx4771), .A0 (nx6576), .A1 (nx7936), .B0 (nx6578)) ;
    dff L0_1_L1_3_Wij_reg_Dout_7 (.Q (WindowDout_1__3__7), .QB (nx6576), .D (
        nx4771), .CLK (CLK)) ;
    oai21 ix5022 (.Y (nx5021), .A0 (nx6582), .A1 (nx7936), .B0 (nx6584)) ;
    dff L0_1_L1_2_Wij_reg_Dout_0 (.Q (WindowDout_1__2__0), .QB (nx6582), .D (
        nx5021), .CLK (CLK)) ;
    nand03 ix6585 (.Y (nx6584), .A0 (nx8086), .A1 (WindowDout_2__2__0), .A2 (
           nx7936)) ;
    oai21 ix5032 (.Y (nx5031), .A0 (nx6588), .A1 (nx7938), .B0 (nx6590)) ;
    dff L0_1_L1_2_Wij_reg_Dout_1 (.Q (WindowDout_1__2__1), .QB (nx6588), .D (
        nx5031), .CLK (CLK)) ;
    nand03 ix6591 (.Y (nx6590), .A0 (nx8086), .A1 (WindowDout_2__2__1), .A2 (
           nx7938)) ;
    oai21 ix5042 (.Y (nx5041), .A0 (nx6594), .A1 (nx7938), .B0 (nx6596)) ;
    dff L0_1_L1_2_Wij_reg_Dout_2 (.Q (WindowDout_1__2__2), .QB (nx6594), .D (
        nx5041), .CLK (CLK)) ;
    nand03 ix6597 (.Y (nx6596), .A0 (nx8086), .A1 (WindowDout_2__2__2), .A2 (
           nx7938)) ;
    oai21 ix5052 (.Y (nx5051), .A0 (nx6600), .A1 (nx7938), .B0 (nx6602)) ;
    dff L0_1_L1_2_Wij_reg_Dout_3 (.Q (WindowDout_1__2__3), .QB (nx6600), .D (
        nx5051), .CLK (CLK)) ;
    nand03 ix6603 (.Y (nx6602), .A0 (nx8086), .A1 (WindowDout_2__2__3), .A2 (
           nx7938)) ;
    oai21 ix5062 (.Y (nx5061), .A0 (nx6606), .A1 (nx7938), .B0 (nx6608)) ;
    dff L0_1_L1_2_Wij_reg_Dout_4 (.Q (WindowDout_1__2__4), .QB (nx6606), .D (
        nx5061), .CLK (CLK)) ;
    nand03 ix6609 (.Y (nx6608), .A0 (nx8086), .A1 (WindowDout_2__2__4), .A2 (
           nx7940)) ;
    oai21 ix5072 (.Y (nx5071), .A0 (nx6612), .A1 (nx7940), .B0 (nx6614)) ;
    dff L0_1_L1_2_Wij_reg_Dout_5 (.Q (WindowDout_1__2__5), .QB (nx6612), .D (
        nx5071), .CLK (CLK)) ;
    nand03 ix6615 (.Y (nx6614), .A0 (nx8086), .A1 (WindowDout_2__2__5), .A2 (
           nx7940)) ;
    oai21 ix5082 (.Y (nx5081), .A0 (nx6618), .A1 (nx7940), .B0 (nx6620)) ;
    dff L0_1_L1_2_Wij_reg_Dout_6 (.Q (WindowDout_1__2__6), .QB (nx6618), .D (
        nx5081), .CLK (CLK)) ;
    nand03 ix6621 (.Y (nx6620), .A0 (nx8088), .A1 (WindowDout_2__2__6), .A2 (
           nx7940)) ;
    oai21 ix5092 (.Y (nx5091), .A0 (nx6624), .A1 (nx7940), .B0 (nx6626)) ;
    dff L0_1_L1_2_Wij_reg_Dout_7 (.Q (WindowDout_1__2__7), .QB (nx6624), .D (
        nx5091), .CLK (CLK)) ;
    nand03 ix6627 (.Y (nx6626), .A0 (nx8088), .A1 (WindowDout_2__2__7), .A2 (
           nx7940)) ;
    oai21 ix5342 (.Y (nx5341), .A0 (nx6630), .A1 (nx7942), .B0 (nx6632)) ;
    dff L0_1_L1_1_Wij_reg_Dout_0 (.Q (WindowDout_1__1__0), .QB (nx6630), .D (
        nx5341), .CLK (CLK)) ;
    nand03 ix6633 (.Y (nx6632), .A0 (nx8088), .A1 (WindowDout_2__1__0), .A2 (
           nx7942)) ;
    oai21 ix5352 (.Y (nx5351), .A0 (nx6636), .A1 (nx7942), .B0 (nx6638)) ;
    dff L0_1_L1_1_Wij_reg_Dout_1 (.Q (WindowDout_1__1__1), .QB (nx6636), .D (
        nx5351), .CLK (CLK)) ;
    nand03 ix6639 (.Y (nx6638), .A0 (nx8088), .A1 (WindowDout_2__1__1), .A2 (
           nx7942)) ;
    oai21 ix5362 (.Y (nx5361), .A0 (nx6642), .A1 (nx7942), .B0 (nx6644)) ;
    dff L0_1_L1_1_Wij_reg_Dout_2 (.Q (WindowDout_1__1__2), .QB (nx6642), .D (
        nx5361), .CLK (CLK)) ;
    nand03 ix6645 (.Y (nx6644), .A0 (nx8088), .A1 (WindowDout_2__1__2), .A2 (
           nx7942)) ;
    oai21 ix5372 (.Y (nx5371), .A0 (nx6648), .A1 (nx7942), .B0 (nx6650)) ;
    dff L0_1_L1_1_Wij_reg_Dout_3 (.Q (WindowDout_1__1__3), .QB (nx6648), .D (
        nx5371), .CLK (CLK)) ;
    nand03 ix6651 (.Y (nx6650), .A0 (nx8088), .A1 (WindowDout_2__1__3), .A2 (
           nx7944)) ;
    oai21 ix5382 (.Y (nx5381), .A0 (nx6654), .A1 (nx7944), .B0 (nx6656)) ;
    dff L0_1_L1_1_Wij_reg_Dout_4 (.Q (WindowDout_1__1__4), .QB (nx6654), .D (
        nx5381), .CLK (CLK)) ;
    nand03 ix6657 (.Y (nx6656), .A0 (nx8088), .A1 (WindowDout_2__1__4), .A2 (
           nx7944)) ;
    oai21 ix5392 (.Y (nx5391), .A0 (nx6660), .A1 (nx7944), .B0 (nx6662)) ;
    dff L0_1_L1_1_Wij_reg_Dout_5 (.Q (WindowDout_1__1__5), .QB (nx6660), .D (
        nx5391), .CLK (CLK)) ;
    nand03 ix6663 (.Y (nx6662), .A0 (nx8090), .A1 (WindowDout_2__1__5), .A2 (
           nx7944)) ;
    oai21 ix5402 (.Y (nx5401), .A0 (nx6666), .A1 (nx7944), .B0 (nx6668)) ;
    dff L0_1_L1_1_Wij_reg_Dout_6 (.Q (WindowDout_1__1__6), .QB (nx6666), .D (
        nx5401), .CLK (CLK)) ;
    nand03 ix6669 (.Y (nx6668), .A0 (nx8090), .A1 (WindowDout_2__1__6), .A2 (
           nx7944)) ;
    oai21 ix5412 (.Y (nx5411), .A0 (nx6672), .A1 (nx7946), .B0 (nx6674)) ;
    dff L0_1_L1_1_Wij_reg_Dout_7 (.Q (WindowDout_1__1__7), .QB (nx6672), .D (
        nx5411), .CLK (CLK)) ;
    nand03 ix6675 (.Y (nx6674), .A0 (nx8090), .A1 (WindowDout_2__1__7), .A2 (
           nx7946)) ;
    oai21 ix5662 (.Y (nx5661), .A0 (nx6678), .A1 (nx7946), .B0 (nx6680)) ;
    dff L0_1_L1_0_Wij_reg_Dout_0 (.Q (WindowDout_1__0__0), .QB (nx6678), .D (
        nx5661), .CLK (CLK)) ;
    nand03 ix6681 (.Y (nx6680), .A0 (nx8090), .A1 (WindowDout_2__0__0), .A2 (
           nx7946)) ;
    oai21 ix5672 (.Y (nx5671), .A0 (nx6684), .A1 (nx7946), .B0 (nx6686)) ;
    dff L0_1_L1_0_Wij_reg_Dout_1 (.Q (WindowDout_1__0__1), .QB (nx6684), .D (
        nx5671), .CLK (CLK)) ;
    nand03 ix6687 (.Y (nx6686), .A0 (nx8090), .A1 (WindowDout_2__0__1), .A2 (
           nx7946)) ;
    oai21 ix5682 (.Y (nx5681), .A0 (nx6690), .A1 (nx7946), .B0 (nx6692)) ;
    dff L0_1_L1_0_Wij_reg_Dout_2 (.Q (WindowDout_1__0__2), .QB (nx6690), .D (
        nx5681), .CLK (CLK)) ;
    nand03 ix6693 (.Y (nx6692), .A0 (nx8090), .A1 (WindowDout_2__0__2), .A2 (
           nx7948)) ;
    oai21 ix5692 (.Y (nx5691), .A0 (nx6696), .A1 (nx7948), .B0 (nx6698)) ;
    dff L0_1_L1_0_Wij_reg_Dout_3 (.Q (WindowDout_1__0__3), .QB (nx6696), .D (
        nx5691), .CLK (CLK)) ;
    nand03 ix6699 (.Y (nx6698), .A0 (nx8090), .A1 (WindowDout_2__0__3), .A2 (
           nx7948)) ;
    oai21 ix5702 (.Y (nx5701), .A0 (nx6702), .A1 (nx7948), .B0 (nx6704)) ;
    dff L0_1_L1_0_Wij_reg_Dout_4 (.Q (WindowDout_1__0__4), .QB (nx6702), .D (
        nx5701), .CLK (CLK)) ;
    nand03 ix6705 (.Y (nx6704), .A0 (nx8092), .A1 (WindowDout_2__0__4), .A2 (
           nx7948)) ;
    oai21 ix5712 (.Y (nx5711), .A0 (nx6708), .A1 (nx7948), .B0 (nx6710)) ;
    dff L0_1_L1_0_Wij_reg_Dout_5 (.Q (WindowDout_1__0__5), .QB (nx6708), .D (
        nx5711), .CLK (CLK)) ;
    nand03 ix6711 (.Y (nx6710), .A0 (nx8092), .A1 (WindowDout_2__0__5), .A2 (
           nx7948)) ;
    oai21 ix5722 (.Y (nx5721), .A0 (nx6714), .A1 (nx7950), .B0 (nx6716)) ;
    dff L0_1_L1_0_Wij_reg_Dout_6 (.Q (WindowDout_1__0__6), .QB (nx6714), .D (
        nx5721), .CLK (CLK)) ;
    nand03 ix6717 (.Y (nx6716), .A0 (nx8092), .A1 (WindowDout_2__0__6), .A2 (
           nx7950)) ;
    oai21 ix5732 (.Y (nx5731), .A0 (nx6720), .A1 (nx7950), .B0 (nx6722)) ;
    dff L0_1_L1_0_Wij_reg_Dout_7 (.Q (WindowDout_1__0__7), .QB (nx6720), .D (
        nx5731), .CLK (CLK)) ;
    nand03 ix6723 (.Y (nx6722), .A0 (nx8092), .A1 (WindowDout_2__0__7), .A2 (
           nx7950)) ;
    oai21 ix4462 (.Y (nx4461), .A0 (nx6726), .A1 (nx7950), .B0 (nx6728)) ;
    dff L0_0_L1_4_Wij_reg_Dout_0 (.Q (WindowDout_0__4__0), .QB (nx6726), .D (
        nx4461), .CLK (CLK)) ;
    oai21 ix4472 (.Y (nx4471), .A0 (nx6732), .A1 (nx7950), .B0 (nx6734)) ;
    dff L0_0_L1_4_Wij_reg_Dout_1 (.Q (WindowDout_0__4__1), .QB (nx6732), .D (
        nx4471), .CLK (CLK)) ;
    oai21 ix4482 (.Y (nx4481), .A0 (nx6738), .A1 (nx7952), .B0 (nx6740)) ;
    dff L0_0_L1_4_Wij_reg_Dout_2 (.Q (WindowDout_0__4__2), .QB (nx6738), .D (
        nx4481), .CLK (CLK)) ;
    oai21 ix4492 (.Y (nx4491), .A0 (nx6744), .A1 (nx7952), .B0 (nx6746)) ;
    dff L0_0_L1_4_Wij_reg_Dout_3 (.Q (WindowDout_0__4__3), .QB (nx6744), .D (
        nx4491), .CLK (CLK)) ;
    oai21 ix4502 (.Y (nx4501), .A0 (nx6750), .A1 (nx7952), .B0 (nx6752)) ;
    dff L0_0_L1_4_Wij_reg_Dout_4 (.Q (WindowDout_0__4__4), .QB (nx6750), .D (
        nx4501), .CLK (CLK)) ;
    oai21 ix4512 (.Y (nx4511), .A0 (nx6756), .A1 (nx7954), .B0 (nx6758)) ;
    dff L0_0_L1_4_Wij_reg_Dout_5 (.Q (WindowDout_0__4__5), .QB (nx6756), .D (
        nx4511), .CLK (CLK)) ;
    oai21 ix4522 (.Y (nx4521), .A0 (nx6762), .A1 (nx7954), .B0 (nx6764)) ;
    dff L0_0_L1_4_Wij_reg_Dout_6 (.Q (WindowDout_0__4__6), .QB (nx6762), .D (
        nx4521), .CLK (CLK)) ;
    oai21 ix4532 (.Y (nx4531), .A0 (nx6768), .A1 (nx7954), .B0 (nx6770)) ;
    dff L0_0_L1_4_Wij_reg_Dout_7 (.Q (WindowDout_0__4__7), .QB (nx6768), .D (
        nx4531), .CLK (CLK)) ;
    oai21 ix4782 (.Y (nx4781), .A0 (nx6774), .A1 (nx7954), .B0 (nx6776)) ;
    dff L0_0_L1_3_Wij_reg_Dout_0 (.Q (WindowDout_0__3__0), .QB (nx6774), .D (
        nx4781), .CLK (CLK)) ;
    oai21 ix4792 (.Y (nx4791), .A0 (nx6780), .A1 (nx7956), .B0 (nx6782)) ;
    dff L0_0_L1_3_Wij_reg_Dout_1 (.Q (WindowDout_0__3__1), .QB (nx6780), .D (
        nx4791), .CLK (CLK)) ;
    oai21 ix4802 (.Y (nx4801), .A0 (nx6786), .A1 (nx7956), .B0 (nx6788)) ;
    dff L0_0_L1_3_Wij_reg_Dout_2 (.Q (WindowDout_0__3__2), .QB (nx6786), .D (
        nx4801), .CLK (CLK)) ;
    oai21 ix4812 (.Y (nx4811), .A0 (nx6792), .A1 (nx7956), .B0 (nx6794)) ;
    dff L0_0_L1_3_Wij_reg_Dout_3 (.Q (WindowDout_0__3__3), .QB (nx6792), .D (
        nx4811), .CLK (CLK)) ;
    oai21 ix4822 (.Y (nx4821), .A0 (nx6798), .A1 (nx7958), .B0 (nx6800)) ;
    dff L0_0_L1_3_Wij_reg_Dout_4 (.Q (WindowDout_0__3__4), .QB (nx6798), .D (
        nx4821), .CLK (CLK)) ;
    oai21 ix4832 (.Y (nx4831), .A0 (nx6804), .A1 (nx7958), .B0 (nx6806)) ;
    dff L0_0_L1_3_Wij_reg_Dout_5 (.Q (WindowDout_0__3__5), .QB (nx6804), .D (
        nx4831), .CLK (CLK)) ;
    oai21 ix4842 (.Y (nx4841), .A0 (nx6810), .A1 (nx7958), .B0 (nx6812)) ;
    dff L0_0_L1_3_Wij_reg_Dout_6 (.Q (WindowDout_0__3__6), .QB (nx6810), .D (
        nx4841), .CLK (CLK)) ;
    oai21 ix4852 (.Y (nx4851), .A0 (nx6816), .A1 (nx7958), .B0 (nx6818)) ;
    dff L0_0_L1_3_Wij_reg_Dout_7 (.Q (WindowDout_0__3__7), .QB (nx6816), .D (
        nx4851), .CLK (CLK)) ;
    oai21 ix5102 (.Y (nx5101), .A0 (nx6822), .A1 (nx7960), .B0 (nx6824)) ;
    dff L0_0_L1_2_Wij_reg_Dout_0 (.Q (WindowDout_0__2__0), .QB (nx6822), .D (
        nx5101), .CLK (CLK)) ;
    oai21 ix5112 (.Y (nx5111), .A0 (nx6828), .A1 (nx7960), .B0 (nx6830)) ;
    dff L0_0_L1_2_Wij_reg_Dout_1 (.Q (WindowDout_0__2__1), .QB (nx6828), .D (
        nx5111), .CLK (CLK)) ;
    oai21 ix5122 (.Y (nx5121), .A0 (nx6834), .A1 (nx7960), .B0 (nx6836)) ;
    dff L0_0_L1_2_Wij_reg_Dout_2 (.Q (WindowDout_0__2__2), .QB (nx6834), .D (
        nx5121), .CLK (CLK)) ;
    oai21 ix5132 (.Y (nx5131), .A0 (nx6840), .A1 (nx7962), .B0 (nx6842)) ;
    dff L0_0_L1_2_Wij_reg_Dout_3 (.Q (WindowDout_0__2__3), .QB (nx6840), .D (
        nx5131), .CLK (CLK)) ;
    oai21 ix5142 (.Y (nx5141), .A0 (nx6846), .A1 (nx7962), .B0 (nx6848)) ;
    dff L0_0_L1_2_Wij_reg_Dout_4 (.Q (WindowDout_0__2__4), .QB (nx6846), .D (
        nx5141), .CLK (CLK)) ;
    oai21 ix5152 (.Y (nx5151), .A0 (nx6852), .A1 (nx7962), .B0 (nx6854)) ;
    dff L0_0_L1_2_Wij_reg_Dout_5 (.Q (WindowDout_0__2__5), .QB (nx6852), .D (
        nx5151), .CLK (CLK)) ;
    oai21 ix5162 (.Y (nx5161), .A0 (nx6858), .A1 (nx7962), .B0 (nx6860)) ;
    dff L0_0_L1_2_Wij_reg_Dout_6 (.Q (WindowDout_0__2__6), .QB (nx6858), .D (
        nx5161), .CLK (CLK)) ;
    oai21 ix5172 (.Y (nx5171), .A0 (nx6864), .A1 (nx7964), .B0 (nx6866)) ;
    dff L0_0_L1_2_Wij_reg_Dout_7 (.Q (WindowDout_0__2__7), .QB (nx6864), .D (
        nx5171), .CLK (CLK)) ;
    oai21 ix5422 (.Y (nx5421), .A0 (nx6870), .A1 (nx7964), .B0 (nx6872)) ;
    dff L0_0_L1_1_Wij_reg_Dout_0 (.Q (WindowDout_0__1__0), .QB (nx6870), .D (
        nx5421), .CLK (CLK)) ;
    oai21 ix5432 (.Y (nx5431), .A0 (nx6876), .A1 (nx7964), .B0 (nx6878)) ;
    dff L0_0_L1_1_Wij_reg_Dout_1 (.Q (WindowDout_0__1__1), .QB (nx6876), .D (
        nx5431), .CLK (CLK)) ;
    oai21 ix5442 (.Y (nx5441), .A0 (nx6882), .A1 (nx7966), .B0 (nx6884)) ;
    dff L0_0_L1_1_Wij_reg_Dout_2 (.Q (WindowDout_0__1__2), .QB (nx6882), .D (
        nx5441), .CLK (CLK)) ;
    oai21 ix5452 (.Y (nx5451), .A0 (nx6888), .A1 (nx7966), .B0 (nx6890)) ;
    dff L0_0_L1_1_Wij_reg_Dout_3 (.Q (WindowDout_0__1__3), .QB (nx6888), .D (
        nx5451), .CLK (CLK)) ;
    oai21 ix5462 (.Y (nx5461), .A0 (nx6894), .A1 (nx7966), .B0 (nx6896)) ;
    dff L0_0_L1_1_Wij_reg_Dout_4 (.Q (WindowDout_0__1__4), .QB (nx6894), .D (
        nx5461), .CLK (CLK)) ;
    oai21 ix5472 (.Y (nx5471), .A0 (nx6900), .A1 (nx7966), .B0 (nx6902)) ;
    dff L0_0_L1_1_Wij_reg_Dout_5 (.Q (WindowDout_0__1__5), .QB (nx6900), .D (
        nx5471), .CLK (CLK)) ;
    oai21 ix5482 (.Y (nx5481), .A0 (nx6906), .A1 (nx7968), .B0 (nx6908)) ;
    dff L0_0_L1_1_Wij_reg_Dout_6 (.Q (WindowDout_0__1__6), .QB (nx6906), .D (
        nx5481), .CLK (CLK)) ;
    oai21 ix5492 (.Y (nx5491), .A0 (nx6912), .A1 (nx7968), .B0 (nx6914)) ;
    dff L0_0_L1_1_Wij_reg_Dout_7 (.Q (WindowDout_0__1__7), .QB (nx6912), .D (
        nx5491), .CLK (CLK)) ;
    oai21 ix5742 (.Y (nx5741), .A0 (nx6918), .A1 (nx7968), .B0 (nx6920)) ;
    dff L0_0_L1_0_Wij_reg_Dout_0 (.Q (WindowDout_0__0__0), .QB (nx6918), .D (
        nx5741), .CLK (CLK)) ;
    oai21 ix5752 (.Y (nx5751), .A0 (nx6924), .A1 (nx7970), .B0 (nx6926)) ;
    dff L0_0_L1_0_Wij_reg_Dout_1 (.Q (WindowDout_0__0__1), .QB (nx6924), .D (
        nx5751), .CLK (CLK)) ;
    oai21 ix5762 (.Y (nx5761), .A0 (nx6930), .A1 (nx7970), .B0 (nx6932)) ;
    dff L0_0_L1_0_Wij_reg_Dout_2 (.Q (WindowDout_0__0__2), .QB (nx6930), .D (
        nx5761), .CLK (CLK)) ;
    oai21 ix5772 (.Y (nx5771), .A0 (nx6936), .A1 (nx7970), .B0 (nx6938)) ;
    dff L0_0_L1_0_Wij_reg_Dout_3 (.Q (WindowDout_0__0__3), .QB (nx6936), .D (
        nx5771), .CLK (CLK)) ;
    oai21 ix5782 (.Y (nx5781), .A0 (nx6942), .A1 (nx7970), .B0 (nx6944)) ;
    dff L0_0_L1_0_Wij_reg_Dout_4 (.Q (WindowDout_0__0__4), .QB (nx6942), .D (
        nx5781), .CLK (CLK)) ;
    oai21 ix5792 (.Y (nx5791), .A0 (nx6948), .A1 (nx7972), .B0 (nx6950)) ;
    dff L0_0_L1_0_Wij_reg_Dout_5 (.Q (WindowDout_0__0__5), .QB (nx6948), .D (
        nx5791), .CLK (CLK)) ;
    oai21 ix5802 (.Y (nx5801), .A0 (nx6954), .A1 (nx7972), .B0 (nx6956)) ;
    dff L0_0_L1_0_Wij_reg_Dout_6 (.Q (WindowDout_0__0__6), .QB (nx6954), .D (
        nx5801), .CLK (CLK)) ;
    oai21 ix5812 (.Y (nx5811), .A0 (nx6960), .A1 (nx7972), .B0 (nx6962)) ;
    dff L0_0_L1_0_Wij_reg_Dout_7 (.Q (WindowDout_0__0__7), .QB (nx6960), .D (
        nx5811), .CLK (CLK)) ;
    dff L0_4_L1_4_Fij_reg_Dout_0 (.Q (FilterDout_4__4__0), .QB (\$dummy [96]), .D (
        nx2061), .CLK (CLK)) ;
    aoi21 ix6967 (.Y (nx6966), .A0 (FilterSize), .A1 (FilterWR), .B0 (RST)) ;
    dff L0_4_L1_4_Fij_reg_Dout_1 (.Q (FilterDout_4__4__1), .QB (\$dummy [97]), .D (
        nx2071), .CLK (CLK)) ;
    dff L0_4_L1_4_Fij_reg_Dout_2 (.Q (FilterDout_4__4__2), .QB (\$dummy [98]), .D (
        nx2081), .CLK (CLK)) ;
    dff L0_4_L1_4_Fij_reg_Dout_3 (.Q (FilterDout_4__4__3), .QB (\$dummy [99]), .D (
        nx2091), .CLK (CLK)) ;
    dff L0_4_L1_4_Fij_reg_Dout_4 (.Q (FilterDout_4__4__4), .QB (\$dummy [100]), 
        .D (nx2101), .CLK (CLK)) ;
    dff L0_4_L1_4_Fij_reg_Dout_5 (.Q (FilterDout_4__4__5), .QB (\$dummy [101]), 
        .D (nx2111), .CLK (CLK)) ;
    dff L0_4_L1_4_Fij_reg_Dout_6 (.Q (FilterDout_4__4__6), .QB (\$dummy [102]), 
        .D (nx2121), .CLK (CLK)) ;
    dff L0_4_L1_4_Fij_reg_Dout_7 (.Q (FilterDout_4__4__7), .QB (\$dummy [103]), 
        .D (nx2131), .CLK (CLK)) ;
    dff L0_4_L1_3_Fij_reg_Dout_0 (.Q (FilterDout_4__3__0), .QB (\$dummy [104]), 
        .D (nx2221), .CLK (CLK)) ;
    dff L0_4_L1_3_Fij_reg_Dout_1 (.Q (FilterDout_4__3__1), .QB (\$dummy [105]), 
        .D (nx2231), .CLK (CLK)) ;
    dff L0_4_L1_3_Fij_reg_Dout_2 (.Q (FilterDout_4__3__2), .QB (\$dummy [106]), 
        .D (nx2241), .CLK (CLK)) ;
    dff L0_4_L1_3_Fij_reg_Dout_3 (.Q (FilterDout_4__3__3), .QB (\$dummy [107]), 
        .D (nx2251), .CLK (CLK)) ;
    dff L0_4_L1_3_Fij_reg_Dout_4 (.Q (FilterDout_4__3__4), .QB (\$dummy [108]), 
        .D (nx2261), .CLK (CLK)) ;
    dff L0_4_L1_3_Fij_reg_Dout_5 (.Q (FilterDout_4__3__5), .QB (\$dummy [109]), 
        .D (nx2271), .CLK (CLK)) ;
    dff L0_4_L1_3_Fij_reg_Dout_6 (.Q (FilterDout_4__3__6), .QB (\$dummy [110]), 
        .D (nx2281), .CLK (CLK)) ;
    dff L0_4_L1_3_Fij_reg_Dout_7 (.Q (FilterDout_4__3__7), .QB (\$dummy [111]), 
        .D (nx2291), .CLK (CLK)) ;
    dff L0_4_L1_2_Fij_reg_Dout_0 (.Q (FilterDout_4__2__0), .QB (\$dummy [112]), 
        .D (nx2381), .CLK (CLK)) ;
    ao32 ix2382 (.Y (nx2381), .A0 (Din[16]), .A1 (nx8104), .A2 (FilterWR), .B0 (
         FilterDout_4__2__0), .B1 (nx8198)) ;
    nor02_2x ix7017 (.Y (nx7016), .A0 (FilterWR), .A1 (RST)) ;
    dff L0_4_L1_2_Fij_reg_Dout_1 (.Q (FilterDout_4__2__1), .QB (\$dummy [113]), 
        .D (nx2391), .CLK (CLK)) ;
    ao32 ix2392 (.Y (nx2391), .A0 (Din[17]), .A1 (nx8104), .A2 (FilterWR), .B0 (
         FilterDout_4__2__1), .B1 (nx8198)) ;
    dff L0_4_L1_2_Fij_reg_Dout_2 (.Q (FilterDout_4__2__2), .QB (\$dummy [114]), 
        .D (nx2401), .CLK (CLK)) ;
    ao32 ix2402 (.Y (nx2401), .A0 (Din[18]), .A1 (nx8104), .A2 (FilterWR), .B0 (
         FilterDout_4__2__2), .B1 (nx8198)) ;
    dff L0_4_L1_2_Fij_reg_Dout_3 (.Q (FilterDout_4__2__3), .QB (\$dummy [115]), 
        .D (nx2411), .CLK (CLK)) ;
    ao32 ix2412 (.Y (nx2411), .A0 (Din[19]), .A1 (nx8104), .A2 (FilterWR), .B0 (
         FilterDout_4__2__3), .B1 (nx8198)) ;
    dff L0_4_L1_2_Fij_reg_Dout_4 (.Q (FilterDout_4__2__4), .QB (\$dummy [116]), 
        .D (nx2421), .CLK (CLK)) ;
    ao32 ix2422 (.Y (nx2421), .A0 (Din[20]), .A1 (nx8104), .A2 (FilterWR), .B0 (
         FilterDout_4__2__4), .B1 (nx8198)) ;
    dff L0_4_L1_2_Fij_reg_Dout_5 (.Q (FilterDout_4__2__5), .QB (\$dummy [117]), 
        .D (nx2431), .CLK (CLK)) ;
    ao32 ix2432 (.Y (nx2431), .A0 (Din[21]), .A1 (nx8106), .A2 (FilterWR), .B0 (
         FilterDout_4__2__5), .B1 (nx8198)) ;
    dff L0_4_L1_2_Fij_reg_Dout_6 (.Q (FilterDout_4__2__6), .QB (\$dummy [118]), 
        .D (nx2441), .CLK (CLK)) ;
    ao32 ix2442 (.Y (nx2441), .A0 (Din[22]), .A1 (nx8106), .A2 (FilterWR), .B0 (
         FilterDout_4__2__6), .B1 (nx8198)) ;
    dff L0_4_L1_2_Fij_reg_Dout_7 (.Q (FilterDout_4__2__7), .QB (\$dummy [119]), 
        .D (nx2451), .CLK (CLK)) ;
    ao32 ix2452 (.Y (nx2451), .A0 (Din[23]), .A1 (nx8106), .A2 (FilterWR), .B0 (
         FilterDout_4__2__7), .B1 (nx8200)) ;
    dff L0_4_L1_1_Fij_reg_Dout_0 (.Q (FilterDout_4__1__0), .QB (\$dummy [120]), 
        .D (nx2541), .CLK (CLK)) ;
    ao32 ix2542 (.Y (nx2541), .A0 (Din[8]), .A1 (nx8106), .A2 (FilterWR), .B0 (
         FilterDout_4__1__0), .B1 (nx8200)) ;
    dff L0_4_L1_1_Fij_reg_Dout_1 (.Q (FilterDout_4__1__1), .QB (\$dummy [121]), 
        .D (nx2551), .CLK (CLK)) ;
    ao32 ix2552 (.Y (nx2551), .A0 (Din[9]), .A1 (nx8106), .A2 (FilterWR), .B0 (
         FilterDout_4__1__1), .B1 (nx8200)) ;
    dff L0_4_L1_1_Fij_reg_Dout_2 (.Q (FilterDout_4__1__2), .QB (\$dummy [122]), 
        .D (nx2561), .CLK (CLK)) ;
    ao32 ix2562 (.Y (nx2561), .A0 (Din[10]), .A1 (nx8106), .A2 (FilterWR), .B0 (
         FilterDout_4__1__2), .B1 (nx8200)) ;
    dff L0_4_L1_1_Fij_reg_Dout_3 (.Q (FilterDout_4__1__3), .QB (\$dummy [123]), 
        .D (nx2571), .CLK (CLK)) ;
    ao32 ix2572 (.Y (nx2571), .A0 (Din[11]), .A1 (nx8106), .A2 (FilterWR), .B0 (
         FilterDout_4__1__3), .B1 (nx8200)) ;
    dff L0_4_L1_1_Fij_reg_Dout_4 (.Q (FilterDout_4__1__4), .QB (\$dummy [124]), 
        .D (nx2581), .CLK (CLK)) ;
    ao32 ix2582 (.Y (nx2581), .A0 (Din[12]), .A1 (nx8108), .A2 (FilterWR), .B0 (
         FilterDout_4__1__4), .B1 (nx8200)) ;
    dff L0_4_L1_1_Fij_reg_Dout_5 (.Q (FilterDout_4__1__5), .QB (\$dummy [125]), 
        .D (nx2591), .CLK (CLK)) ;
    ao32 ix2592 (.Y (nx2591), .A0 (Din[13]), .A1 (nx8108), .A2 (FilterWR), .B0 (
         FilterDout_4__1__5), .B1 (nx8200)) ;
    dff L0_4_L1_1_Fij_reg_Dout_6 (.Q (FilterDout_4__1__6), .QB (\$dummy [126]), 
        .D (nx2601), .CLK (CLK)) ;
    ao32 ix2602 (.Y (nx2601), .A0 (Din[14]), .A1 (nx8108), .A2 (FilterWR), .B0 (
         FilterDout_4__1__6), .B1 (nx8202)) ;
    dff L0_4_L1_1_Fij_reg_Dout_7 (.Q (FilterDout_4__1__7), .QB (\$dummy [127]), 
        .D (nx2611), .CLK (CLK)) ;
    ao32 ix2612 (.Y (nx2611), .A0 (Din[15]), .A1 (nx8108), .A2 (FilterWR), .B0 (
         FilterDout_4__1__7), .B1 (nx8202)) ;
    dff L0_4_L1_0_Fij_reg_Dout_0 (.Q (FilterDout_4__0__0), .QB (\$dummy [128]), 
        .D (nx2701), .CLK (CLK)) ;
    ao32 ix2702 (.Y (nx2701), .A0 (Din[0]), .A1 (nx8108), .A2 (FilterWR), .B0 (
         FilterDout_4__0__0), .B1 (nx8202)) ;
    dff L0_4_L1_0_Fij_reg_Dout_1 (.Q (FilterDout_4__0__1), .QB (\$dummy [129]), 
        .D (nx2711), .CLK (CLK)) ;
    ao32 ix2712 (.Y (nx2711), .A0 (Din[1]), .A1 (nx8108), .A2 (FilterWR), .B0 (
         FilterDout_4__0__1), .B1 (nx8202)) ;
    dff L0_4_L1_0_Fij_reg_Dout_2 (.Q (FilterDout_4__0__2), .QB (\$dummy [130]), 
        .D (nx2721), .CLK (CLK)) ;
    ao32 ix2722 (.Y (nx2721), .A0 (Din[2]), .A1 (nx8108), .A2 (FilterWR), .B0 (
         FilterDout_4__0__2), .B1 (nx8202)) ;
    dff L0_4_L1_0_Fij_reg_Dout_3 (.Q (FilterDout_4__0__3), .QB (\$dummy [131]), 
        .D (nx2731), .CLK (CLK)) ;
    ao32 ix2732 (.Y (nx2731), .A0 (Din[3]), .A1 (nx8110), .A2 (FilterWR), .B0 (
         FilterDout_4__0__3), .B1 (nx8202)) ;
    dff L0_4_L1_0_Fij_reg_Dout_4 (.Q (FilterDout_4__0__4), .QB (\$dummy [132]), 
        .D (nx2741), .CLK (CLK)) ;
    ao32 ix2742 (.Y (nx2741), .A0 (Din[4]), .A1 (nx8110), .A2 (FilterWR), .B0 (
         FilterDout_4__0__4), .B1 (nx8202)) ;
    dff L0_4_L1_0_Fij_reg_Dout_5 (.Q (FilterDout_4__0__5), .QB (\$dummy [133]), 
        .D (nx2751), .CLK (CLK)) ;
    ao32 ix2752 (.Y (nx2751), .A0 (Din[5]), .A1 (nx8110), .A2 (FilterWR), .B0 (
         FilterDout_4__0__5), .B1 (nx8204)) ;
    dff L0_4_L1_0_Fij_reg_Dout_6 (.Q (FilterDout_4__0__6), .QB (\$dummy [134]), 
        .D (nx2761), .CLK (CLK)) ;
    ao32 ix2762 (.Y (nx2761), .A0 (Din[6]), .A1 (nx8110), .A2 (FilterWR), .B0 (
         FilterDout_4__0__6), .B1 (nx8204)) ;
    dff L0_4_L1_0_Fij_reg_Dout_7 (.Q (FilterDout_4__0__7), .QB (\$dummy [135]), 
        .D (nx2771), .CLK (CLK)) ;
    ao32 ix2772 (.Y (nx2771), .A0 (Din[7]), .A1 (nx8110), .A2 (FilterWR), .B0 (
         FilterDout_4__0__7), .B1 (nx8204)) ;
    oai21 ix2862 (.Y (nx2861), .A0 (nx7090), .A1 (nx7974), .B0 (nx7093)) ;
    dff L0_3_L1_4_Fij_reg_Dout_0 (.Q (FilterDout_3__4__0), .QB (nx7090), .D (
        nx2861), .CLK (CLK)) ;
    nand03 ix7094 (.Y (nx7093), .A0 (nx8110), .A1 (FilterDout_4__4__0), .A2 (
           nx7974)) ;
    oai21 ix2872 (.Y (nx2871), .A0 (nx7097), .A1 (nx7974), .B0 (nx7099)) ;
    dff L0_3_L1_4_Fij_reg_Dout_1 (.Q (FilterDout_3__4__1), .QB (nx7097), .D (
        nx2871), .CLK (CLK)) ;
    nand03 ix7100 (.Y (nx7099), .A0 (nx8110), .A1 (FilterDout_4__4__1), .A2 (
           nx7974)) ;
    oai21 ix2882 (.Y (nx2881), .A0 (nx7103), .A1 (nx7974), .B0 (nx7105)) ;
    dff L0_3_L1_4_Fij_reg_Dout_2 (.Q (FilterDout_3__4__2), .QB (nx7103), .D (
        nx2881), .CLK (CLK)) ;
    nand03 ix7106 (.Y (nx7105), .A0 (nx8112), .A1 (FilterDout_4__4__2), .A2 (
           nx7974)) ;
    oai21 ix2892 (.Y (nx2891), .A0 (nx7109), .A1 (nx7974), .B0 (nx7111)) ;
    dff L0_3_L1_4_Fij_reg_Dout_3 (.Q (FilterDout_3__4__3), .QB (nx7109), .D (
        nx2891), .CLK (CLK)) ;
    nand03 ix7112 (.Y (nx7111), .A0 (nx8112), .A1 (FilterDout_4__4__3), .A2 (
           nx7976)) ;
    oai21 ix2902 (.Y (nx2901), .A0 (nx7115), .A1 (nx7976), .B0 (nx7117)) ;
    dff L0_3_L1_4_Fij_reg_Dout_4 (.Q (FilterDout_3__4__4), .QB (nx7115), .D (
        nx2901), .CLK (CLK)) ;
    nand03 ix7118 (.Y (nx7117), .A0 (nx8112), .A1 (FilterDout_4__4__4), .A2 (
           nx7976)) ;
    oai21 ix2912 (.Y (nx2911), .A0 (nx7121), .A1 (nx7976), .B0 (nx7123)) ;
    dff L0_3_L1_4_Fij_reg_Dout_5 (.Q (FilterDout_3__4__5), .QB (nx7121), .D (
        nx2911), .CLK (CLK)) ;
    nand03 ix7124 (.Y (nx7123), .A0 (nx8112), .A1 (FilterDout_4__4__5), .A2 (
           nx7976)) ;
    oai21 ix2922 (.Y (nx2921), .A0 (nx7127), .A1 (nx7976), .B0 (nx7129)) ;
    dff L0_3_L1_4_Fij_reg_Dout_6 (.Q (FilterDout_3__4__6), .QB (nx7127), .D (
        nx2921), .CLK (CLK)) ;
    nand03 ix7130 (.Y (nx7129), .A0 (nx8112), .A1 (FilterDout_4__4__6), .A2 (
           nx7976)) ;
    oai21 ix2932 (.Y (nx2931), .A0 (nx7133), .A1 (nx7978), .B0 (nx7135)) ;
    dff L0_3_L1_4_Fij_reg_Dout_7 (.Q (FilterDout_3__4__7), .QB (nx7133), .D (
        nx2931), .CLK (CLK)) ;
    nand03 ix7136 (.Y (nx7135), .A0 (nx8112), .A1 (FilterDout_4__4__7), .A2 (
           nx7978)) ;
    oai21 ix3022 (.Y (nx3021), .A0 (nx7139), .A1 (nx7978), .B0 (nx7141)) ;
    dff L0_3_L1_3_Fij_reg_Dout_0 (.Q (FilterDout_3__3__0), .QB (nx7139), .D (
        nx3021), .CLK (CLK)) ;
    nand03 ix7142 (.Y (nx7141), .A0 (nx8112), .A1 (FilterDout_4__3__0), .A2 (
           nx7978)) ;
    oai21 ix3032 (.Y (nx3031), .A0 (nx7145), .A1 (nx7978), .B0 (nx7147)) ;
    dff L0_3_L1_3_Fij_reg_Dout_1 (.Q (FilterDout_3__3__1), .QB (nx7145), .D (
        nx3031), .CLK (CLK)) ;
    nand03 ix7148 (.Y (nx7147), .A0 (nx8114), .A1 (FilterDout_4__3__1), .A2 (
           nx7978)) ;
    oai21 ix3042 (.Y (nx3041), .A0 (nx7151), .A1 (nx7978), .B0 (nx7153)) ;
    dff L0_3_L1_3_Fij_reg_Dout_2 (.Q (FilterDout_3__3__2), .QB (nx7151), .D (
        nx3041), .CLK (CLK)) ;
    nand03 ix7154 (.Y (nx7153), .A0 (nx8114), .A1 (FilterDout_4__3__2), .A2 (
           nx7980)) ;
    oai21 ix3052 (.Y (nx3051), .A0 (nx7157), .A1 (nx7980), .B0 (nx7159)) ;
    dff L0_3_L1_3_Fij_reg_Dout_3 (.Q (FilterDout_3__3__3), .QB (nx7157), .D (
        nx3051), .CLK (CLK)) ;
    nand03 ix7160 (.Y (nx7159), .A0 (nx8114), .A1 (FilterDout_4__3__3), .A2 (
           nx7980)) ;
    oai21 ix3062 (.Y (nx3061), .A0 (nx7163), .A1 (nx7980), .B0 (nx7165)) ;
    dff L0_3_L1_3_Fij_reg_Dout_4 (.Q (FilterDout_3__3__4), .QB (nx7163), .D (
        nx3061), .CLK (CLK)) ;
    nand03 ix7166 (.Y (nx7165), .A0 (nx8114), .A1 (FilterDout_4__3__4), .A2 (
           nx7980)) ;
    oai21 ix3072 (.Y (nx3071), .A0 (nx7169), .A1 (nx7980), .B0 (nx7171)) ;
    dff L0_3_L1_3_Fij_reg_Dout_5 (.Q (FilterDout_3__3__5), .QB (nx7169), .D (
        nx3071), .CLK (CLK)) ;
    nand03 ix7172 (.Y (nx7171), .A0 (nx8114), .A1 (FilterDout_4__3__5), .A2 (
           nx7980)) ;
    oai21 ix3082 (.Y (nx3081), .A0 (nx7175), .A1 (nx7982), .B0 (nx7177)) ;
    dff L0_3_L1_3_Fij_reg_Dout_6 (.Q (FilterDout_3__3__6), .QB (nx7175), .D (
        nx3081), .CLK (CLK)) ;
    nand03 ix7178 (.Y (nx7177), .A0 (nx8114), .A1 (FilterDout_4__3__6), .A2 (
           nx7982)) ;
    oai21 ix3092 (.Y (nx3091), .A0 (nx7181), .A1 (nx7982), .B0 (nx7183)) ;
    dff L0_3_L1_3_Fij_reg_Dout_7 (.Q (FilterDout_3__3__7), .QB (nx7181), .D (
        nx3091), .CLK (CLK)) ;
    nand03 ix7184 (.Y (nx7183), .A0 (nx8114), .A1 (FilterDout_4__3__7), .A2 (
           nx7982)) ;
    dff L0_3_L1_2_Fij_reg_Dout_0 (.Q (FilterDout_3__2__0), .QB (\$dummy [136]), 
        .D (nx3181), .CLK (CLK)) ;
    ao32 ix3182 (.Y (nx3181), .A0 (nx8116), .A1 (FilterDout_4__2__0), .A2 (
         FilterWR), .B0 (FilterDout_3__2__0), .B1 (nx8204)) ;
    dff L0_3_L1_2_Fij_reg_Dout_1 (.Q (FilterDout_3__2__1), .QB (\$dummy [137]), 
        .D (nx3191), .CLK (CLK)) ;
    ao32 ix3192 (.Y (nx3191), .A0 (nx8116), .A1 (FilterDout_4__2__1), .A2 (
         FilterWR), .B0 (FilterDout_3__2__1), .B1 (nx8204)) ;
    dff L0_3_L1_2_Fij_reg_Dout_2 (.Q (FilterDout_3__2__2), .QB (\$dummy [138]), 
        .D (nx3201), .CLK (CLK)) ;
    ao32 ix3202 (.Y (nx3201), .A0 (nx8116), .A1 (FilterDout_4__2__2), .A2 (
         FilterWR), .B0 (FilterDout_3__2__2), .B1 (nx8204)) ;
    dff L0_3_L1_2_Fij_reg_Dout_3 (.Q (FilterDout_3__2__3), .QB (\$dummy [139]), 
        .D (nx3211), .CLK (CLK)) ;
    ao32 ix3212 (.Y (nx3211), .A0 (nx8116), .A1 (FilterDout_4__2__3), .A2 (
         FilterWR), .B0 (FilterDout_3__2__3), .B1 (nx8204)) ;
    dff L0_3_L1_2_Fij_reg_Dout_4 (.Q (FilterDout_3__2__4), .QB (\$dummy [140]), 
        .D (nx3221), .CLK (CLK)) ;
    ao32 ix3222 (.Y (nx3221), .A0 (nx8116), .A1 (FilterDout_4__2__4), .A2 (
         FilterWR), .B0 (FilterDout_3__2__4), .B1 (nx8206)) ;
    dff L0_3_L1_2_Fij_reg_Dout_5 (.Q (FilterDout_3__2__5), .QB (\$dummy [141]), 
        .D (nx3231), .CLK (CLK)) ;
    ao32 ix3232 (.Y (nx3231), .A0 (nx8116), .A1 (FilterDout_4__2__5), .A2 (
         FilterWR), .B0 (FilterDout_3__2__5), .B1 (nx8206)) ;
    dff L0_3_L1_2_Fij_reg_Dout_6 (.Q (FilterDout_3__2__6), .QB (\$dummy [142]), 
        .D (nx3241), .CLK (CLK)) ;
    ao32 ix3242 (.Y (nx3241), .A0 (nx8116), .A1 (FilterDout_4__2__6), .A2 (
         FilterWR), .B0 (FilterDout_3__2__6), .B1 (nx8206)) ;
    dff L0_3_L1_2_Fij_reg_Dout_7 (.Q (FilterDout_3__2__7), .QB (\$dummy [143]), 
        .D (nx3251), .CLK (CLK)) ;
    ao32 ix3252 (.Y (nx3251), .A0 (nx8118), .A1 (FilterDout_4__2__7), .A2 (
         FilterWR), .B0 (FilterDout_3__2__7), .B1 (nx8206)) ;
    dff L0_3_L1_1_Fij_reg_Dout_0 (.Q (FilterDout_3__1__0), .QB (\$dummy [144]), 
        .D (nx3341), .CLK (CLK)) ;
    ao32 ix3342 (.Y (nx3341), .A0 (nx8118), .A1 (FilterDout_4__1__0), .A2 (
         FilterWR), .B0 (FilterDout_3__1__0), .B1 (nx8206)) ;
    dff L0_3_L1_1_Fij_reg_Dout_1 (.Q (FilterDout_3__1__1), .QB (\$dummy [145]), 
        .D (nx3351), .CLK (CLK)) ;
    ao32 ix3352 (.Y (nx3351), .A0 (nx8118), .A1 (FilterDout_4__1__1), .A2 (
         FilterWR), .B0 (FilterDout_3__1__1), .B1 (nx8206)) ;
    dff L0_3_L1_1_Fij_reg_Dout_2 (.Q (FilterDout_3__1__2), .QB (\$dummy [146]), 
        .D (nx3361), .CLK (CLK)) ;
    ao32 ix3362 (.Y (nx3361), .A0 (nx8118), .A1 (FilterDout_4__1__2), .A2 (
         FilterWR), .B0 (FilterDout_3__1__2), .B1 (nx8206)) ;
    dff L0_3_L1_1_Fij_reg_Dout_3 (.Q (FilterDout_3__1__3), .QB (\$dummy [147]), 
        .D (nx3371), .CLK (CLK)) ;
    ao32 ix3372 (.Y (nx3371), .A0 (nx8118), .A1 (FilterDout_4__1__3), .A2 (
         FilterWR), .B0 (FilterDout_3__1__3), .B1 (nx8208)) ;
    dff L0_3_L1_1_Fij_reg_Dout_4 (.Q (FilterDout_3__1__4), .QB (\$dummy [148]), 
        .D (nx3381), .CLK (CLK)) ;
    ao32 ix3382 (.Y (nx3381), .A0 (nx8118), .A1 (FilterDout_4__1__4), .A2 (
         FilterWR), .B0 (FilterDout_3__1__4), .B1 (nx8208)) ;
    dff L0_3_L1_1_Fij_reg_Dout_5 (.Q (FilterDout_3__1__5), .QB (\$dummy [149]), 
        .D (nx3391), .CLK (CLK)) ;
    ao32 ix3392 (.Y (nx3391), .A0 (nx8118), .A1 (FilterDout_4__1__5), .A2 (
         FilterWR), .B0 (FilterDout_3__1__5), .B1 (nx8208)) ;
    dff L0_3_L1_1_Fij_reg_Dout_6 (.Q (FilterDout_3__1__6), .QB (\$dummy [150]), 
        .D (nx3401), .CLK (CLK)) ;
    ao32 ix3402 (.Y (nx3401), .A0 (nx8120), .A1 (FilterDout_4__1__6), .A2 (
         FilterWR), .B0 (FilterDout_3__1__6), .B1 (nx8208)) ;
    dff L0_3_L1_1_Fij_reg_Dout_7 (.Q (FilterDout_3__1__7), .QB (\$dummy [151]), 
        .D (nx3411), .CLK (CLK)) ;
    ao32 ix3412 (.Y (nx3411), .A0 (nx8120), .A1 (FilterDout_4__1__7), .A2 (
         FilterWR), .B0 (FilterDout_3__1__7), .B1 (nx8208)) ;
    dff L0_3_L1_0_Fij_reg_Dout_0 (.Q (FilterDout_3__0__0), .QB (\$dummy [152]), 
        .D (nx3501), .CLK (CLK)) ;
    ao32 ix3502 (.Y (nx3501), .A0 (nx8120), .A1 (FilterDout_4__0__0), .A2 (
         FilterWR), .B0 (FilterDout_3__0__0), .B1 (nx8208)) ;
    dff L0_3_L1_0_Fij_reg_Dout_1 (.Q (FilterDout_3__0__1), .QB (\$dummy [153]), 
        .D (nx3511), .CLK (CLK)) ;
    ao32 ix3512 (.Y (nx3511), .A0 (nx8120), .A1 (FilterDout_4__0__1), .A2 (
         FilterWR), .B0 (FilterDout_3__0__1), .B1 (nx8208)) ;
    dff L0_3_L1_0_Fij_reg_Dout_2 (.Q (FilterDout_3__0__2), .QB (\$dummy [154]), 
        .D (nx3521), .CLK (CLK)) ;
    ao32 ix3522 (.Y (nx3521), .A0 (nx8120), .A1 (FilterDout_4__0__2), .A2 (
         FilterWR), .B0 (FilterDout_3__0__2), .B1 (nx8210)) ;
    dff L0_3_L1_0_Fij_reg_Dout_3 (.Q (FilterDout_3__0__3), .QB (\$dummy [155]), 
        .D (nx3531), .CLK (CLK)) ;
    ao32 ix3532 (.Y (nx3531), .A0 (nx8120), .A1 (FilterDout_4__0__3), .A2 (
         FilterWR), .B0 (FilterDout_3__0__3), .B1 (nx8210)) ;
    dff L0_3_L1_0_Fij_reg_Dout_4 (.Q (FilterDout_3__0__4), .QB (\$dummy [156]), 
        .D (nx3541), .CLK (CLK)) ;
    ao32 ix3542 (.Y (nx3541), .A0 (nx8120), .A1 (FilterDout_4__0__4), .A2 (
         FilterWR), .B0 (FilterDout_3__0__4), .B1 (nx8210)) ;
    dff L0_3_L1_0_Fij_reg_Dout_5 (.Q (FilterDout_3__0__5), .QB (\$dummy [157]), 
        .D (nx3551), .CLK (CLK)) ;
    ao32 ix3552 (.Y (nx3551), .A0 (nx8122), .A1 (FilterDout_4__0__5), .A2 (
         FilterWR), .B0 (FilterDout_3__0__5), .B1 (nx8210)) ;
    dff L0_3_L1_0_Fij_reg_Dout_6 (.Q (FilterDout_3__0__6), .QB (\$dummy [158]), 
        .D (nx3561), .CLK (CLK)) ;
    ao32 ix3562 (.Y (nx3561), .A0 (nx8122), .A1 (FilterDout_4__0__6), .A2 (
         FilterWR), .B0 (FilterDout_3__0__6), .B1 (nx8210)) ;
    dff L0_3_L1_0_Fij_reg_Dout_7 (.Q (FilterDout_3__0__7), .QB (\$dummy [159]), 
        .D (nx3571), .CLK (CLK)) ;
    ao32 ix3572 (.Y (nx3571), .A0 (nx8122), .A1 (FilterDout_4__0__7), .A2 (
         FilterWR), .B0 (FilterDout_3__0__7), .B1 (nx8210)) ;
    oai21 ix3662 (.Y (nx3661), .A0 (nx7259), .A1 (nx7982), .B0 (nx7261)) ;
    dff L0_2_L1_4_Fij_reg_Dout_0 (.Q (FilterDout_2__4__0), .QB (nx7259), .D (
        nx3661), .CLK (CLK)) ;
    oai21 ix3672 (.Y (nx3671), .A0 (nx7265), .A1 (nx7982), .B0 (nx7267)) ;
    dff L0_2_L1_4_Fij_reg_Dout_1 (.Q (FilterDout_2__4__1), .QB (nx7265), .D (
        nx3671), .CLK (CLK)) ;
    oai21 ix3682 (.Y (nx3681), .A0 (nx7271), .A1 (nx7984), .B0 (nx7273)) ;
    dff L0_2_L1_4_Fij_reg_Dout_2 (.Q (FilterDout_2__4__2), .QB (nx7271), .D (
        nx3681), .CLK (CLK)) ;
    oai21 ix3692 (.Y (nx3691), .A0 (nx7277), .A1 (nx7984), .B0 (nx7279)) ;
    dff L0_2_L1_4_Fij_reg_Dout_3 (.Q (FilterDout_2__4__3), .QB (nx7277), .D (
        nx3691), .CLK (CLK)) ;
    oai21 ix3702 (.Y (nx3701), .A0 (nx7283), .A1 (nx7984), .B0 (nx7285)) ;
    dff L0_2_L1_4_Fij_reg_Dout_4 (.Q (FilterDout_2__4__4), .QB (nx7283), .D (
        nx3701), .CLK (CLK)) ;
    oai21 ix3712 (.Y (nx3711), .A0 (nx7289), .A1 (nx7986), .B0 (nx7291)) ;
    dff L0_2_L1_4_Fij_reg_Dout_5 (.Q (FilterDout_2__4__5), .QB (nx7289), .D (
        nx3711), .CLK (CLK)) ;
    oai21 ix3722 (.Y (nx3721), .A0 (nx7295), .A1 (nx7986), .B0 (nx7297)) ;
    dff L0_2_L1_4_Fij_reg_Dout_6 (.Q (FilterDout_2__4__6), .QB (nx7295), .D (
        nx3721), .CLK (CLK)) ;
    oai21 ix3732 (.Y (nx3731), .A0 (nx7301), .A1 (nx7986), .B0 (nx7303)) ;
    dff L0_2_L1_4_Fij_reg_Dout_7 (.Q (FilterDout_2__4__7), .QB (nx7301), .D (
        nx3731), .CLK (CLK)) ;
    oai21 ix3822 (.Y (nx3821), .A0 (nx7307), .A1 (nx7986), .B0 (nx7309)) ;
    dff L0_2_L1_3_Fij_reg_Dout_0 (.Q (FilterDout_2__3__0), .QB (nx7307), .D (
        nx3821), .CLK (CLK)) ;
    oai21 ix3832 (.Y (nx3831), .A0 (nx7313), .A1 (nx7988), .B0 (nx7315)) ;
    dff L0_2_L1_3_Fij_reg_Dout_1 (.Q (FilterDout_2__3__1), .QB (nx7313), .D (
        nx3831), .CLK (CLK)) ;
    oai21 ix3842 (.Y (nx3841), .A0 (nx7319), .A1 (nx7988), .B0 (nx7321)) ;
    dff L0_2_L1_3_Fij_reg_Dout_2 (.Q (FilterDout_2__3__2), .QB (nx7319), .D (
        nx3841), .CLK (CLK)) ;
    oai21 ix3852 (.Y (nx3851), .A0 (nx7325), .A1 (nx7988), .B0 (nx7327)) ;
    dff L0_2_L1_3_Fij_reg_Dout_3 (.Q (FilterDout_2__3__3), .QB (nx7325), .D (
        nx3851), .CLK (CLK)) ;
    oai21 ix3862 (.Y (nx3861), .A0 (nx7331), .A1 (nx7990), .B0 (nx7333)) ;
    dff L0_2_L1_3_Fij_reg_Dout_4 (.Q (FilterDout_2__3__4), .QB (nx7331), .D (
        nx3861), .CLK (CLK)) ;
    oai21 ix3872 (.Y (nx3871), .A0 (nx7337), .A1 (nx7990), .B0 (nx7339)) ;
    dff L0_2_L1_3_Fij_reg_Dout_5 (.Q (FilterDout_2__3__5), .QB (nx7337), .D (
        nx3871), .CLK (CLK)) ;
    oai21 ix3882 (.Y (nx3881), .A0 (nx7343), .A1 (nx7990), .B0 (nx7345)) ;
    dff L0_2_L1_3_Fij_reg_Dout_6 (.Q (FilterDout_2__3__6), .QB (nx7343), .D (
        nx3881), .CLK (CLK)) ;
    oai21 ix3892 (.Y (nx3891), .A0 (nx7349), .A1 (nx7990), .B0 (nx7351)) ;
    dff L0_2_L1_3_Fij_reg_Dout_7 (.Q (FilterDout_2__3__7), .QB (nx7349), .D (
        nx3891), .CLK (CLK)) ;
    dff L0_2_L1_2_Fij_reg_Dout_0 (.Q (FilterDout_2__2__0), .QB (\$dummy [160]), 
        .D (nx3981), .CLK (CLK)) ;
    ao32 ix3982 (.Y (nx3981), .A0 (nx8126), .A1 (FilterDout_3__2__0), .A2 (
         FilterWR), .B0 (FilterDout_2__2__0), .B1 (nx8210)) ;
    dff L0_2_L1_2_Fij_reg_Dout_1 (.Q (FilterDout_2__2__1), .QB (\$dummy [161]), 
        .D (nx3991), .CLK (CLK)) ;
    ao32 ix3992 (.Y (nx3991), .A0 (nx8126), .A1 (FilterDout_3__2__1), .A2 (
         FilterWR), .B0 (FilterDout_2__2__1), .B1 (nx8212)) ;
    dff L0_2_L1_2_Fij_reg_Dout_2 (.Q (FilterDout_2__2__2), .QB (\$dummy [162]), 
        .D (nx4001), .CLK (CLK)) ;
    ao32 ix4002 (.Y (nx4001), .A0 (nx8128), .A1 (FilterDout_3__2__2), .A2 (
         FilterWR), .B0 (FilterDout_2__2__2), .B1 (nx8212)) ;
    dff L0_2_L1_2_Fij_reg_Dout_3 (.Q (FilterDout_2__2__3), .QB (\$dummy [163]), 
        .D (nx4011), .CLK (CLK)) ;
    ao32 ix4012 (.Y (nx4011), .A0 (nx8128), .A1 (FilterDout_3__2__3), .A2 (
         FilterWR), .B0 (FilterDout_2__2__3), .B1 (nx8212)) ;
    dff L0_2_L1_2_Fij_reg_Dout_4 (.Q (FilterDout_2__2__4), .QB (\$dummy [164]), 
        .D (nx4021), .CLK (CLK)) ;
    ao32 ix4022 (.Y (nx4021), .A0 (nx8128), .A1 (FilterDout_3__2__4), .A2 (
         FilterWR), .B0 (FilterDout_2__2__4), .B1 (nx8212)) ;
    dff L0_2_L1_2_Fij_reg_Dout_5 (.Q (FilterDout_2__2__5), .QB (\$dummy [165]), 
        .D (nx4031), .CLK (CLK)) ;
    ao32 ix4032 (.Y (nx4031), .A0 (nx8128), .A1 (FilterDout_3__2__5), .A2 (
         FilterWR), .B0 (FilterDout_2__2__5), .B1 (nx8212)) ;
    dff L0_2_L1_2_Fij_reg_Dout_6 (.Q (FilterDout_2__2__6), .QB (\$dummy [166]), 
        .D (nx4041), .CLK (CLK)) ;
    ao32 ix4042 (.Y (nx4041), .A0 (nx8128), .A1 (FilterDout_3__2__6), .A2 (
         FilterWR), .B0 (FilterDout_2__2__6), .B1 (nx8212)) ;
    dff L0_2_L1_2_Fij_reg_Dout_7 (.Q (FilterDout_2__2__7), .QB (\$dummy [167]), 
        .D (nx4051), .CLK (CLK)) ;
    ao32 ix4052 (.Y (nx4051), .A0 (nx8128), .A1 (FilterDout_3__2__7), .A2 (
         FilterWR), .B0 (FilterDout_2__2__7), .B1 (nx8212)) ;
    dff L0_2_L1_1_Fij_reg_Dout_0 (.Q (FilterDout_2__1__0), .QB (\$dummy [168]), 
        .D (nx4141), .CLK (CLK)) ;
    ao32 ix4142 (.Y (nx4141), .A0 (nx8128), .A1 (FilterDout_3__1__0), .A2 (
         FilterWR), .B0 (FilterDout_2__1__0), .B1 (nx8214)) ;
    dff L0_2_L1_1_Fij_reg_Dout_1 (.Q (FilterDout_2__1__1), .QB (\$dummy [169]), 
        .D (nx4151), .CLK (CLK)) ;
    ao32 ix4152 (.Y (nx4151), .A0 (nx8130), .A1 (FilterDout_3__1__1), .A2 (
         FilterWR), .B0 (FilterDout_2__1__1), .B1 (nx8214)) ;
    dff L0_2_L1_1_Fij_reg_Dout_2 (.Q (FilterDout_2__1__2), .QB (\$dummy [170]), 
        .D (nx4161), .CLK (CLK)) ;
    ao32 ix4162 (.Y (nx4161), .A0 (nx8130), .A1 (FilterDout_3__1__2), .A2 (
         FilterWR), .B0 (FilterDout_2__1__2), .B1 (nx8214)) ;
    dff L0_2_L1_1_Fij_reg_Dout_3 (.Q (FilterDout_2__1__3), .QB (\$dummy [171]), 
        .D (nx4171), .CLK (CLK)) ;
    ao32 ix4172 (.Y (nx4171), .A0 (nx8130), .A1 (FilterDout_3__1__3), .A2 (
         FilterWR), .B0 (FilterDout_2__1__3), .B1 (nx8214)) ;
    dff L0_2_L1_1_Fij_reg_Dout_4 (.Q (FilterDout_2__1__4), .QB (\$dummy [172]), 
        .D (nx4181), .CLK (CLK)) ;
    ao32 ix4182 (.Y (nx4181), .A0 (nx8130), .A1 (FilterDout_3__1__4), .A2 (
         FilterWR), .B0 (FilterDout_2__1__4), .B1 (nx8214)) ;
    dff L0_2_L1_1_Fij_reg_Dout_5 (.Q (FilterDout_2__1__5), .QB (\$dummy [173]), 
        .D (nx4191), .CLK (CLK)) ;
    ao32 ix4192 (.Y (nx4191), .A0 (nx8130), .A1 (FilterDout_3__1__5), .A2 (
         FilterWR), .B0 (FilterDout_2__1__5), .B1 (nx8214)) ;
    dff L0_2_L1_1_Fij_reg_Dout_6 (.Q (FilterDout_2__1__6), .QB (\$dummy [174]), 
        .D (nx4201), .CLK (CLK)) ;
    ao32 ix4202 (.Y (nx4201), .A0 (nx8130), .A1 (FilterDout_3__1__6), .A2 (
         FilterWR), .B0 (FilterDout_2__1__6), .B1 (nx8214)) ;
    dff L0_2_L1_1_Fij_reg_Dout_7 (.Q (FilterDout_2__1__7), .QB (\$dummy [175]), 
        .D (nx4211), .CLK (CLK)) ;
    ao32 ix4212 (.Y (nx4211), .A0 (nx8130), .A1 (FilterDout_3__1__7), .A2 (
         FilterWR), .B0 (FilterDout_2__1__7), .B1 (nx8216)) ;
    dff L0_2_L1_0_Fij_reg_Dout_0 (.Q (FilterDout_2__0__0), .QB (\$dummy [176]), 
        .D (nx4301), .CLK (CLK)) ;
    ao32 ix4302 (.Y (nx4301), .A0 (nx8132), .A1 (FilterDout_3__0__0), .A2 (
         FilterWR), .B0 (FilterDout_2__0__0), .B1 (nx8216)) ;
    dff L0_2_L1_0_Fij_reg_Dout_1 (.Q (FilterDout_2__0__1), .QB (\$dummy [177]), 
        .D (nx4311), .CLK (CLK)) ;
    ao32 ix4312 (.Y (nx4311), .A0 (nx8132), .A1 (FilterDout_3__0__1), .A2 (
         FilterWR), .B0 (FilterDout_2__0__1), .B1 (nx8216)) ;
    dff L0_2_L1_0_Fij_reg_Dout_2 (.Q (FilterDout_2__0__2), .QB (\$dummy [178]), 
        .D (nx4321), .CLK (CLK)) ;
    ao32 ix4322 (.Y (nx4321), .A0 (nx8132), .A1 (FilterDout_3__0__2), .A2 (
         FilterWR), .B0 (FilterDout_2__0__2), .B1 (nx8216)) ;
    dff L0_2_L1_0_Fij_reg_Dout_3 (.Q (FilterDout_2__0__3), .QB (\$dummy [179]), 
        .D (nx4331), .CLK (CLK)) ;
    ao32 ix4332 (.Y (nx4331), .A0 (nx8132), .A1 (FilterDout_3__0__3), .A2 (
         FilterWR), .B0 (FilterDout_2__0__3), .B1 (nx8216)) ;
    dff L0_2_L1_0_Fij_reg_Dout_4 (.Q (FilterDout_2__0__4), .QB (\$dummy [180]), 
        .D (nx4341), .CLK (CLK)) ;
    ao32 ix4342 (.Y (nx4341), .A0 (nx8132), .A1 (FilterDout_3__0__4), .A2 (
         FilterWR), .B0 (FilterDout_2__0__4), .B1 (nx8216)) ;
    dff L0_2_L1_0_Fij_reg_Dout_5 (.Q (FilterDout_2__0__5), .QB (\$dummy [181]), 
        .D (nx4351), .CLK (CLK)) ;
    ao32 ix4352 (.Y (nx4351), .A0 (nx8132), .A1 (FilterDout_3__0__5), .A2 (
         FilterWR), .B0 (FilterDout_2__0__5), .B1 (nx8216)) ;
    dff L0_2_L1_0_Fij_reg_Dout_6 (.Q (FilterDout_2__0__6), .QB (\$dummy [182]), 
        .D (nx4361), .CLK (CLK)) ;
    ao32 ix4362 (.Y (nx4361), .A0 (nx8132), .A1 (FilterDout_3__0__6), .A2 (
         FilterWR), .B0 (FilterDout_2__0__6), .B1 (nx8218)) ;
    dff L0_2_L1_0_Fij_reg_Dout_7 (.Q (FilterDout_2__0__7), .QB (\$dummy [183]), 
        .D (nx4371), .CLK (CLK)) ;
    ao32 ix4372 (.Y (nx4371), .A0 (nx8134), .A1 (FilterDout_3__0__7), .A2 (
         FilterWR), .B0 (FilterDout_2__0__7), .B1 (nx8218)) ;
    oai21 ix4542 (.Y (nx4541), .A0 (nx7427), .A1 (nx7992), .B0 (nx7429)) ;
    dff L0_1_L1_4_Fij_reg_Dout_0 (.Q (FilterDout_1__4__0), .QB (nx7427), .D (
        nx4541), .CLK (CLK)) ;
    oai21 ix4552 (.Y (nx4551), .A0 (nx7433), .A1 (nx7992), .B0 (nx7435)) ;
    dff L0_1_L1_4_Fij_reg_Dout_1 (.Q (FilterDout_1__4__1), .QB (nx7433), .D (
        nx4551), .CLK (CLK)) ;
    oai21 ix4562 (.Y (nx4561), .A0 (nx7439), .A1 (nx7992), .B0 (nx7441)) ;
    dff L0_1_L1_4_Fij_reg_Dout_2 (.Q (FilterDout_1__4__2), .QB (nx7439), .D (
        nx4561), .CLK (CLK)) ;
    oai21 ix4572 (.Y (nx4571), .A0 (nx7445), .A1 (nx7994), .B0 (nx7447)) ;
    dff L0_1_L1_4_Fij_reg_Dout_3 (.Q (FilterDout_1__4__3), .QB (nx7445), .D (
        nx4571), .CLK (CLK)) ;
    oai21 ix4582 (.Y (nx4581), .A0 (nx7451), .A1 (nx7994), .B0 (nx7453)) ;
    dff L0_1_L1_4_Fij_reg_Dout_4 (.Q (FilterDout_1__4__4), .QB (nx7451), .D (
        nx4581), .CLK (CLK)) ;
    oai21 ix4592 (.Y (nx4591), .A0 (nx7457), .A1 (nx7994), .B0 (nx7459)) ;
    dff L0_1_L1_4_Fij_reg_Dout_5 (.Q (FilterDout_1__4__5), .QB (nx7457), .D (
        nx4591), .CLK (CLK)) ;
    oai21 ix4602 (.Y (nx4601), .A0 (nx7463), .A1 (nx7994), .B0 (nx7465)) ;
    dff L0_1_L1_4_Fij_reg_Dout_6 (.Q (FilterDout_1__4__6), .QB (nx7463), .D (
        nx4601), .CLK (CLK)) ;
    oai21 ix4612 (.Y (nx4611), .A0 (nx7469), .A1 (nx7996), .B0 (nx7471)) ;
    dff L0_1_L1_4_Fij_reg_Dout_7 (.Q (FilterDout_1__4__7), .QB (nx7469), .D (
        nx4611), .CLK (CLK)) ;
    oai21 ix4862 (.Y (nx4861), .A0 (nx7475), .A1 (nx7996), .B0 (nx7477)) ;
    dff L0_1_L1_3_Fij_reg_Dout_0 (.Q (FilterDout_1__3__0), .QB (nx7475), .D (
        nx4861), .CLK (CLK)) ;
    oai21 ix4872 (.Y (nx4871), .A0 (nx7481), .A1 (nx7996), .B0 (nx7483)) ;
    dff L0_1_L1_3_Fij_reg_Dout_1 (.Q (FilterDout_1__3__1), .QB (nx7481), .D (
        nx4871), .CLK (CLK)) ;
    oai21 ix4882 (.Y (nx4881), .A0 (nx7487), .A1 (nx7998), .B0 (nx7489)) ;
    dff L0_1_L1_3_Fij_reg_Dout_2 (.Q (FilterDout_1__3__2), .QB (nx7487), .D (
        nx4881), .CLK (CLK)) ;
    oai21 ix4892 (.Y (nx4891), .A0 (nx7493), .A1 (nx7998), .B0 (nx7495)) ;
    dff L0_1_L1_3_Fij_reg_Dout_3 (.Q (FilterDout_1__3__3), .QB (nx7493), .D (
        nx4891), .CLK (CLK)) ;
    oai21 ix4902 (.Y (nx4901), .A0 (nx7499), .A1 (nx7998), .B0 (nx7501)) ;
    dff L0_1_L1_3_Fij_reg_Dout_4 (.Q (FilterDout_1__3__4), .QB (nx7499), .D (
        nx4901), .CLK (CLK)) ;
    oai21 ix4912 (.Y (nx4911), .A0 (nx7505), .A1 (nx7998), .B0 (nx7507)) ;
    dff L0_1_L1_3_Fij_reg_Dout_5 (.Q (FilterDout_1__3__5), .QB (nx7505), .D (
        nx4911), .CLK (CLK)) ;
    oai21 ix4922 (.Y (nx4921), .A0 (nx7511), .A1 (nx8000), .B0 (nx7513)) ;
    dff L0_1_L1_3_Fij_reg_Dout_6 (.Q (FilterDout_1__3__6), .QB (nx7511), .D (
        nx4921), .CLK (CLK)) ;
    oai21 ix4932 (.Y (nx4931), .A0 (nx7517), .A1 (nx8000), .B0 (nx7519)) ;
    dff L0_1_L1_3_Fij_reg_Dout_7 (.Q (FilterDout_1__3__7), .QB (nx7517), .D (
        nx4931), .CLK (CLK)) ;
    oai21 ix5182 (.Y (nx5181), .A0 (nx7523), .A1 (nx8000), .B0 (nx7525)) ;
    dff L0_1_L1_2_Fij_reg_Dout_0 (.Q (FilterDout_1__2__0), .QB (nx7523), .D (
        nx5181), .CLK (CLK)) ;
    nand03 ix7526 (.Y (nx7525), .A0 (nx8138), .A1 (FilterDout_2__2__0), .A2 (
           nx8000)) ;
    oai21 ix5192 (.Y (nx5191), .A0 (nx7529), .A1 (nx8002), .B0 (nx7531)) ;
    dff L0_1_L1_2_Fij_reg_Dout_1 (.Q (FilterDout_1__2__1), .QB (nx7529), .D (
        nx5191), .CLK (CLK)) ;
    nand03 ix7532 (.Y (nx7531), .A0 (nx8138), .A1 (FilterDout_2__2__1), .A2 (
           nx8002)) ;
    oai21 ix5202 (.Y (nx5201), .A0 (nx7535), .A1 (nx8002), .B0 (nx7537)) ;
    dff L0_1_L1_2_Fij_reg_Dout_2 (.Q (FilterDout_1__2__2), .QB (nx7535), .D (
        nx5201), .CLK (CLK)) ;
    nand03 ix7538 (.Y (nx7537), .A0 (nx8138), .A1 (FilterDout_2__2__2), .A2 (
           nx8002)) ;
    oai21 ix5212 (.Y (nx5211), .A0 (nx7541), .A1 (nx8002), .B0 (nx7543)) ;
    dff L0_1_L1_2_Fij_reg_Dout_3 (.Q (FilterDout_1__2__3), .QB (nx7541), .D (
        nx5211), .CLK (CLK)) ;
    nand03 ix7544 (.Y (nx7543), .A0 (nx8138), .A1 (FilterDout_2__2__3), .A2 (
           nx8002)) ;
    oai21 ix5222 (.Y (nx5221), .A0 (nx7547), .A1 (nx8002), .B0 (nx7549)) ;
    dff L0_1_L1_2_Fij_reg_Dout_4 (.Q (FilterDout_1__2__4), .QB (nx7547), .D (
        nx5221), .CLK (CLK)) ;
    nand03 ix7550 (.Y (nx7549), .A0 (nx8140), .A1 (FilterDout_2__2__4), .A2 (
           nx8004)) ;
    oai21 ix5232 (.Y (nx5231), .A0 (nx7553), .A1 (nx8004), .B0 (nx7555)) ;
    dff L0_1_L1_2_Fij_reg_Dout_5 (.Q (FilterDout_1__2__5), .QB (nx7553), .D (
        nx5231), .CLK (CLK)) ;
    nand03 ix7556 (.Y (nx7555), .A0 (nx8140), .A1 (FilterDout_2__2__5), .A2 (
           nx8004)) ;
    oai21 ix5242 (.Y (nx5241), .A0 (nx7559), .A1 (nx8004), .B0 (nx7561)) ;
    dff L0_1_L1_2_Fij_reg_Dout_6 (.Q (FilterDout_1__2__6), .QB (nx7559), .D (
        nx5241), .CLK (CLK)) ;
    nand03 ix7562 (.Y (nx7561), .A0 (nx8140), .A1 (FilterDout_2__2__6), .A2 (
           nx8004)) ;
    oai21 ix5252 (.Y (nx5251), .A0 (nx7565), .A1 (nx8004), .B0 (nx7567)) ;
    dff L0_1_L1_2_Fij_reg_Dout_7 (.Q (FilterDout_1__2__7), .QB (nx7565), .D (
        nx5251), .CLK (CLK)) ;
    nand03 ix7568 (.Y (nx7567), .A0 (nx8140), .A1 (FilterDout_2__2__7), .A2 (
           nx8004)) ;
    oai21 ix5502 (.Y (nx5501), .A0 (nx7571), .A1 (nx8006), .B0 (nx7573)) ;
    dff L0_1_L1_1_Fij_reg_Dout_0 (.Q (FilterDout_1__1__0), .QB (nx7571), .D (
        nx5501), .CLK (CLK)) ;
    nand03 ix7574 (.Y (nx7573), .A0 (nx8140), .A1 (FilterDout_2__1__0), .A2 (
           nx8006)) ;
    oai21 ix5512 (.Y (nx5511), .A0 (nx7577), .A1 (nx8006), .B0 (nx7579)) ;
    dff L0_1_L1_1_Fij_reg_Dout_1 (.Q (FilterDout_1__1__1), .QB (nx7577), .D (
        nx5511), .CLK (CLK)) ;
    nand03 ix7580 (.Y (nx7579), .A0 (nx8140), .A1 (FilterDout_2__1__1), .A2 (
           nx8006)) ;
    oai21 ix5522 (.Y (nx5521), .A0 (nx7583), .A1 (nx8006), .B0 (nx7585)) ;
    dff L0_1_L1_1_Fij_reg_Dout_2 (.Q (FilterDout_1__1__2), .QB (nx7583), .D (
        nx5521), .CLK (CLK)) ;
    nand03 ix7586 (.Y (nx7585), .A0 (nx8140), .A1 (FilterDout_2__1__2), .A2 (
           nx8006)) ;
    oai21 ix5532 (.Y (nx5531), .A0 (nx7589), .A1 (nx8006), .B0 (nx7591)) ;
    dff L0_1_L1_1_Fij_reg_Dout_3 (.Q (FilterDout_1__1__3), .QB (nx7589), .D (
        nx5531), .CLK (CLK)) ;
    nand03 ix7592 (.Y (nx7591), .A0 (nx8142), .A1 (FilterDout_2__1__3), .A2 (
           nx8008)) ;
    oai21 ix5542 (.Y (nx5541), .A0 (nx7595), .A1 (nx8008), .B0 (nx7597)) ;
    dff L0_1_L1_1_Fij_reg_Dout_4 (.Q (FilterDout_1__1__4), .QB (nx7595), .D (
        nx5541), .CLK (CLK)) ;
    nand03 ix7598 (.Y (nx7597), .A0 (nx8142), .A1 (FilterDout_2__1__4), .A2 (
           nx8008)) ;
    oai21 ix5552 (.Y (nx5551), .A0 (nx7601), .A1 (nx8008), .B0 (nx7603)) ;
    dff L0_1_L1_1_Fij_reg_Dout_5 (.Q (FilterDout_1__1__5), .QB (nx7601), .D (
        nx5551), .CLK (CLK)) ;
    nand03 ix7604 (.Y (nx7603), .A0 (nx8142), .A1 (FilterDout_2__1__5), .A2 (
           nx8008)) ;
    oai21 ix5562 (.Y (nx5561), .A0 (nx7607), .A1 (nx8008), .B0 (nx7609)) ;
    dff L0_1_L1_1_Fij_reg_Dout_6 (.Q (FilterDout_1__1__6), .QB (nx7607), .D (
        nx5561), .CLK (CLK)) ;
    nand03 ix7610 (.Y (nx7609), .A0 (nx8142), .A1 (FilterDout_2__1__6), .A2 (
           nx8008)) ;
    oai21 ix5572 (.Y (nx5571), .A0 (nx7613), .A1 (nx8010), .B0 (nx7615)) ;
    dff L0_1_L1_1_Fij_reg_Dout_7 (.Q (FilterDout_1__1__7), .QB (nx7613), .D (
        nx5571), .CLK (CLK)) ;
    nand03 ix7616 (.Y (nx7615), .A0 (nx8142), .A1 (FilterDout_2__1__7), .A2 (
           nx8010)) ;
    oai21 ix5822 (.Y (nx5821), .A0 (nx7619), .A1 (nx8010), .B0 (nx7621)) ;
    dff L0_1_L1_0_Fij_reg_Dout_0 (.Q (FilterDout_1__0__0), .QB (nx7619), .D (
        nx5821), .CLK (CLK)) ;
    nand03 ix7622 (.Y (nx7621), .A0 (nx8142), .A1 (FilterDout_2__0__0), .A2 (
           nx8010)) ;
    oai21 ix5832 (.Y (nx5831), .A0 (nx7625), .A1 (nx8010), .B0 (nx7627)) ;
    dff L0_1_L1_0_Fij_reg_Dout_1 (.Q (FilterDout_1__0__1), .QB (nx7625), .D (
        nx5831), .CLK (CLK)) ;
    nand03 ix7628 (.Y (nx7627), .A0 (nx8142), .A1 (FilterDout_2__0__1), .A2 (
           nx8010)) ;
    oai21 ix5842 (.Y (nx5841), .A0 (nx7631), .A1 (nx8010), .B0 (nx7633)) ;
    dff L0_1_L1_0_Fij_reg_Dout_2 (.Q (FilterDout_1__0__2), .QB (nx7631), .D (
        nx5841), .CLK (CLK)) ;
    nand03 ix7634 (.Y (nx7633), .A0 (nx8144), .A1 (FilterDout_2__0__2), .A2 (
           nx8012)) ;
    oai21 ix5852 (.Y (nx5851), .A0 (nx7637), .A1 (nx8012), .B0 (nx7639)) ;
    dff L0_1_L1_0_Fij_reg_Dout_3 (.Q (FilterDout_1__0__3), .QB (nx7637), .D (
        nx5851), .CLK (CLK)) ;
    nand03 ix7640 (.Y (nx7639), .A0 (nx8144), .A1 (FilterDout_2__0__3), .A2 (
           nx8012)) ;
    oai21 ix5862 (.Y (nx5861), .A0 (nx7643), .A1 (nx8012), .B0 (nx7645)) ;
    dff L0_1_L1_0_Fij_reg_Dout_4 (.Q (FilterDout_1__0__4), .QB (nx7643), .D (
        nx5861), .CLK (CLK)) ;
    nand03 ix7646 (.Y (nx7645), .A0 (nx8144), .A1 (FilterDout_2__0__4), .A2 (
           nx8012)) ;
    oai21 ix5872 (.Y (nx5871), .A0 (nx7649), .A1 (nx8012), .B0 (nx7651)) ;
    dff L0_1_L1_0_Fij_reg_Dout_5 (.Q (FilterDout_1__0__5), .QB (nx7649), .D (
        nx5871), .CLK (CLK)) ;
    nand03 ix7652 (.Y (nx7651), .A0 (nx8144), .A1 (FilterDout_2__0__5), .A2 (
           nx8012)) ;
    oai21 ix5882 (.Y (nx5881), .A0 (nx7655), .A1 (nx8014), .B0 (nx7657)) ;
    dff L0_1_L1_0_Fij_reg_Dout_6 (.Q (FilterDout_1__0__6), .QB (nx7655), .D (
        nx5881), .CLK (CLK)) ;
    nand03 ix7658 (.Y (nx7657), .A0 (nx8144), .A1 (FilterDout_2__0__6), .A2 (
           nx8014)) ;
    oai21 ix5892 (.Y (nx5891), .A0 (nx7661), .A1 (nx8014), .B0 (nx7663)) ;
    dff L0_1_L1_0_Fij_reg_Dout_7 (.Q (FilterDout_1__0__7), .QB (nx7661), .D (
        nx5891), .CLK (CLK)) ;
    nand03 ix7664 (.Y (nx7663), .A0 (nx8144), .A1 (FilterDout_2__0__7), .A2 (
           nx8014)) ;
    oai21 ix4622 (.Y (nx4621), .A0 (nx7667), .A1 (nx8014), .B0 (nx7669)) ;
    dff L0_0_L1_4_Fij_reg_Dout_0 (.Q (FilterDout_0__4__0), .QB (nx7667), .D (
        nx4621), .CLK (CLK)) ;
    oai21 ix4632 (.Y (nx4631), .A0 (nx7673), .A1 (nx8014), .B0 (nx7675)) ;
    dff L0_0_L1_4_Fij_reg_Dout_1 (.Q (FilterDout_0__4__1), .QB (nx7673), .D (
        nx4631), .CLK (CLK)) ;
    oai21 ix4642 (.Y (nx4641), .A0 (nx7679), .A1 (nx8016), .B0 (nx7681)) ;
    dff L0_0_L1_4_Fij_reg_Dout_2 (.Q (FilterDout_0__4__2), .QB (nx7679), .D (
        nx4641), .CLK (CLK)) ;
    oai21 ix4652 (.Y (nx4651), .A0 (nx7685), .A1 (nx8016), .B0 (nx7687)) ;
    dff L0_0_L1_4_Fij_reg_Dout_3 (.Q (FilterDout_0__4__3), .QB (nx7685), .D (
        nx4651), .CLK (CLK)) ;
    oai21 ix4662 (.Y (nx4661), .A0 (nx7691), .A1 (nx8016), .B0 (nx7693)) ;
    dff L0_0_L1_4_Fij_reg_Dout_4 (.Q (FilterDout_0__4__4), .QB (nx7691), .D (
        nx4661), .CLK (CLK)) ;
    oai21 ix4672 (.Y (nx4671), .A0 (nx7697), .A1 (nx8018), .B0 (nx7699)) ;
    dff L0_0_L1_4_Fij_reg_Dout_5 (.Q (FilterDout_0__4__5), .QB (nx7697), .D (
        nx4671), .CLK (CLK)) ;
    oai21 ix4682 (.Y (nx4681), .A0 (nx7703), .A1 (nx8018), .B0 (nx7705)) ;
    dff L0_0_L1_4_Fij_reg_Dout_6 (.Q (FilterDout_0__4__6), .QB (nx7703), .D (
        nx4681), .CLK (CLK)) ;
    oai21 ix4692 (.Y (nx4691), .A0 (nx7709), .A1 (nx8018), .B0 (nx7711)) ;
    dff L0_0_L1_4_Fij_reg_Dout_7 (.Q (FilterDout_0__4__7), .QB (nx7709), .D (
        nx4691), .CLK (CLK)) ;
    oai21 ix4942 (.Y (nx4941), .A0 (nx7715), .A1 (nx8018), .B0 (nx7717)) ;
    dff L0_0_L1_3_Fij_reg_Dout_0 (.Q (FilterDout_0__3__0), .QB (nx7715), .D (
        nx4941), .CLK (CLK)) ;
    oai21 ix4952 (.Y (nx4951), .A0 (nx7721), .A1 (nx8020), .B0 (nx7723)) ;
    dff L0_0_L1_3_Fij_reg_Dout_1 (.Q (FilterDout_0__3__1), .QB (nx7721), .D (
        nx4951), .CLK (CLK)) ;
    oai21 ix4962 (.Y (nx4961), .A0 (nx7727), .A1 (nx8020), .B0 (nx7729)) ;
    dff L0_0_L1_3_Fij_reg_Dout_2 (.Q (FilterDout_0__3__2), .QB (nx7727), .D (
        nx4961), .CLK (CLK)) ;
    oai21 ix4972 (.Y (nx4971), .A0 (nx7733), .A1 (nx8020), .B0 (nx7735)) ;
    dff L0_0_L1_3_Fij_reg_Dout_3 (.Q (FilterDout_0__3__3), .QB (nx7733), .D (
        nx4971), .CLK (CLK)) ;
    oai21 ix4982 (.Y (nx4981), .A0 (nx7739), .A1 (nx8022), .B0 (nx7741)) ;
    dff L0_0_L1_3_Fij_reg_Dout_4 (.Q (FilterDout_0__3__4), .QB (nx7739), .D (
        nx4981), .CLK (CLK)) ;
    oai21 ix4992 (.Y (nx4991), .A0 (nx7745), .A1 (nx8022), .B0 (nx7747)) ;
    dff L0_0_L1_3_Fij_reg_Dout_5 (.Q (FilterDout_0__3__5), .QB (nx7745), .D (
        nx4991), .CLK (CLK)) ;
    oai21 ix5002 (.Y (nx5001), .A0 (nx7751), .A1 (nx8022), .B0 (nx7753)) ;
    dff L0_0_L1_3_Fij_reg_Dout_6 (.Q (FilterDout_0__3__6), .QB (nx7751), .D (
        nx5001), .CLK (CLK)) ;
    oai21 ix5012 (.Y (nx5011), .A0 (nx7757), .A1 (nx8022), .B0 (nx7759)) ;
    dff L0_0_L1_3_Fij_reg_Dout_7 (.Q (FilterDout_0__3__7), .QB (nx7757), .D (
        nx5011), .CLK (CLK)) ;
    oai21 ix5262 (.Y (nx5261), .A0 (nx7763), .A1 (nx8024), .B0 (nx7765)) ;
    dff L0_0_L1_2_Fij_reg_Dout_0 (.Q (FilterDout_0__2__0), .QB (nx7763), .D (
        nx5261), .CLK (CLK)) ;
    oai21 ix5272 (.Y (nx5271), .A0 (nx7769), .A1 (nx8024), .B0 (nx7771)) ;
    dff L0_0_L1_2_Fij_reg_Dout_1 (.Q (FilterDout_0__2__1), .QB (nx7769), .D (
        nx5271), .CLK (CLK)) ;
    oai21 ix5282 (.Y (nx5281), .A0 (nx7775), .A1 (nx8024), .B0 (nx7777)) ;
    dff L0_0_L1_2_Fij_reg_Dout_2 (.Q (FilterDout_0__2__2), .QB (nx7775), .D (
        nx5281), .CLK (CLK)) ;
    oai21 ix5292 (.Y (nx5291), .A0 (nx7781), .A1 (nx8026), .B0 (nx7783)) ;
    dff L0_0_L1_2_Fij_reg_Dout_3 (.Q (FilterDout_0__2__3), .QB (nx7781), .D (
        nx5291), .CLK (CLK)) ;
    oai21 ix5302 (.Y (nx5301), .A0 (nx7787), .A1 (nx8026), .B0 (nx7789)) ;
    dff L0_0_L1_2_Fij_reg_Dout_4 (.Q (FilterDout_0__2__4), .QB (nx7787), .D (
        nx5301), .CLK (CLK)) ;
    oai21 ix5312 (.Y (nx5311), .A0 (nx7793), .A1 (nx8026), .B0 (nx7795)) ;
    dff L0_0_L1_2_Fij_reg_Dout_5 (.Q (FilterDout_0__2__5), .QB (nx7793), .D (
        nx5311), .CLK (CLK)) ;
    oai21 ix5322 (.Y (nx5321), .A0 (nx7799), .A1 (nx8026), .B0 (nx7801)) ;
    dff L0_0_L1_2_Fij_reg_Dout_6 (.Q (FilterDout_0__2__6), .QB (nx7799), .D (
        nx5321), .CLK (CLK)) ;
    oai21 ix5332 (.Y (nx5331), .A0 (nx7805), .A1 (nx8028), .B0 (nx7807)) ;
    dff L0_0_L1_2_Fij_reg_Dout_7 (.Q (FilterDout_0__2__7), .QB (nx7805), .D (
        nx5331), .CLK (CLK)) ;
    oai21 ix5582 (.Y (nx5581), .A0 (nx7811), .A1 (nx8028), .B0 (nx7813)) ;
    dff L0_0_L1_1_Fij_reg_Dout_0 (.Q (FilterDout_0__1__0), .QB (nx7811), .D (
        nx5581), .CLK (CLK)) ;
    oai21 ix5592 (.Y (nx5591), .A0 (nx7817), .A1 (nx8028), .B0 (nx7819)) ;
    dff L0_0_L1_1_Fij_reg_Dout_1 (.Q (FilterDout_0__1__1), .QB (nx7817), .D (
        nx5591), .CLK (CLK)) ;
    oai21 ix5602 (.Y (nx5601), .A0 (nx7823), .A1 (nx8030), .B0 (nx7825)) ;
    dff L0_0_L1_1_Fij_reg_Dout_2 (.Q (FilterDout_0__1__2), .QB (nx7823), .D (
        nx5601), .CLK (CLK)) ;
    oai21 ix5612 (.Y (nx5611), .A0 (nx7829), .A1 (nx8030), .B0 (nx7831)) ;
    dff L0_0_L1_1_Fij_reg_Dout_3 (.Q (FilterDout_0__1__3), .QB (nx7829), .D (
        nx5611), .CLK (CLK)) ;
    oai21 ix5622 (.Y (nx5621), .A0 (nx7835), .A1 (nx8030), .B0 (nx7837)) ;
    dff L0_0_L1_1_Fij_reg_Dout_4 (.Q (FilterDout_0__1__4), .QB (nx7835), .D (
        nx5621), .CLK (CLK)) ;
    oai21 ix5632 (.Y (nx5631), .A0 (nx7841), .A1 (nx8030), .B0 (nx7843)) ;
    dff L0_0_L1_1_Fij_reg_Dout_5 (.Q (FilterDout_0__1__5), .QB (nx7841), .D (
        nx5631), .CLK (CLK)) ;
    oai21 ix5642 (.Y (nx5641), .A0 (nx7847), .A1 (nx8032), .B0 (nx7849)) ;
    dff L0_0_L1_1_Fij_reg_Dout_6 (.Q (FilterDout_0__1__6), .QB (nx7847), .D (
        nx5641), .CLK (CLK)) ;
    oai21 ix5652 (.Y (nx5651), .A0 (nx7853), .A1 (nx8032), .B0 (nx7855)) ;
    dff L0_0_L1_1_Fij_reg_Dout_7 (.Q (FilterDout_0__1__7), .QB (nx7853), .D (
        nx5651), .CLK (CLK)) ;
    oai21 ix5902 (.Y (nx5901), .A0 (nx7859), .A1 (nx8032), .B0 (nx7861)) ;
    dff L0_0_L1_0_Fij_reg_Dout_0 (.Q (FilterDout_0__0__0), .QB (nx7859), .D (
        nx5901), .CLK (CLK)) ;
    oai21 ix5912 (.Y (nx5911), .A0 (nx7865), .A1 (nx8034), .B0 (nx7867)) ;
    dff L0_0_L1_0_Fij_reg_Dout_1 (.Q (FilterDout_0__0__1), .QB (nx7865), .D (
        nx5911), .CLK (CLK)) ;
    oai21 ix5922 (.Y (nx5921), .A0 (nx7871), .A1 (nx8034), .B0 (nx7873)) ;
    dff L0_0_L1_0_Fij_reg_Dout_2 (.Q (FilterDout_0__0__2), .QB (nx7871), .D (
        nx5921), .CLK (CLK)) ;
    oai21 ix5932 (.Y (nx5931), .A0 (nx7877), .A1 (nx8034), .B0 (nx7879)) ;
    dff L0_0_L1_0_Fij_reg_Dout_3 (.Q (FilterDout_0__0__3), .QB (nx7877), .D (
        nx5931), .CLK (CLK)) ;
    oai21 ix5942 (.Y (nx5941), .A0 (nx7883), .A1 (nx8034), .B0 (nx7885)) ;
    dff L0_0_L1_0_Fij_reg_Dout_4 (.Q (FilterDout_0__0__4), .QB (nx7883), .D (
        nx5941), .CLK (CLK)) ;
    oai21 ix5952 (.Y (nx5951), .A0 (nx7889), .A1 (nx8036), .B0 (nx7891)) ;
    dff L0_0_L1_0_Fij_reg_Dout_5 (.Q (FilterDout_0__0__5), .QB (nx7889), .D (
        nx5951), .CLK (CLK)) ;
    oai21 ix5962 (.Y (nx5961), .A0 (nx7895), .A1 (nx8036), .B0 (nx7897)) ;
    dff L0_0_L1_0_Fij_reg_Dout_6 (.Q (FilterDout_0__0__6), .QB (nx7895), .D (
        nx5961), .CLK (CLK)) ;
    oai21 ix5972 (.Y (nx5971), .A0 (nx7901), .A1 (nx8036), .B0 (nx7903)) ;
    dff L0_0_L1_0_Fij_reg_Dout_7 (.Q (FilterDout_0__0__7), .QB (nx7901), .D (
        nx5971), .CLK (CLK)) ;
    inv02 ix167 (.Y (nx166), .A (nx6966)) ;
    inv02 ix83 (.Y (nx82), .A (nx6008)) ;
    inv02 ix7909 (.Y (nx7910), .A (nx8042)) ;
    inv02 ix7911 (.Y (nx7912), .A (nx8042)) ;
    inv02 ix7913 (.Y (nx7914), .A (nx8042)) ;
    inv02 ix7915 (.Y (nx7916), .A (nx8042)) ;
    inv02 ix7917 (.Y (nx7918), .A (nx8042)) ;
    inv02 ix7919 (.Y (nx7920), .A (nx8244)) ;
    inv02 ix7921 (.Y (nx7922), .A (nx8244)) ;
    inv02 ix7923 (.Y (nx7924), .A (nx8244)) ;
    inv02 ix7925 (.Y (nx7926), .A (nx8244)) ;
    inv02 ix7927 (.Y (nx7928), .A (nx8244)) ;
    inv02 ix7929 (.Y (nx7930), .A (nx8244)) ;
    inv02 ix7931 (.Y (nx7932), .A (nx8244)) ;
    inv02 ix7933 (.Y (nx7934), .A (nx8252)) ;
    inv02 ix7935 (.Y (nx7936), .A (nx8252)) ;
    inv02 ix7937 (.Y (nx7938), .A (nx8252)) ;
    inv02 ix7939 (.Y (nx7940), .A (nx8252)) ;
    inv02 ix7941 (.Y (nx7942), .A (nx8252)) ;
    inv02 ix7943 (.Y (nx7944), .A (nx8252)) ;
    inv02 ix7945 (.Y (nx7946), .A (nx8252)) ;
    inv02 ix7947 (.Y (nx7948), .A (nx8254)) ;
    inv02 ix7949 (.Y (nx7950), .A (nx8254)) ;
    inv02 ix7951 (.Y (nx7952), .A (nx8254)) ;
    inv02 ix7953 (.Y (nx7954), .A (nx8254)) ;
    inv02 ix7955 (.Y (nx7956), .A (nx8254)) ;
    inv02 ix7957 (.Y (nx7958), .A (nx8254)) ;
    inv02 ix7959 (.Y (nx7960), .A (nx8254)) ;
    inv02 ix7961 (.Y (nx7962), .A (nx8260)) ;
    inv02 ix7963 (.Y (nx7964), .A (nx8260)) ;
    inv02 ix7965 (.Y (nx7966), .A (nx8260)) ;
    inv02 ix7967 (.Y (nx7968), .A (nx8260)) ;
    inv02 ix7969 (.Y (nx7970), .A (nx8260)) ;
    inv02 ix7971 (.Y (nx7972), .A (nx8260)) ;
    inv02 ix7973 (.Y (nx7974), .A (nx8186)) ;
    inv02 ix7975 (.Y (nx7976), .A (nx8186)) ;
    inv02 ix7977 (.Y (nx7978), .A (nx8186)) ;
    inv02 ix7979 (.Y (nx7980), .A (nx8186)) ;
    inv02 ix7981 (.Y (nx7982), .A (nx8186)) ;
    inv02 ix7983 (.Y (nx7984), .A (nx8266)) ;
    inv02 ix7985 (.Y (nx7986), .A (nx8266)) ;
    inv02 ix7987 (.Y (nx7988), .A (nx8266)) ;
    inv02 ix7989 (.Y (nx7990), .A (nx8266)) ;
    inv02 ix7991 (.Y (nx7992), .A (nx8266)) ;
    inv02 ix7993 (.Y (nx7994), .A (nx8266)) ;
    inv02 ix7995 (.Y (nx7996), .A (nx8266)) ;
    inv02 ix7997 (.Y (nx7998), .A (nx8274)) ;
    inv02 ix7999 (.Y (nx8000), .A (nx8274)) ;
    inv02 ix8001 (.Y (nx8002), .A (nx8274)) ;
    inv02 ix8003 (.Y (nx8004), .A (nx8274)) ;
    inv02 ix8005 (.Y (nx8006), .A (nx8274)) ;
    inv02 ix8007 (.Y (nx8008), .A (nx8274)) ;
    inv02 ix8009 (.Y (nx8010), .A (nx8274)) ;
    inv02 ix8011 (.Y (nx8012), .A (nx8276)) ;
    inv02 ix8013 (.Y (nx8014), .A (nx8276)) ;
    inv02 ix8015 (.Y (nx8016), .A (nx8276)) ;
    inv02 ix8017 (.Y (nx8018), .A (nx8276)) ;
    inv02 ix8019 (.Y (nx8020), .A (nx8276)) ;
    inv02 ix8021 (.Y (nx8022), .A (nx8276)) ;
    inv02 ix8023 (.Y (nx8024), .A (nx8276)) ;
    inv02 ix8025 (.Y (nx8026), .A (nx8282)) ;
    inv02 ix8027 (.Y (nx8028), .A (nx8282)) ;
    inv02 ix8029 (.Y (nx8030), .A (nx8282)) ;
    inv02 ix8031 (.Y (nx8032), .A (nx8282)) ;
    inv02 ix8033 (.Y (nx8034), .A (nx8282)) ;
    inv02 ix8035 (.Y (nx8036), .A (nx8282)) ;
    inv02 ix8041 (.Y (nx8042), .A (nx8288)) ;
    inv02 ix8043 (.Y (nx8044), .A (nx8288)) ;
    inv02 ix8045 (.Y (nx8046), .A (nx8288)) ;
    inv02 ix8047 (.Y (nx8048), .A (nx8288)) ;
    inv02 ix8049 (.Y (nx8050), .A (nx8288)) ;
    inv02 ix8051 (.Y (nx8052), .A (RST)) ;
    inv02 ix8053 (.Y (nx8054), .A (RST)) ;
    inv02 ix8055 (.Y (nx8056), .A (RST)) ;
    inv02 ix8057 (.Y (nx8058), .A (RST)) ;
    inv02 ix8059 (.Y (nx8060), .A (RST)) ;
    inv02 ix8061 (.Y (nx8062), .A (RST)) ;
    inv02 ix8063 (.Y (nx8064), .A (RST)) ;
    inv02 ix8065 (.Y (nx8066), .A (RST)) ;
    inv02 ix8067 (.Y (nx8068), .A (RST)) ;
    inv02 ix8069 (.Y (nx8070), .A (RST)) ;
    inv02 ix8073 (.Y (nx8074), .A (RST)) ;
    inv02 ix8075 (.Y (nx8076), .A (RST)) ;
    inv02 ix8077 (.Y (nx8078), .A (RST)) ;
    inv02 ix8079 (.Y (nx8080), .A (RST)) ;
    inv02 ix8085 (.Y (nx8086), .A (RST)) ;
    inv02 ix8087 (.Y (nx8088), .A (RST)) ;
    inv02 ix8089 (.Y (nx8090), .A (RST)) ;
    inv02 ix8091 (.Y (nx8092), .A (RST)) ;
    inv02 ix8103 (.Y (nx8104), .A (RST)) ;
    inv02 ix8105 (.Y (nx8106), .A (RST)) ;
    inv02 ix8107 (.Y (nx8108), .A (RST)) ;
    inv02 ix8109 (.Y (nx8110), .A (RST)) ;
    inv02 ix8111 (.Y (nx8112), .A (RST)) ;
    inv02 ix8113 (.Y (nx8114), .A (RST)) ;
    inv02 ix8115 (.Y (nx8116), .A (RST)) ;
    inv02 ix8117 (.Y (nx8118), .A (RST)) ;
    inv02 ix8119 (.Y (nx8120), .A (RST)) ;
    inv02 ix8121 (.Y (nx8122), .A (RST)) ;
    inv02 ix8125 (.Y (nx8126), .A (RST)) ;
    inv02 ix8127 (.Y (nx8128), .A (RST)) ;
    inv02 ix8129 (.Y (nx8130), .A (RST)) ;
    inv02 ix8131 (.Y (nx8132), .A (RST)) ;
    inv02 ix8133 (.Y (nx8134), .A (RST)) ;
    inv02 ix8137 (.Y (nx8138), .A (RST)) ;
    inv02 ix8139 (.Y (nx8140), .A (RST)) ;
    inv02 ix8141 (.Y (nx8142), .A (RST)) ;
    inv02 ix8143 (.Y (nx8144), .A (RST)) ;
    inv02 ix8159 (.Y (nx8160), .A (nx8220)) ;
    inv02 ix8161 (.Y (nx8162), .A (nx8220)) ;
    inv02 ix8163 (.Y (nx8164), .A (nx8220)) ;
    inv02 ix8165 (.Y (nx8166), .A (nx8220)) ;
    inv02 ix8167 (.Y (nx8168), .A (nx8220)) ;
    inv02 ix8169 (.Y (nx8170), .A (nx8220)) ;
    inv02 ix8171 (.Y (nx8172), .A (nx8220)) ;
    inv02 ix8173 (.Y (nx8174), .A (nx8222)) ;
    inv02 ix8175 (.Y (nx8176), .A (nx8222)) ;
    inv02 ix8177 (.Y (nx8178), .A (nx8222)) ;
    inv02 ix8179 (.Y (nx8180), .A (nx8222)) ;
    inv02 ix8185 (.Y (nx8186), .A (nx8292)) ;
    inv02 ix8187 (.Y (nx8188), .A (nx8292)) ;
    inv02 ix8189 (.Y (nx8190), .A (nx8292)) ;
    inv02 ix8191 (.Y (nx8192), .A (nx8292)) ;
    inv02 ix8193 (.Y (nx8194), .A (nx8292)) ;
    inv02 ix8197 (.Y (nx8198), .A (nx8224)) ;
    inv02 ix8199 (.Y (nx8200), .A (nx8224)) ;
    inv02 ix8201 (.Y (nx8202), .A (nx8224)) ;
    inv02 ix8203 (.Y (nx8204), .A (nx8224)) ;
    inv02 ix8205 (.Y (nx8206), .A (nx8224)) ;
    inv02 ix8207 (.Y (nx8208), .A (nx8224)) ;
    inv02 ix8209 (.Y (nx8210), .A (nx8224)) ;
    inv02 ix8211 (.Y (nx8212), .A (nx8226)) ;
    inv02 ix8213 (.Y (nx8214), .A (nx8226)) ;
    inv02 ix8215 (.Y (nx8216), .A (nx8226)) ;
    inv02 ix8217 (.Y (nx8218), .A (nx8226)) ;
    inv02 ix8219 (.Y (nx8220), .A (nx6075)) ;
    inv02 ix8221 (.Y (nx8222), .A (nx6075)) ;
    inv02 ix8223 (.Y (nx8224), .A (nx7016)) ;
    inv02 ix8225 (.Y (nx8226), .A (nx7016)) ;
    mux21_ni ix1982 (.Y (nx1981), .A0 (WindowDout_4__4__0), .A1 (nx86), .S0 (
             nx8288)) ;
    mux21_ni ix1992 (.Y (nx1991), .A0 (WindowDout_4__4__1), .A1 (nx96), .S0 (
             nx8288)) ;
    mux21_ni ix2002 (.Y (nx2001), .A0 (WindowDout_4__4__2), .A1 (nx106), .S0 (
             nx8238)) ;
    mux21_ni ix2012 (.Y (nx2011), .A0 (WindowDout_4__4__3), .A1 (nx116), .S0 (
             nx8238)) ;
    mux21_ni ix2022 (.Y (nx2021), .A0 (WindowDout_4__4__4), .A1 (nx126), .S0 (
             nx8238)) ;
    mux21_ni ix2032 (.Y (nx2031), .A0 (WindowDout_4__4__5), .A1 (nx136), .S0 (
             nx8238)) ;
    mux21_ni ix2042 (.Y (nx2041), .A0 (WindowDout_4__4__6), .A1 (nx146), .S0 (
             nx8238)) ;
    mux21_ni ix2052 (.Y (nx2051), .A0 (WindowDout_4__4__7), .A1 (nx156), .S0 (
             nx8238)) ;
    mux21_ni ix2142 (.Y (nx2141), .A0 (WindowDout_4__3__0), .A1 (nx218), .S0 (
             nx8238)) ;
    mux21_ni ix2152 (.Y (nx2151), .A0 (WindowDout_4__3__1), .A1 (nx228), .S0 (
             nx82)) ;
    mux21_ni ix2162 (.Y (nx2161), .A0 (WindowDout_4__3__2), .A1 (nx238), .S0 (
             nx82)) ;
    mux21_ni ix2172 (.Y (nx2171), .A0 (WindowDout_4__3__3), .A1 (nx248), .S0 (
             nx82)) ;
    mux21_ni ix2182 (.Y (nx2181), .A0 (WindowDout_4__3__4), .A1 (nx258), .S0 (
             nx82)) ;
    mux21_ni ix2192 (.Y (nx2191), .A0 (WindowDout_4__3__5), .A1 (nx268), .S0 (
             nx82)) ;
    mux21_ni ix2202 (.Y (nx2201), .A0 (WindowDout_4__3__6), .A1 (nx278), .S0 (
             nx82)) ;
    mux21_ni ix2212 (.Y (nx2211), .A0 (WindowDout_4__3__7), .A1 (nx288), .S0 (
             nx82)) ;
    or03 ix6321 (.Y (nx6320), .A0 (RST), .A1 (nx6149), .A2 (nx8042)) ;
    or03 ix6327 (.Y (nx6326), .A0 (RST), .A1 (nx6156), .A2 (nx8246)) ;
    or03 ix6333 (.Y (nx6332), .A0 (RST), .A1 (nx6162), .A2 (nx8246)) ;
    or03 ix6339 (.Y (nx6338), .A0 (RST), .A1 (nx6168), .A2 (nx8246)) ;
    or03 ix6345 (.Y (nx6344), .A0 (RST), .A1 (nx6174), .A2 (nx8246)) ;
    or03 ix6351 (.Y (nx6350), .A0 (RST), .A1 (nx6180), .A2 (nx8246)) ;
    or03 ix6357 (.Y (nx6356), .A0 (RST), .A1 (nx6186), .A2 (nx8246)) ;
    or03 ix6363 (.Y (nx6362), .A0 (RST), .A1 (nx6192), .A2 (nx8246)) ;
    or03 ix6369 (.Y (nx6368), .A0 (RST), .A1 (nx6198), .A2 (nx8248)) ;
    or03 ix6375 (.Y (nx6374), .A0 (RST), .A1 (nx6204), .A2 (nx8248)) ;
    or03 ix6381 (.Y (nx6380), .A0 (RST), .A1 (nx6210), .A2 (nx8248)) ;
    or03 ix6387 (.Y (nx6386), .A0 (RST), .A1 (nx6216), .A2 (nx8248)) ;
    or03 ix6393 (.Y (nx6392), .A0 (RST), .A1 (nx6222), .A2 (nx8248)) ;
    or03 ix6399 (.Y (nx6398), .A0 (RST), .A1 (nx6228), .A2 (nx8248)) ;
    or03 ix6405 (.Y (nx6404), .A0 (RST), .A1 (nx6234), .A2 (nx8248)) ;
    or03 ix6411 (.Y (nx6410), .A0 (RST), .A1 (nx6240), .A2 (nx8250)) ;
    or03 ix6489 (.Y (nx6488), .A0 (RST), .A1 (nx6318), .A2 (nx8250)) ;
    or03 ix6495 (.Y (nx6494), .A0 (RST), .A1 (nx6324), .A2 (nx8250)) ;
    or03 ix6501 (.Y (nx6500), .A0 (RST), .A1 (nx6330), .A2 (nx8250)) ;
    or03 ix6507 (.Y (nx6506), .A0 (RST), .A1 (nx6336), .A2 (nx8250)) ;
    or03 ix6513 (.Y (nx6512), .A0 (RST), .A1 (nx6342), .A2 (nx8250)) ;
    or03 ix6519 (.Y (nx6518), .A0 (RST), .A1 (nx6348), .A2 (nx8250)) ;
    or03 ix6525 (.Y (nx6524), .A0 (RST), .A1 (nx6354), .A2 (nx8044)) ;
    or03 ix6531 (.Y (nx6530), .A0 (RST), .A1 (nx6360), .A2 (nx8044)) ;
    or03 ix6537 (.Y (nx6536), .A0 (RST), .A1 (nx6366), .A2 (nx8044)) ;
    or03 ix6543 (.Y (nx6542), .A0 (RST), .A1 (nx6372), .A2 (nx8044)) ;
    or03 ix6549 (.Y (nx6548), .A0 (RST), .A1 (nx6378), .A2 (nx8046)) ;
    or03 ix6555 (.Y (nx6554), .A0 (RST), .A1 (nx6384), .A2 (nx8046)) ;
    or03 ix6561 (.Y (nx6560), .A0 (RST), .A1 (nx6390), .A2 (nx8046)) ;
    or03 ix6567 (.Y (nx6566), .A0 (RST), .A1 (nx6396), .A2 (nx8046)) ;
    or03 ix6573 (.Y (nx6572), .A0 (RST), .A1 (nx6402), .A2 (nx8046)) ;
    or03 ix6579 (.Y (nx6578), .A0 (RST), .A1 (nx6408), .A2 (nx8046)) ;
    or03 ix6729 (.Y (nx6728), .A0 (RST), .A1 (nx6486), .A2 (nx8256)) ;
    or03 ix6735 (.Y (nx6734), .A0 (RST), .A1 (nx6492), .A2 (nx8256)) ;
    or03 ix6741 (.Y (nx6740), .A0 (RST), .A1 (nx6498), .A2 (nx8256)) ;
    or03 ix6747 (.Y (nx6746), .A0 (RST), .A1 (nx6504), .A2 (nx8256)) ;
    or03 ix6753 (.Y (nx6752), .A0 (RST), .A1 (nx6510), .A2 (nx8256)) ;
    or03 ix6759 (.Y (nx6758), .A0 (RST), .A1 (nx6516), .A2 (nx8256)) ;
    or03 ix6765 (.Y (nx6764), .A0 (RST), .A1 (nx6522), .A2 (nx8256)) ;
    or03 ix6771 (.Y (nx6770), .A0 (RST), .A1 (nx6528), .A2 (nx8258)) ;
    or03 ix6777 (.Y (nx6776), .A0 (RST), .A1 (nx6534), .A2 (nx8258)) ;
    or03 ix6783 (.Y (nx6782), .A0 (RST), .A1 (nx6540), .A2 (nx8258)) ;
    or03 ix6789 (.Y (nx6788), .A0 (RST), .A1 (nx6546), .A2 (nx8258)) ;
    or03 ix6795 (.Y (nx6794), .A0 (RST), .A1 (nx6552), .A2 (nx8258)) ;
    or03 ix6801 (.Y (nx6800), .A0 (RST), .A1 (nx6558), .A2 (nx8258)) ;
    or03 ix6807 (.Y (nx6806), .A0 (RST), .A1 (nx6564), .A2 (nx8258)) ;
    or03 ix6813 (.Y (nx6812), .A0 (RST), .A1 (nx6570), .A2 (nx8048)) ;
    or03 ix6819 (.Y (nx6818), .A0 (RST), .A1 (nx6576), .A2 (nx8048)) ;
    or03 ix6825 (.Y (nx6824), .A0 (RST), .A1 (nx6582), .A2 (nx8048)) ;
    or03 ix6831 (.Y (nx6830), .A0 (RST), .A1 (nx6588), .A2 (nx8048)) ;
    or03 ix6837 (.Y (nx6836), .A0 (RST), .A1 (nx6594), .A2 (nx8048)) ;
    or03 ix6843 (.Y (nx6842), .A0 (RST), .A1 (nx6600), .A2 (nx8260)) ;
    or03 ix6849 (.Y (nx6848), .A0 (RST), .A1 (nx6606), .A2 (nx8262)) ;
    or03 ix6855 (.Y (nx6854), .A0 (RST), .A1 (nx6612), .A2 (nx8262)) ;
    or03 ix6861 (.Y (nx6860), .A0 (RST), .A1 (nx6618), .A2 (nx8262)) ;
    or03 ix6867 (.Y (nx6866), .A0 (RST), .A1 (nx6624), .A2 (nx8262)) ;
    or03 ix6873 (.Y (nx6872), .A0 (RST), .A1 (nx6630), .A2 (nx8262)) ;
    or03 ix6879 (.Y (nx6878), .A0 (RST), .A1 (nx6636), .A2 (nx8262)) ;
    or03 ix6885 (.Y (nx6884), .A0 (RST), .A1 (nx6642), .A2 (nx8262)) ;
    or03 ix6891 (.Y (nx6890), .A0 (RST), .A1 (nx6648), .A2 (nx8264)) ;
    or03 ix6897 (.Y (nx6896), .A0 (RST), .A1 (nx6654), .A2 (nx8264)) ;
    or03 ix6903 (.Y (nx6902), .A0 (RST), .A1 (nx6660), .A2 (nx8264)) ;
    or03 ix6909 (.Y (nx6908), .A0 (RST), .A1 (nx6666), .A2 (nx8264)) ;
    or03 ix6915 (.Y (nx6914), .A0 (RST), .A1 (nx6672), .A2 (nx8264)) ;
    or03 ix6921 (.Y (nx6920), .A0 (RST), .A1 (nx6678), .A2 (nx8264)) ;
    or03 ix6927 (.Y (nx6926), .A0 (RST), .A1 (nx6684), .A2 (nx8264)) ;
    or03 ix6933 (.Y (nx6932), .A0 (RST), .A1 (nx6690), .A2 (nx8050)) ;
    or03 ix6939 (.Y (nx6938), .A0 (RST), .A1 (nx6696), .A2 (nx8050)) ;
    or03 ix6945 (.Y (nx6944), .A0 (RST), .A1 (nx6702), .A2 (nx8050)) ;
    or03 ix6951 (.Y (nx6950), .A0 (RST), .A1 (nx6708), .A2 (nx8050)) ;
    or03 ix6957 (.Y (nx6956), .A0 (RST), .A1 (nx6714), .A2 (nx8050)) ;
    or03 ix6963 (.Y (nx6962), .A0 (RST), .A1 (nx6720), .A2 (nx8050)) ;
    mux21_ni ix2062 (.Y (nx2061), .A0 (FilterDout_4__4__0), .A1 (nx86), .S0 (
             nx8292)) ;
    mux21_ni ix2072 (.Y (nx2071), .A0 (FilterDout_4__4__1), .A1 (nx96), .S0 (
             nx8292)) ;
    mux21_ni ix2082 (.Y (nx2081), .A0 (FilterDout_4__4__2), .A1 (nx106), .S0 (
             nx8242)) ;
    mux21_ni ix2092 (.Y (nx2091), .A0 (FilterDout_4__4__3), .A1 (nx116), .S0 (
             nx8242)) ;
    mux21_ni ix2102 (.Y (nx2101), .A0 (FilterDout_4__4__4), .A1 (nx126), .S0 (
             nx8242)) ;
    mux21_ni ix2112 (.Y (nx2111), .A0 (FilterDout_4__4__5), .A1 (nx136), .S0 (
             nx8242)) ;
    mux21_ni ix2122 (.Y (nx2121), .A0 (FilterDout_4__4__6), .A1 (nx146), .S0 (
             nx8242)) ;
    mux21_ni ix2132 (.Y (nx2131), .A0 (FilterDout_4__4__7), .A1 (nx156), .S0 (
             nx8242)) ;
    mux21_ni ix2222 (.Y (nx2221), .A0 (FilterDout_4__3__0), .A1 (nx218), .S0 (
             nx8242)) ;
    mux21_ni ix2232 (.Y (nx2231), .A0 (FilterDout_4__3__1), .A1 (nx228), .S0 (
             nx166)) ;
    mux21_ni ix2242 (.Y (nx2241), .A0 (FilterDout_4__3__2), .A1 (nx238), .S0 (
             nx166)) ;
    mux21_ni ix2252 (.Y (nx2251), .A0 (FilterDout_4__3__3), .A1 (nx248), .S0 (
             nx166)) ;
    mux21_ni ix2262 (.Y (nx2261), .A0 (FilterDout_4__3__4), .A1 (nx258), .S0 (
             nx166)) ;
    mux21_ni ix2272 (.Y (nx2271), .A0 (FilterDout_4__3__5), .A1 (nx268), .S0 (
             nx166)) ;
    mux21_ni ix2282 (.Y (nx2281), .A0 (FilterDout_4__3__6), .A1 (nx278), .S0 (
             nx166)) ;
    mux21_ni ix2292 (.Y (nx2291), .A0 (FilterDout_4__3__7), .A1 (nx288), .S0 (
             nx166)) ;
    or03 ix7262 (.Y (nx7261), .A0 (RST), .A1 (nx7090), .A2 (nx8186)) ;
    or03 ix7268 (.Y (nx7267), .A0 (RST), .A1 (nx7097), .A2 (nx8268)) ;
    or03 ix7274 (.Y (nx7273), .A0 (RST), .A1 (nx7103), .A2 (nx8268)) ;
    or03 ix7280 (.Y (nx7279), .A0 (RST), .A1 (nx7109), .A2 (nx8268)) ;
    or03 ix7286 (.Y (nx7285), .A0 (RST), .A1 (nx7115), .A2 (nx8268)) ;
    or03 ix7292 (.Y (nx7291), .A0 (RST), .A1 (nx7121), .A2 (nx8268)) ;
    or03 ix7298 (.Y (nx7297), .A0 (RST), .A1 (nx7127), .A2 (nx8268)) ;
    or03 ix7304 (.Y (nx7303), .A0 (RST), .A1 (nx7133), .A2 (nx8268)) ;
    or03 ix7310 (.Y (nx7309), .A0 (RST), .A1 (nx7139), .A2 (nx8270)) ;
    or03 ix7316 (.Y (nx7315), .A0 (RST), .A1 (nx7145), .A2 (nx8270)) ;
    or03 ix7322 (.Y (nx7321), .A0 (RST), .A1 (nx7151), .A2 (nx8270)) ;
    or03 ix7328 (.Y (nx7327), .A0 (RST), .A1 (nx7157), .A2 (nx8270)) ;
    or03 ix7334 (.Y (nx7333), .A0 (RST), .A1 (nx7163), .A2 (nx8270)) ;
    or03 ix7340 (.Y (nx7339), .A0 (RST), .A1 (nx7169), .A2 (nx8270)) ;
    or03 ix7346 (.Y (nx7345), .A0 (RST), .A1 (nx7175), .A2 (nx8270)) ;
    or03 ix7352 (.Y (nx7351), .A0 (RST), .A1 (nx7181), .A2 (nx8272)) ;
    or03 ix7430 (.Y (nx7429), .A0 (RST), .A1 (nx7259), .A2 (nx8272)) ;
    or03 ix7436 (.Y (nx7435), .A0 (RST), .A1 (nx7265), .A2 (nx8272)) ;
    or03 ix7442 (.Y (nx7441), .A0 (RST), .A1 (nx7271), .A2 (nx8272)) ;
    or03 ix7448 (.Y (nx7447), .A0 (RST), .A1 (nx7277), .A2 (nx8272)) ;
    or03 ix7454 (.Y (nx7453), .A0 (RST), .A1 (nx7283), .A2 (nx8272)) ;
    or03 ix7460 (.Y (nx7459), .A0 (RST), .A1 (nx7289), .A2 (nx8272)) ;
    or03 ix7466 (.Y (nx7465), .A0 (RST), .A1 (nx7295), .A2 (nx8188)) ;
    or03 ix7472 (.Y (nx7471), .A0 (RST), .A1 (nx7301), .A2 (nx8188)) ;
    or03 ix7478 (.Y (nx7477), .A0 (RST), .A1 (nx7307), .A2 (nx8188)) ;
    or03 ix7484 (.Y (nx7483), .A0 (RST), .A1 (nx7313), .A2 (nx8188)) ;
    or03 ix7490 (.Y (nx7489), .A0 (RST), .A1 (nx7319), .A2 (nx8190)) ;
    or03 ix7496 (.Y (nx7495), .A0 (RST), .A1 (nx7325), .A2 (nx8190)) ;
    or03 ix7502 (.Y (nx7501), .A0 (RST), .A1 (nx7331), .A2 (nx8190)) ;
    or03 ix7508 (.Y (nx7507), .A0 (RST), .A1 (nx7337), .A2 (nx8190)) ;
    or03 ix7514 (.Y (nx7513), .A0 (RST), .A1 (nx7343), .A2 (nx8190)) ;
    or03 ix7520 (.Y (nx7519), .A0 (RST), .A1 (nx7349), .A2 (nx8190)) ;
    or03 ix7670 (.Y (nx7669), .A0 (RST), .A1 (nx7427), .A2 (nx8278)) ;
    or03 ix7676 (.Y (nx7675), .A0 (RST), .A1 (nx7433), .A2 (nx8278)) ;
    or03 ix7682 (.Y (nx7681), .A0 (RST), .A1 (nx7439), .A2 (nx8278)) ;
    or03 ix7688 (.Y (nx7687), .A0 (RST), .A1 (nx7445), .A2 (nx8278)) ;
    or03 ix7694 (.Y (nx7693), .A0 (RST), .A1 (nx7451), .A2 (nx8278)) ;
    or03 ix7700 (.Y (nx7699), .A0 (RST), .A1 (nx7457), .A2 (nx8278)) ;
    or03 ix7706 (.Y (nx7705), .A0 (RST), .A1 (nx7463), .A2 (nx8278)) ;
    or03 ix7712 (.Y (nx7711), .A0 (RST), .A1 (nx7469), .A2 (nx8280)) ;
    or03 ix7718 (.Y (nx7717), .A0 (RST), .A1 (nx7475), .A2 (nx8280)) ;
    or03 ix7724 (.Y (nx7723), .A0 (RST), .A1 (nx7481), .A2 (nx8280)) ;
    or03 ix7730 (.Y (nx7729), .A0 (RST), .A1 (nx7487), .A2 (nx8280)) ;
    or03 ix7736 (.Y (nx7735), .A0 (RST), .A1 (nx7493), .A2 (nx8280)) ;
    or03 ix7742 (.Y (nx7741), .A0 (RST), .A1 (nx7499), .A2 (nx8280)) ;
    or03 ix7748 (.Y (nx7747), .A0 (RST), .A1 (nx7505), .A2 (nx8280)) ;
    or03 ix7754 (.Y (nx7753), .A0 (RST), .A1 (nx7511), .A2 (nx8192)) ;
    or03 ix7760 (.Y (nx7759), .A0 (RST), .A1 (nx7517), .A2 (nx8192)) ;
    or03 ix7766 (.Y (nx7765), .A0 (RST), .A1 (nx7523), .A2 (nx8192)) ;
    or03 ix7772 (.Y (nx7771), .A0 (RST), .A1 (nx7529), .A2 (nx8192)) ;
    or03 ix7778 (.Y (nx7777), .A0 (RST), .A1 (nx7535), .A2 (nx8192)) ;
    or03 ix7784 (.Y (nx7783), .A0 (RST), .A1 (nx7541), .A2 (nx8282)) ;
    or03 ix7790 (.Y (nx7789), .A0 (RST), .A1 (nx7547), .A2 (nx8284)) ;
    or03 ix7796 (.Y (nx7795), .A0 (RST), .A1 (nx7553), .A2 (nx8284)) ;
    or03 ix7802 (.Y (nx7801), .A0 (RST), .A1 (nx7559), .A2 (nx8284)) ;
    or03 ix7808 (.Y (nx7807), .A0 (RST), .A1 (nx7565), .A2 (nx8284)) ;
    or03 ix7814 (.Y (nx7813), .A0 (RST), .A1 (nx7571), .A2 (nx8284)) ;
    or03 ix7820 (.Y (nx7819), .A0 (RST), .A1 (nx7577), .A2 (nx8284)) ;
    or03 ix7826 (.Y (nx7825), .A0 (RST), .A1 (nx7583), .A2 (nx8284)) ;
    or03 ix7832 (.Y (nx7831), .A0 (RST), .A1 (nx7589), .A2 (nx8286)) ;
    or03 ix7838 (.Y (nx7837), .A0 (RST), .A1 (nx7595), .A2 (nx8286)) ;
    or03 ix7844 (.Y (nx7843), .A0 (RST), .A1 (nx7601), .A2 (nx8286)) ;
    or03 ix7850 (.Y (nx7849), .A0 (RST), .A1 (nx7607), .A2 (nx8286)) ;
    or03 ix7856 (.Y (nx7855), .A0 (RST), .A1 (nx7613), .A2 (nx8286)) ;
    or03 ix7862 (.Y (nx7861), .A0 (RST), .A1 (nx7619), .A2 (nx8286)) ;
    or03 ix7868 (.Y (nx7867), .A0 (RST), .A1 (nx7625), .A2 (nx8286)) ;
    or03 ix7874 (.Y (nx7873), .A0 (RST), .A1 (nx7631), .A2 (nx8194)) ;
    or03 ix7880 (.Y (nx7879), .A0 (RST), .A1 (nx7637), .A2 (nx8194)) ;
    or03 ix7886 (.Y (nx7885), .A0 (RST), .A1 (nx7643), .A2 (nx8194)) ;
    or03 ix7892 (.Y (nx7891), .A0 (RST), .A1 (nx7649), .A2 (nx8194)) ;
    or03 ix7898 (.Y (nx7897), .A0 (RST), .A1 (nx7655), .A2 (nx8194)) ;
    or03 ix7904 (.Y (nx7903), .A0 (RST), .A1 (nx7661), .A2 (nx8194)) ;
    inv02 ix8235 (.Y (nx8236), .A (nx8300)) ;
    inv02 ix8237 (.Y (nx8238), .A (nx8300)) ;
    inv02 ix8239 (.Y (nx8240), .A (nx8302)) ;
    inv02 ix8241 (.Y (nx8242), .A (nx8302)) ;
    inv02 ix8243 (.Y (nx8244), .A (nx8290)) ;
    inv02 ix8245 (.Y (nx8246), .A (nx8290)) ;
    inv02 ix8247 (.Y (nx8248), .A (nx8290)) ;
    inv02 ix8249 (.Y (nx8250), .A (nx8290)) ;
    inv02 ix8251 (.Y (nx8252), .A (nx8290)) ;
    inv02 ix8253 (.Y (nx8254), .A (nx8290)) ;
    inv02 ix8255 (.Y (nx8256), .A (nx8290)) ;
    inv02 ix8257 (.Y (nx8258), .A (nx8236)) ;
    inv02 ix8259 (.Y (nx8260), .A (nx8236)) ;
    inv02 ix8261 (.Y (nx8262), .A (nx8236)) ;
    inv02 ix8263 (.Y (nx8264), .A (nx8236)) ;
    inv02 ix8265 (.Y (nx8266), .A (nx8294)) ;
    inv02 ix8267 (.Y (nx8268), .A (nx8294)) ;
    inv02 ix8269 (.Y (nx8270), .A (nx8294)) ;
    inv02 ix8271 (.Y (nx8272), .A (nx8294)) ;
    inv02 ix8273 (.Y (nx8274), .A (nx8294)) ;
    inv02 ix8275 (.Y (nx8276), .A (nx8294)) ;
    inv02 ix8277 (.Y (nx8278), .A (nx8294)) ;
    inv02 ix8279 (.Y (nx8280), .A (nx8240)) ;
    inv02 ix8281 (.Y (nx8282), .A (nx8240)) ;
    inv02 ix8283 (.Y (nx8284), .A (nx8240)) ;
    inv02 ix8285 (.Y (nx8286), .A (nx8240)) ;
    inv02 ix8287 (.Y (nx8288), .A (nx8300)) ;
    inv02 ix8289 (.Y (nx8290), .A (nx8300)) ;
    inv02 ix8291 (.Y (nx8292), .A (nx8302)) ;
    inv02 ix8293 (.Y (nx8294), .A (nx8302)) ;
    inv01 ix8299 (.Y (nx8300), .A (nx82)) ;
    inv01 ix8301 (.Y (nx8302), .A (nx166)) ;
endmodule


module RAM_8_18 ( CLK, WR, Address, Din, Dout ) ;

    input CLK ;
    input WR ;
    input [17:0]Address ;
    input [7:0]Din ;
    output [39:0]Dout ;




endmodule


module accelerator ( CLK, RST, Start, FilterSize, Instr, FilterDin_0__0__7, 
                     FilterDin_0__0__6, FilterDin_0__0__5, FilterDin_0__0__4, 
                     FilterDin_0__0__3, FilterDin_0__0__2, FilterDin_0__0__1, 
                     FilterDin_0__0__0, FilterDin_0__1__7, FilterDin_0__1__6, 
                     FilterDin_0__1__5, FilterDin_0__1__4, FilterDin_0__1__3, 
                     FilterDin_0__1__2, FilterDin_0__1__1, FilterDin_0__1__0, 
                     FilterDin_0__2__7, FilterDin_0__2__6, FilterDin_0__2__5, 
                     FilterDin_0__2__4, FilterDin_0__2__3, FilterDin_0__2__2, 
                     FilterDin_0__2__1, FilterDin_0__2__0, FilterDin_0__3__7, 
                     FilterDin_0__3__6, FilterDin_0__3__5, FilterDin_0__3__4, 
                     FilterDin_0__3__3, FilterDin_0__3__2, FilterDin_0__3__1, 
                     FilterDin_0__3__0, FilterDin_0__4__7, FilterDin_0__4__6, 
                     FilterDin_0__4__5, FilterDin_0__4__4, FilterDin_0__4__3, 
                     FilterDin_0__4__2, FilterDin_0__4__1, FilterDin_0__4__0, 
                     FilterDin_1__0__7, FilterDin_1__0__6, FilterDin_1__0__5, 
                     FilterDin_1__0__4, FilterDin_1__0__3, FilterDin_1__0__2, 
                     FilterDin_1__0__1, FilterDin_1__0__0, FilterDin_1__1__7, 
                     FilterDin_1__1__6, FilterDin_1__1__5, FilterDin_1__1__4, 
                     FilterDin_1__1__3, FilterDin_1__1__2, FilterDin_1__1__1, 
                     FilterDin_1__1__0, FilterDin_1__2__7, FilterDin_1__2__6, 
                     FilterDin_1__2__5, FilterDin_1__2__4, FilterDin_1__2__3, 
                     FilterDin_1__2__2, FilterDin_1__2__1, FilterDin_1__2__0, 
                     FilterDin_1__3__7, FilterDin_1__3__6, FilterDin_1__3__5, 
                     FilterDin_1__3__4, FilterDin_1__3__3, FilterDin_1__3__2, 
                     FilterDin_1__3__1, FilterDin_1__3__0, FilterDin_1__4__7, 
                     FilterDin_1__4__6, FilterDin_1__4__5, FilterDin_1__4__4, 
                     FilterDin_1__4__3, FilterDin_1__4__2, FilterDin_1__4__1, 
                     FilterDin_1__4__0, FilterDin_2__0__7, FilterDin_2__0__6, 
                     FilterDin_2__0__5, FilterDin_2__0__4, FilterDin_2__0__3, 
                     FilterDin_2__0__2, FilterDin_2__0__1, FilterDin_2__0__0, 
                     FilterDin_2__1__7, FilterDin_2__1__6, FilterDin_2__1__5, 
                     FilterDin_2__1__4, FilterDin_2__1__3, FilterDin_2__1__2, 
                     FilterDin_2__1__1, FilterDin_2__1__0, FilterDin_2__2__7, 
                     FilterDin_2__2__6, FilterDin_2__2__5, FilterDin_2__2__4, 
                     FilterDin_2__2__3, FilterDin_2__2__2, FilterDin_2__2__1, 
                     FilterDin_2__2__0, FilterDin_2__3__7, FilterDin_2__3__6, 
                     FilterDin_2__3__5, FilterDin_2__3__4, FilterDin_2__3__3, 
                     FilterDin_2__3__2, FilterDin_2__3__1, FilterDin_2__3__0, 
                     FilterDin_2__4__7, FilterDin_2__4__6, FilterDin_2__4__5, 
                     FilterDin_2__4__4, FilterDin_2__4__3, FilterDin_2__4__2, 
                     FilterDin_2__4__1, FilterDin_2__4__0, FilterDin_3__0__7, 
                     FilterDin_3__0__6, FilterDin_3__0__5, FilterDin_3__0__4, 
                     FilterDin_3__0__3, FilterDin_3__0__2, FilterDin_3__0__1, 
                     FilterDin_3__0__0, FilterDin_3__1__7, FilterDin_3__1__6, 
                     FilterDin_3__1__5, FilterDin_3__1__4, FilterDin_3__1__3, 
                     FilterDin_3__1__2, FilterDin_3__1__1, FilterDin_3__1__0, 
                     FilterDin_3__2__7, FilterDin_3__2__6, FilterDin_3__2__5, 
                     FilterDin_3__2__4, FilterDin_3__2__3, FilterDin_3__2__2, 
                     FilterDin_3__2__1, FilterDin_3__2__0, FilterDin_3__3__7, 
                     FilterDin_3__3__6, FilterDin_3__3__5, FilterDin_3__3__4, 
                     FilterDin_3__3__3, FilterDin_3__3__2, FilterDin_3__3__1, 
                     FilterDin_3__3__0, FilterDin_3__4__7, FilterDin_3__4__6, 
                     FilterDin_3__4__5, FilterDin_3__4__4, FilterDin_3__4__3, 
                     FilterDin_3__4__2, FilterDin_3__4__1, FilterDin_3__4__0, 
                     FilterDin_4__0__7, FilterDin_4__0__6, FilterDin_4__0__5, 
                     FilterDin_4__0__4, FilterDin_4__0__3, FilterDin_4__0__2, 
                     FilterDin_4__0__1, FilterDin_4__0__0, FilterDin_4__1__7, 
                     FilterDin_4__1__6, FilterDin_4__1__5, FilterDin_4__1__4, 
                     FilterDin_4__1__3, FilterDin_4__1__2, FilterDin_4__1__1, 
                     FilterDin_4__1__0, FilterDin_4__2__7, FilterDin_4__2__6, 
                     FilterDin_4__2__5, FilterDin_4__2__4, FilterDin_4__2__3, 
                     FilterDin_4__2__2, FilterDin_4__2__1, FilterDin_4__2__0, 
                     FilterDin_4__3__7, FilterDin_4__3__6, FilterDin_4__3__5, 
                     FilterDin_4__3__4, FilterDin_4__3__3, FilterDin_4__3__2, 
                     FilterDin_4__3__1, FilterDin_4__3__0, FilterDin_4__4__7, 
                     FilterDin_4__4__6, FilterDin_4__4__5, FilterDin_4__4__4, 
                     FilterDin_4__4__3, FilterDin_4__4__2, FilterDin_4__4__1, 
                     FilterDin_4__4__0, WindowDin_0__0__7, WindowDin_0__0__6, 
                     WindowDin_0__0__5, WindowDin_0__0__4, WindowDin_0__0__3, 
                     WindowDin_0__0__2, WindowDin_0__0__1, WindowDin_0__0__0, 
                     WindowDin_0__1__7, WindowDin_0__1__6, WindowDin_0__1__5, 
                     WindowDin_0__1__4, WindowDin_0__1__3, WindowDin_0__1__2, 
                     WindowDin_0__1__1, WindowDin_0__1__0, WindowDin_0__2__7, 
                     WindowDin_0__2__6, WindowDin_0__2__5, WindowDin_0__2__4, 
                     WindowDin_0__2__3, WindowDin_0__2__2, WindowDin_0__2__1, 
                     WindowDin_0__2__0, WindowDin_0__3__7, WindowDin_0__3__6, 
                     WindowDin_0__3__5, WindowDin_0__3__4, WindowDin_0__3__3, 
                     WindowDin_0__3__2, WindowDin_0__3__1, WindowDin_0__3__0, 
                     WindowDin_0__4__7, WindowDin_0__4__6, WindowDin_0__4__5, 
                     WindowDin_0__4__4, WindowDin_0__4__3, WindowDin_0__4__2, 
                     WindowDin_0__4__1, WindowDin_0__4__0, WindowDin_1__0__7, 
                     WindowDin_1__0__6, WindowDin_1__0__5, WindowDin_1__0__4, 
                     WindowDin_1__0__3, WindowDin_1__0__2, WindowDin_1__0__1, 
                     WindowDin_1__0__0, WindowDin_1__1__7, WindowDin_1__1__6, 
                     WindowDin_1__1__5, WindowDin_1__1__4, WindowDin_1__1__3, 
                     WindowDin_1__1__2, WindowDin_1__1__1, WindowDin_1__1__0, 
                     WindowDin_1__2__7, WindowDin_1__2__6, WindowDin_1__2__5, 
                     WindowDin_1__2__4, WindowDin_1__2__3, WindowDin_1__2__2, 
                     WindowDin_1__2__1, WindowDin_1__2__0, WindowDin_1__3__7, 
                     WindowDin_1__3__6, WindowDin_1__3__5, WindowDin_1__3__4, 
                     WindowDin_1__3__3, WindowDin_1__3__2, WindowDin_1__3__1, 
                     WindowDin_1__3__0, WindowDin_1__4__7, WindowDin_1__4__6, 
                     WindowDin_1__4__5, WindowDin_1__4__4, WindowDin_1__4__3, 
                     WindowDin_1__4__2, WindowDin_1__4__1, WindowDin_1__4__0, 
                     WindowDin_2__0__7, WindowDin_2__0__6, WindowDin_2__0__5, 
                     WindowDin_2__0__4, WindowDin_2__0__3, WindowDin_2__0__2, 
                     WindowDin_2__0__1, WindowDin_2__0__0, WindowDin_2__1__7, 
                     WindowDin_2__1__6, WindowDin_2__1__5, WindowDin_2__1__4, 
                     WindowDin_2__1__3, WindowDin_2__1__2, WindowDin_2__1__1, 
                     WindowDin_2__1__0, WindowDin_2__2__7, WindowDin_2__2__6, 
                     WindowDin_2__2__5, WindowDin_2__2__4, WindowDin_2__2__3, 
                     WindowDin_2__2__2, WindowDin_2__2__1, WindowDin_2__2__0, 
                     WindowDin_2__3__7, WindowDin_2__3__6, WindowDin_2__3__5, 
                     WindowDin_2__3__4, WindowDin_2__3__3, WindowDin_2__3__2, 
                     WindowDin_2__3__1, WindowDin_2__3__0, WindowDin_2__4__7, 
                     WindowDin_2__4__6, WindowDin_2__4__5, WindowDin_2__4__4, 
                     WindowDin_2__4__3, WindowDin_2__4__2, WindowDin_2__4__1, 
                     WindowDin_2__4__0, WindowDin_3__0__7, WindowDin_3__0__6, 
                     WindowDin_3__0__5, WindowDin_3__0__4, WindowDin_3__0__3, 
                     WindowDin_3__0__2, WindowDin_3__0__1, WindowDin_3__0__0, 
                     WindowDin_3__1__7, WindowDin_3__1__6, WindowDin_3__1__5, 
                     WindowDin_3__1__4, WindowDin_3__1__3, WindowDin_3__1__2, 
                     WindowDin_3__1__1, WindowDin_3__1__0, WindowDin_3__2__7, 
                     WindowDin_3__2__6, WindowDin_3__2__5, WindowDin_3__2__4, 
                     WindowDin_3__2__3, WindowDin_3__2__2, WindowDin_3__2__1, 
                     WindowDin_3__2__0, WindowDin_3__3__7, WindowDin_3__3__6, 
                     WindowDin_3__3__5, WindowDin_3__3__4, WindowDin_3__3__3, 
                     WindowDin_3__3__2, WindowDin_3__3__1, WindowDin_3__3__0, 
                     WindowDin_3__4__7, WindowDin_3__4__6, WindowDin_3__4__5, 
                     WindowDin_3__4__4, WindowDin_3__4__3, WindowDin_3__4__2, 
                     WindowDin_3__4__1, WindowDin_3__4__0, WindowDin_4__0__7, 
                     WindowDin_4__0__6, WindowDin_4__0__5, WindowDin_4__0__4, 
                     WindowDin_4__0__3, WindowDin_4__0__2, WindowDin_4__0__1, 
                     WindowDin_4__0__0, WindowDin_4__1__7, WindowDin_4__1__6, 
                     WindowDin_4__1__5, WindowDin_4__1__4, WindowDin_4__1__3, 
                     WindowDin_4__1__2, WindowDin_4__1__1, WindowDin_4__1__0, 
                     WindowDin_4__2__7, WindowDin_4__2__6, WindowDin_4__2__5, 
                     WindowDin_4__2__4, WindowDin_4__2__3, WindowDin_4__2__2, 
                     WindowDin_4__2__1, WindowDin_4__2__0, WindowDin_4__3__7, 
                     WindowDin_4__3__6, WindowDin_4__3__5, WindowDin_4__3__4, 
                     WindowDin_4__3__3, WindowDin_4__3__2, WindowDin_4__3__1, 
                     WindowDin_4__3__0, WindowDin_4__4__7, WindowDin_4__4__6, 
                     WindowDin_4__4__5, WindowDin_4__4__4, WindowDin_4__4__3, 
                     WindowDin_4__4__2, WindowDin_4__4__1, WindowDin_4__4__0, 
                     Done, Result ) ;

    input CLK ;
    input RST ;
    input Start ;
    input FilterSize ;
    input Instr ;
    input FilterDin_0__0__7 ;
    input FilterDin_0__0__6 ;
    input FilterDin_0__0__5 ;
    input FilterDin_0__0__4 ;
    input FilterDin_0__0__3 ;
    input FilterDin_0__0__2 ;
    input FilterDin_0__0__1 ;
    input FilterDin_0__0__0 ;
    input FilterDin_0__1__7 ;
    input FilterDin_0__1__6 ;
    input FilterDin_0__1__5 ;
    input FilterDin_0__1__4 ;
    input FilterDin_0__1__3 ;
    input FilterDin_0__1__2 ;
    input FilterDin_0__1__1 ;
    input FilterDin_0__1__0 ;
    input FilterDin_0__2__7 ;
    input FilterDin_0__2__6 ;
    input FilterDin_0__2__5 ;
    input FilterDin_0__2__4 ;
    input FilterDin_0__2__3 ;
    input FilterDin_0__2__2 ;
    input FilterDin_0__2__1 ;
    input FilterDin_0__2__0 ;
    input FilterDin_0__3__7 ;
    input FilterDin_0__3__6 ;
    input FilterDin_0__3__5 ;
    input FilterDin_0__3__4 ;
    input FilterDin_0__3__3 ;
    input FilterDin_0__3__2 ;
    input FilterDin_0__3__1 ;
    input FilterDin_0__3__0 ;
    input FilterDin_0__4__7 ;
    input FilterDin_0__4__6 ;
    input FilterDin_0__4__5 ;
    input FilterDin_0__4__4 ;
    input FilterDin_0__4__3 ;
    input FilterDin_0__4__2 ;
    input FilterDin_0__4__1 ;
    input FilterDin_0__4__0 ;
    input FilterDin_1__0__7 ;
    input FilterDin_1__0__6 ;
    input FilterDin_1__0__5 ;
    input FilterDin_1__0__4 ;
    input FilterDin_1__0__3 ;
    input FilterDin_1__0__2 ;
    input FilterDin_1__0__1 ;
    input FilterDin_1__0__0 ;
    input FilterDin_1__1__7 ;
    input FilterDin_1__1__6 ;
    input FilterDin_1__1__5 ;
    input FilterDin_1__1__4 ;
    input FilterDin_1__1__3 ;
    input FilterDin_1__1__2 ;
    input FilterDin_1__1__1 ;
    input FilterDin_1__1__0 ;
    input FilterDin_1__2__7 ;
    input FilterDin_1__2__6 ;
    input FilterDin_1__2__5 ;
    input FilterDin_1__2__4 ;
    input FilterDin_1__2__3 ;
    input FilterDin_1__2__2 ;
    input FilterDin_1__2__1 ;
    input FilterDin_1__2__0 ;
    input FilterDin_1__3__7 ;
    input FilterDin_1__3__6 ;
    input FilterDin_1__3__5 ;
    input FilterDin_1__3__4 ;
    input FilterDin_1__3__3 ;
    input FilterDin_1__3__2 ;
    input FilterDin_1__3__1 ;
    input FilterDin_1__3__0 ;
    input FilterDin_1__4__7 ;
    input FilterDin_1__4__6 ;
    input FilterDin_1__4__5 ;
    input FilterDin_1__4__4 ;
    input FilterDin_1__4__3 ;
    input FilterDin_1__4__2 ;
    input FilterDin_1__4__1 ;
    input FilterDin_1__4__0 ;
    input FilterDin_2__0__7 ;
    input FilterDin_2__0__6 ;
    input FilterDin_2__0__5 ;
    input FilterDin_2__0__4 ;
    input FilterDin_2__0__3 ;
    input FilterDin_2__0__2 ;
    input FilterDin_2__0__1 ;
    input FilterDin_2__0__0 ;
    input FilterDin_2__1__7 ;
    input FilterDin_2__1__6 ;
    input FilterDin_2__1__5 ;
    input FilterDin_2__1__4 ;
    input FilterDin_2__1__3 ;
    input FilterDin_2__1__2 ;
    input FilterDin_2__1__1 ;
    input FilterDin_2__1__0 ;
    input FilterDin_2__2__7 ;
    input FilterDin_2__2__6 ;
    input FilterDin_2__2__5 ;
    input FilterDin_2__2__4 ;
    input FilterDin_2__2__3 ;
    input FilterDin_2__2__2 ;
    input FilterDin_2__2__1 ;
    input FilterDin_2__2__0 ;
    input FilterDin_2__3__7 ;
    input FilterDin_2__3__6 ;
    input FilterDin_2__3__5 ;
    input FilterDin_2__3__4 ;
    input FilterDin_2__3__3 ;
    input FilterDin_2__3__2 ;
    input FilterDin_2__3__1 ;
    input FilterDin_2__3__0 ;
    input FilterDin_2__4__7 ;
    input FilterDin_2__4__6 ;
    input FilterDin_2__4__5 ;
    input FilterDin_2__4__4 ;
    input FilterDin_2__4__3 ;
    input FilterDin_2__4__2 ;
    input FilterDin_2__4__1 ;
    input FilterDin_2__4__0 ;
    input FilterDin_3__0__7 ;
    input FilterDin_3__0__6 ;
    input FilterDin_3__0__5 ;
    input FilterDin_3__0__4 ;
    input FilterDin_3__0__3 ;
    input FilterDin_3__0__2 ;
    input FilterDin_3__0__1 ;
    input FilterDin_3__0__0 ;
    input FilterDin_3__1__7 ;
    input FilterDin_3__1__6 ;
    input FilterDin_3__1__5 ;
    input FilterDin_3__1__4 ;
    input FilterDin_3__1__3 ;
    input FilterDin_3__1__2 ;
    input FilterDin_3__1__1 ;
    input FilterDin_3__1__0 ;
    input FilterDin_3__2__7 ;
    input FilterDin_3__2__6 ;
    input FilterDin_3__2__5 ;
    input FilterDin_3__2__4 ;
    input FilterDin_3__2__3 ;
    input FilterDin_3__2__2 ;
    input FilterDin_3__2__1 ;
    input FilterDin_3__2__0 ;
    input FilterDin_3__3__7 ;
    input FilterDin_3__3__6 ;
    input FilterDin_3__3__5 ;
    input FilterDin_3__3__4 ;
    input FilterDin_3__3__3 ;
    input FilterDin_3__3__2 ;
    input FilterDin_3__3__1 ;
    input FilterDin_3__3__0 ;
    input FilterDin_3__4__7 ;
    input FilterDin_3__4__6 ;
    input FilterDin_3__4__5 ;
    input FilterDin_3__4__4 ;
    input FilterDin_3__4__3 ;
    input FilterDin_3__4__2 ;
    input FilterDin_3__4__1 ;
    input FilterDin_3__4__0 ;
    input FilterDin_4__0__7 ;
    input FilterDin_4__0__6 ;
    input FilterDin_4__0__5 ;
    input FilterDin_4__0__4 ;
    input FilterDin_4__0__3 ;
    input FilterDin_4__0__2 ;
    input FilterDin_4__0__1 ;
    input FilterDin_4__0__0 ;
    input FilterDin_4__1__7 ;
    input FilterDin_4__1__6 ;
    input FilterDin_4__1__5 ;
    input FilterDin_4__1__4 ;
    input FilterDin_4__1__3 ;
    input FilterDin_4__1__2 ;
    input FilterDin_4__1__1 ;
    input FilterDin_4__1__0 ;
    input FilterDin_4__2__7 ;
    input FilterDin_4__2__6 ;
    input FilterDin_4__2__5 ;
    input FilterDin_4__2__4 ;
    input FilterDin_4__2__3 ;
    input FilterDin_4__2__2 ;
    input FilterDin_4__2__1 ;
    input FilterDin_4__2__0 ;
    input FilterDin_4__3__7 ;
    input FilterDin_4__3__6 ;
    input FilterDin_4__3__5 ;
    input FilterDin_4__3__4 ;
    input FilterDin_4__3__3 ;
    input FilterDin_4__3__2 ;
    input FilterDin_4__3__1 ;
    input FilterDin_4__3__0 ;
    input FilterDin_4__4__7 ;
    input FilterDin_4__4__6 ;
    input FilterDin_4__4__5 ;
    input FilterDin_4__4__4 ;
    input FilterDin_4__4__3 ;
    input FilterDin_4__4__2 ;
    input FilterDin_4__4__1 ;
    input FilterDin_4__4__0 ;
    input WindowDin_0__0__7 ;
    input WindowDin_0__0__6 ;
    input WindowDin_0__0__5 ;
    input WindowDin_0__0__4 ;
    input WindowDin_0__0__3 ;
    input WindowDin_0__0__2 ;
    input WindowDin_0__0__1 ;
    input WindowDin_0__0__0 ;
    input WindowDin_0__1__7 ;
    input WindowDin_0__1__6 ;
    input WindowDin_0__1__5 ;
    input WindowDin_0__1__4 ;
    input WindowDin_0__1__3 ;
    input WindowDin_0__1__2 ;
    input WindowDin_0__1__1 ;
    input WindowDin_0__1__0 ;
    input WindowDin_0__2__7 ;
    input WindowDin_0__2__6 ;
    input WindowDin_0__2__5 ;
    input WindowDin_0__2__4 ;
    input WindowDin_0__2__3 ;
    input WindowDin_0__2__2 ;
    input WindowDin_0__2__1 ;
    input WindowDin_0__2__0 ;
    input WindowDin_0__3__7 ;
    input WindowDin_0__3__6 ;
    input WindowDin_0__3__5 ;
    input WindowDin_0__3__4 ;
    input WindowDin_0__3__3 ;
    input WindowDin_0__3__2 ;
    input WindowDin_0__3__1 ;
    input WindowDin_0__3__0 ;
    input WindowDin_0__4__7 ;
    input WindowDin_0__4__6 ;
    input WindowDin_0__4__5 ;
    input WindowDin_0__4__4 ;
    input WindowDin_0__4__3 ;
    input WindowDin_0__4__2 ;
    input WindowDin_0__4__1 ;
    input WindowDin_0__4__0 ;
    input WindowDin_1__0__7 ;
    input WindowDin_1__0__6 ;
    input WindowDin_1__0__5 ;
    input WindowDin_1__0__4 ;
    input WindowDin_1__0__3 ;
    input WindowDin_1__0__2 ;
    input WindowDin_1__0__1 ;
    input WindowDin_1__0__0 ;
    input WindowDin_1__1__7 ;
    input WindowDin_1__1__6 ;
    input WindowDin_1__1__5 ;
    input WindowDin_1__1__4 ;
    input WindowDin_1__1__3 ;
    input WindowDin_1__1__2 ;
    input WindowDin_1__1__1 ;
    input WindowDin_1__1__0 ;
    input WindowDin_1__2__7 ;
    input WindowDin_1__2__6 ;
    input WindowDin_1__2__5 ;
    input WindowDin_1__2__4 ;
    input WindowDin_1__2__3 ;
    input WindowDin_1__2__2 ;
    input WindowDin_1__2__1 ;
    input WindowDin_1__2__0 ;
    input WindowDin_1__3__7 ;
    input WindowDin_1__3__6 ;
    input WindowDin_1__3__5 ;
    input WindowDin_1__3__4 ;
    input WindowDin_1__3__3 ;
    input WindowDin_1__3__2 ;
    input WindowDin_1__3__1 ;
    input WindowDin_1__3__0 ;
    input WindowDin_1__4__7 ;
    input WindowDin_1__4__6 ;
    input WindowDin_1__4__5 ;
    input WindowDin_1__4__4 ;
    input WindowDin_1__4__3 ;
    input WindowDin_1__4__2 ;
    input WindowDin_1__4__1 ;
    input WindowDin_1__4__0 ;
    input WindowDin_2__0__7 ;
    input WindowDin_2__0__6 ;
    input WindowDin_2__0__5 ;
    input WindowDin_2__0__4 ;
    input WindowDin_2__0__3 ;
    input WindowDin_2__0__2 ;
    input WindowDin_2__0__1 ;
    input WindowDin_2__0__0 ;
    input WindowDin_2__1__7 ;
    input WindowDin_2__1__6 ;
    input WindowDin_2__1__5 ;
    input WindowDin_2__1__4 ;
    input WindowDin_2__1__3 ;
    input WindowDin_2__1__2 ;
    input WindowDin_2__1__1 ;
    input WindowDin_2__1__0 ;
    input WindowDin_2__2__7 ;
    input WindowDin_2__2__6 ;
    input WindowDin_2__2__5 ;
    input WindowDin_2__2__4 ;
    input WindowDin_2__2__3 ;
    input WindowDin_2__2__2 ;
    input WindowDin_2__2__1 ;
    input WindowDin_2__2__0 ;
    input WindowDin_2__3__7 ;
    input WindowDin_2__3__6 ;
    input WindowDin_2__3__5 ;
    input WindowDin_2__3__4 ;
    input WindowDin_2__3__3 ;
    input WindowDin_2__3__2 ;
    input WindowDin_2__3__1 ;
    input WindowDin_2__3__0 ;
    input WindowDin_2__4__7 ;
    input WindowDin_2__4__6 ;
    input WindowDin_2__4__5 ;
    input WindowDin_2__4__4 ;
    input WindowDin_2__4__3 ;
    input WindowDin_2__4__2 ;
    input WindowDin_2__4__1 ;
    input WindowDin_2__4__0 ;
    input WindowDin_3__0__7 ;
    input WindowDin_3__0__6 ;
    input WindowDin_3__0__5 ;
    input WindowDin_3__0__4 ;
    input WindowDin_3__0__3 ;
    input WindowDin_3__0__2 ;
    input WindowDin_3__0__1 ;
    input WindowDin_3__0__0 ;
    input WindowDin_3__1__7 ;
    input WindowDin_3__1__6 ;
    input WindowDin_3__1__5 ;
    input WindowDin_3__1__4 ;
    input WindowDin_3__1__3 ;
    input WindowDin_3__1__2 ;
    input WindowDin_3__1__1 ;
    input WindowDin_3__1__0 ;
    input WindowDin_3__2__7 ;
    input WindowDin_3__2__6 ;
    input WindowDin_3__2__5 ;
    input WindowDin_3__2__4 ;
    input WindowDin_3__2__3 ;
    input WindowDin_3__2__2 ;
    input WindowDin_3__2__1 ;
    input WindowDin_3__2__0 ;
    input WindowDin_3__3__7 ;
    input WindowDin_3__3__6 ;
    input WindowDin_3__3__5 ;
    input WindowDin_3__3__4 ;
    input WindowDin_3__3__3 ;
    input WindowDin_3__3__2 ;
    input WindowDin_3__3__1 ;
    input WindowDin_3__3__0 ;
    input WindowDin_3__4__7 ;
    input WindowDin_3__4__6 ;
    input WindowDin_3__4__5 ;
    input WindowDin_3__4__4 ;
    input WindowDin_3__4__3 ;
    input WindowDin_3__4__2 ;
    input WindowDin_3__4__1 ;
    input WindowDin_3__4__0 ;
    input WindowDin_4__0__7 ;
    input WindowDin_4__0__6 ;
    input WindowDin_4__0__5 ;
    input WindowDin_4__0__4 ;
    input WindowDin_4__0__3 ;
    input WindowDin_4__0__2 ;
    input WindowDin_4__0__1 ;
    input WindowDin_4__0__0 ;
    input WindowDin_4__1__7 ;
    input WindowDin_4__1__6 ;
    input WindowDin_4__1__5 ;
    input WindowDin_4__1__4 ;
    input WindowDin_4__1__3 ;
    input WindowDin_4__1__2 ;
    input WindowDin_4__1__1 ;
    input WindowDin_4__1__0 ;
    input WindowDin_4__2__7 ;
    input WindowDin_4__2__6 ;
    input WindowDin_4__2__5 ;
    input WindowDin_4__2__4 ;
    input WindowDin_4__2__3 ;
    input WindowDin_4__2__2 ;
    input WindowDin_4__2__1 ;
    input WindowDin_4__2__0 ;
    input WindowDin_4__3__7 ;
    input WindowDin_4__3__6 ;
    input WindowDin_4__3__5 ;
    input WindowDin_4__3__4 ;
    input WindowDin_4__3__3 ;
    input WindowDin_4__3__2 ;
    input WindowDin_4__3__1 ;
    input WindowDin_4__3__0 ;
    input WindowDin_4__4__7 ;
    input WindowDin_4__4__6 ;
    input WindowDin_4__4__5 ;
    input WindowDin_4__4__4 ;
    input WindowDin_4__4__3 ;
    input WindowDin_4__4__2 ;
    input WindowDin_4__4__1 ;
    input WindowDin_4__4__0 ;
    output Done ;
    output [7:0]Result ;

    wire LoopingAndResultNotReady, L1FirstOperands_0__15, L1FirstOperands_0__14, 
         L1FirstOperands_0__13, L1FirstOperands_0__12, L1FirstOperands_0__11, 
         L1FirstOperands_0__10, L1FirstOperands_0__9, L1FirstOperands_0__8, 
         L1FirstOperands_0__7, L1FirstOperands_0__6, L1FirstOperands_0__5, 
         L1FirstOperands_0__4, L1FirstOperands_0__3, L1FirstOperands_0__2, 
         L1FirstOperands_0__1, L1FirstOperands_0__0, L1FirstOperands_2__15, 
         L1FirstOperands_2__14, L1FirstOperands_2__13, L1FirstOperands_2__12, 
         L1FirstOperands_2__11, L1FirstOperands_2__10, L1FirstOperands_2__9, 
         L1FirstOperands_2__8, L1FirstOperands_2__7, L1FirstOperands_2__6, 
         L1FirstOperands_2__5, L1FirstOperands_2__4, L1FirstOperands_2__3, 
         L1FirstOperands_2__2, L1FirstOperands_2__1, L1FirstOperands_2__0, 
         L1FirstOperands_3__15, L1FirstOperands_3__14, L1FirstOperands_3__13, 
         L1FirstOperands_3__12, L1FirstOperands_3__11, L1FirstOperands_3__10, 
         L1FirstOperands_3__9, L1FirstOperands_3__8, L1FirstOperands_3__7, 
         L1FirstOperands_3__6, L1FirstOperands_3__5, L1FirstOperands_3__4, 
         L1FirstOperands_3__3, L1FirstOperands_3__2, L1FirstOperands_3__1, 
         L1FirstOperands_3__0, L1FirstOperands_4__15, L1FirstOperands_4__14, 
         L1FirstOperands_4__13, L1FirstOperands_4__12, L1FirstOperands_4__11, 
         L1FirstOperands_4__10, L1FirstOperands_4__9, L1FirstOperands_4__8, 
         L1FirstOperands_4__7, L1FirstOperands_4__6, L1FirstOperands_4__5, 
         L1FirstOperands_4__4, L1FirstOperands_4__3, L1FirstOperands_4__2, 
         L1FirstOperands_4__1, L1FirstOperands_4__0, L1FirstOperands_6__15, 
         L1FirstOperands_6__14, L1FirstOperands_6__13, L1FirstOperands_6__12, 
         L1FirstOperands_6__11, L1FirstOperands_6__10, L1FirstOperands_6__9, 
         L1FirstOperands_6__8, L1FirstOperands_6__7, L1FirstOperands_6__6, 
         L1FirstOperands_6__5, L1FirstOperands_6__4, L1FirstOperands_6__3, 
         L1FirstOperands_6__2, L1FirstOperands_6__1, L1FirstOperands_6__0, 
         L1FirstOperands_7__15, L1FirstOperands_7__14, L1FirstOperands_7__13, 
         L1FirstOperands_7__12, L1FirstOperands_7__11, L1FirstOperands_7__10, 
         L1FirstOperands_7__9, L1FirstOperands_7__8, L1FirstOperands_7__7, 
         L1FirstOperands_7__6, L1FirstOperands_7__5, L1FirstOperands_7__4, 
         L1FirstOperands_7__3, L1FirstOperands_7__2, L1FirstOperands_7__1, 
         L1FirstOperands_7__0, L1FirstOperands_8__15, L1FirstOperands_8__14, 
         L1FirstOperands_8__13, L1FirstOperands_8__12, L1FirstOperands_8__11, 
         L1FirstOperands_8__10, L1FirstOperands_8__9, L1FirstOperands_8__8, 
         L1FirstOperands_8__7, L1FirstOperands_8__6, L1FirstOperands_8__5, 
         L1FirstOperands_8__4, L1FirstOperands_8__3, L1FirstOperands_8__2, 
         L1FirstOperands_8__1, L1FirstOperands_8__0, L1FirstOperands_10__15, 
         L1FirstOperands_10__14, L1FirstOperands_10__13, L1FirstOperands_10__12, 
         L1FirstOperands_10__11, L1FirstOperands_10__10, L1FirstOperands_10__9, 
         L1FirstOperands_10__8, L1FirstOperands_10__7, L1FirstOperands_10__6, 
         L1FirstOperands_10__5, L1FirstOperands_10__4, L1FirstOperands_10__3, 
         L1FirstOperands_10__2, L1FirstOperands_10__1, L1FirstOperands_10__0, 
         L1FirstOperands_11__15, L1FirstOperands_11__14, L1FirstOperands_11__13, 
         L1FirstOperands_11__12, L1FirstOperands_11__11, L1FirstOperands_11__10, 
         L1FirstOperands_11__9, L1FirstOperands_11__8, L1FirstOperands_11__7, 
         L1FirstOperands_11__6, L1FirstOperands_11__5, L1FirstOperands_11__4, 
         L1FirstOperands_11__3, L1FirstOperands_11__2, L1FirstOperands_11__1, 
         L1FirstOperands_11__0, L1ResultsLarge_0__16, L1ResultsLarge_0__15, 
         L1ResultsLarge_0__14, L1ResultsLarge_0__13, L1ResultsLarge_0__12, 
         L1ResultsLarge_0__11, L1ResultsLarge_0__10, L1ResultsLarge_0__9, 
         L1ResultsLarge_0__8, L1ResultsLarge_0__7, L1ResultsLarge_0__6, 
         L1ResultsLarge_0__5, L1ResultsLarge_0__4, L1ResultsLarge_0__3, 
         L1ResultsLarge_0__2, L1ResultsLarge_0__1, L1ResultsLarge_0__0, 
         L1ResultsLarge_1__16, L1ResultsLarge_1__15, L1ResultsLarge_1__14, 
         L1ResultsLarge_1__13, L1ResultsLarge_1__12, L1ResultsLarge_1__11, 
         L1ResultsLarge_1__10, L1ResultsLarge_1__9, L1ResultsLarge_1__8, 
         L1ResultsLarge_1__7, L1ResultsLarge_1__6, L1ResultsLarge_1__5, 
         L1ResultsLarge_1__4, L1ResultsLarge_1__3, L1ResultsLarge_1__2, 
         L1ResultsLarge_1__1, L1ResultsLarge_1__0, L1ResultsLarge_2__16, 
         L1ResultsLarge_2__15, L1ResultsLarge_2__14, L1ResultsLarge_2__13, 
         L1ResultsLarge_2__12, L1ResultsLarge_2__11, L1ResultsLarge_2__10, 
         L1ResultsLarge_2__9, L1ResultsLarge_2__8, L1ResultsLarge_2__7, 
         L1ResultsLarge_2__6, L1ResultsLarge_2__5, L1ResultsLarge_2__4, 
         L1ResultsLarge_2__3, L1ResultsLarge_2__2, L1ResultsLarge_2__1, 
         L1ResultsLarge_2__0, L1ResultsLarge_3__16, L1ResultsLarge_3__15, 
         L1ResultsLarge_3__14, L1ResultsLarge_3__13, L1ResultsLarge_3__12, 
         L1ResultsLarge_3__11, L1ResultsLarge_3__10, L1ResultsLarge_3__9, 
         L1ResultsLarge_3__8, L1ResultsLarge_3__7, L1ResultsLarge_3__6, 
         L1ResultsLarge_3__5, L1ResultsLarge_3__4, L1ResultsLarge_3__3, 
         L1ResultsLarge_3__2, L1ResultsLarge_3__1, L1ResultsLarge_3__0, 
         L1ResultsLarge_4__16, L1ResultsLarge_4__15, L1ResultsLarge_4__14, 
         L1ResultsLarge_4__13, L1ResultsLarge_4__12, L1ResultsLarge_4__11, 
         L1ResultsLarge_4__10, L1ResultsLarge_4__9, L1ResultsLarge_4__8, 
         L1ResultsLarge_4__7, L1ResultsLarge_4__6, L1ResultsLarge_4__5, 
         L1ResultsLarge_4__4, L1ResultsLarge_4__3, L1ResultsLarge_4__2, 
         L1ResultsLarge_4__1, L1ResultsLarge_4__0, L1ResultsLarge_5__16, 
         L1ResultsLarge_5__15, L1ResultsLarge_5__14, L1ResultsLarge_5__13, 
         L1ResultsLarge_5__12, L1ResultsLarge_5__11, L1ResultsLarge_5__10, 
         L1ResultsLarge_5__9, L1ResultsLarge_5__8, L1ResultsLarge_5__7, 
         L1ResultsLarge_5__6, L1ResultsLarge_5__5, L1ResultsLarge_5__4, 
         L1ResultsLarge_5__3, L1ResultsLarge_5__2, L1ResultsLarge_5__1, 
         L1ResultsLarge_5__0, L1ResultsLarge_6__16, L1ResultsLarge_6__15, 
         L1ResultsLarge_6__14, L1ResultsLarge_6__13, L1ResultsLarge_6__12, 
         L1ResultsLarge_6__11, L1ResultsLarge_6__10, L1ResultsLarge_6__9, 
         L1ResultsLarge_6__8, L1ResultsLarge_6__7, L1ResultsLarge_6__6, 
         L1ResultsLarge_6__5, L1ResultsLarge_6__4, L1ResultsLarge_6__3, 
         L1ResultsLarge_6__2, L1ResultsLarge_6__1, L1ResultsLarge_6__0, 
         L1ResultsLarge_7__16, L1ResultsLarge_7__15, L1ResultsLarge_7__14, 
         L1ResultsLarge_7__13, L1ResultsLarge_7__12, L1ResultsLarge_7__11, 
         L1ResultsLarge_7__10, L1ResultsLarge_7__9, L1ResultsLarge_7__8, 
         L1ResultsLarge_7__7, L1ResultsLarge_7__6, L1ResultsLarge_7__5, 
         L1ResultsLarge_7__4, L1ResultsLarge_7__3, L1ResultsLarge_7__2, 
         L1ResultsLarge_7__1, L1ResultsLarge_7__0, L1ResultsLarge_8__16, 
         L1ResultsLarge_8__15, L1ResultsLarge_8__14, L1ResultsLarge_8__13, 
         L1ResultsLarge_8__12, L1ResultsLarge_8__11, L1ResultsLarge_8__10, 
         L1ResultsLarge_8__9, L1ResultsLarge_8__8, L1ResultsLarge_8__7, 
         L1ResultsLarge_8__6, L1ResultsLarge_8__5, L1ResultsLarge_8__4, 
         L1ResultsLarge_8__3, L1ResultsLarge_8__2, L1ResultsLarge_8__1, 
         L1ResultsLarge_8__0, L1ResultsLarge_9__16, L1ResultsLarge_9__15, 
         L1ResultsLarge_9__14, L1ResultsLarge_9__13, L1ResultsLarge_9__12, 
         L1ResultsLarge_9__11, L1ResultsLarge_9__10, L1ResultsLarge_9__9, 
         L1ResultsLarge_9__8, L1ResultsLarge_9__7, L1ResultsLarge_9__6, 
         L1ResultsLarge_9__5, L1ResultsLarge_9__4, L1ResultsLarge_9__3, 
         L1ResultsLarge_9__2, L1ResultsLarge_9__1, L1ResultsLarge_9__0, 
         L1ResultsLarge_10__16, L1ResultsLarge_10__15, L1ResultsLarge_10__14, 
         L1ResultsLarge_10__13, L1ResultsLarge_10__12, L1ResultsLarge_10__11, 
         L1ResultsLarge_10__10, L1ResultsLarge_10__9, L1ResultsLarge_10__8, 
         L1ResultsLarge_10__7, L1ResultsLarge_10__6, L1ResultsLarge_10__5, 
         L1ResultsLarge_10__4, L1ResultsLarge_10__3, L1ResultsLarge_10__2, 
         L1ResultsLarge_10__1, L1ResultsLarge_10__0, L1ResultsLarge_11__16, 
         L1ResultsLarge_11__15, L1ResultsLarge_11__14, L1ResultsLarge_11__13, 
         L1ResultsLarge_11__12, L1ResultsLarge_11__11, L1ResultsLarge_11__10, 
         L1ResultsLarge_11__9, L1ResultsLarge_11__8, L1ResultsLarge_11__7, 
         L1ResultsLarge_11__6, L1ResultsLarge_11__5, L1ResultsLarge_11__4, 
         L1ResultsLarge_11__3, L1ResultsLarge_11__2, L1ResultsLarge_11__1, 
         L1ResultsLarge_11__0, L2ResultsLarge_0__16, L2ResultsLarge_0__15, 
         L2ResultsLarge_0__14, L2ResultsLarge_0__13, L2ResultsLarge_0__12, 
         L2ResultsLarge_0__11, L2ResultsLarge_0__10, L2ResultsLarge_0__9, 
         L2ResultsLarge_0__8, L2ResultsLarge_0__7, L2ResultsLarge_0__6, 
         L2ResultsLarge_0__5, L2ResultsLarge_0__4, L2ResultsLarge_0__3, 
         L2ResultsLarge_0__2, L2ResultsLarge_0__1, L2ResultsLarge_0__0, 
         L2ResultsLarge_1__16, L2ResultsLarge_1__15, L2ResultsLarge_1__14, 
         L2ResultsLarge_1__13, L2ResultsLarge_1__12, L2ResultsLarge_1__11, 
         L2ResultsLarge_1__10, L2ResultsLarge_1__9, L2ResultsLarge_1__8, 
         L2ResultsLarge_1__7, L2ResultsLarge_1__6, L2ResultsLarge_1__5, 
         L2ResultsLarge_1__4, L2ResultsLarge_1__3, L2ResultsLarge_1__2, 
         L2ResultsLarge_1__1, L2ResultsLarge_1__0, L2ResultsLarge_2__16, 
         L2ResultsLarge_2__15, L2ResultsLarge_2__14, L2ResultsLarge_2__13, 
         L2ResultsLarge_2__12, L2ResultsLarge_2__11, L2ResultsLarge_2__10, 
         L2ResultsLarge_2__9, L2ResultsLarge_2__8, L2ResultsLarge_2__7, 
         L2ResultsLarge_2__6, L2ResultsLarge_2__5, L2ResultsLarge_2__4, 
         L2ResultsLarge_2__3, L2ResultsLarge_2__2, L2ResultsLarge_2__1, 
         L2ResultsLarge_2__0, L2ResultsLarge_3__16, L2ResultsLarge_3__15, 
         L2ResultsLarge_3__14, L2ResultsLarge_3__13, L2ResultsLarge_3__12, 
         L2ResultsLarge_3__11, L2ResultsLarge_3__10, L2ResultsLarge_3__9, 
         L2ResultsLarge_3__8, L2ResultsLarge_3__7, L2ResultsLarge_3__6, 
         L2ResultsLarge_3__5, L2ResultsLarge_3__4, L2ResultsLarge_3__3, 
         L2ResultsLarge_3__2, L2ResultsLarge_3__1, L2ResultsLarge_3__0, 
         L2ResultsLarge_4__16, L2ResultsLarge_4__15, L2ResultsLarge_4__14, 
         L2ResultsLarge_4__13, L2ResultsLarge_4__12, L2ResultsLarge_4__11, 
         L2ResultsLarge_4__10, L2ResultsLarge_4__9, L2ResultsLarge_4__8, 
         L2ResultsLarge_4__7, L2ResultsLarge_4__6, L2ResultsLarge_4__5, 
         L2ResultsLarge_4__4, L2ResultsLarge_4__3, L2ResultsLarge_4__2, 
         L2ResultsLarge_4__1, L2ResultsLarge_4__0, L2ResultsLarge_5__16, 
         L2ResultsLarge_5__15, L2ResultsLarge_5__14, L2ResultsLarge_5__13, 
         L2ResultsLarge_5__12, L2ResultsLarge_5__11, L2ResultsLarge_5__10, 
         L2ResultsLarge_5__9, L2ResultsLarge_5__8, L2ResultsLarge_5__7, 
         L2ResultsLarge_5__6, L2ResultsLarge_5__5, L2ResultsLarge_5__4, 
         L2ResultsLarge_5__3, L2ResultsLarge_5__2, L2ResultsLarge_5__1, 
         L2ResultsLarge_5__0, L3ResultsLarge_0__16, L3ResultsLarge_0__15, 
         L3ResultsLarge_0__14, L3ResultsLarge_0__13, L3ResultsLarge_0__12, 
         L3ResultsLarge_0__11, L3ResultsLarge_0__10, L3ResultsLarge_0__9, 
         L3ResultsLarge_0__8, L3ResultsLarge_0__7, L3ResultsLarge_0__6, 
         L3ResultsLarge_0__5, L3ResultsLarge_0__4, L3ResultsLarge_0__3, 
         L3ResultsLarge_0__2, L3ResultsLarge_0__1, L3ResultsLarge_0__0, 
         L3ResultsLarge_1__16, L3ResultsLarge_1__15, L3ResultsLarge_1__14, 
         L3ResultsLarge_1__13, L3ResultsLarge_1__12, L3ResultsLarge_1__11, 
         L3ResultsLarge_1__10, L3ResultsLarge_1__9, L3ResultsLarge_1__8, 
         L3ResultsLarge_1__7, L3ResultsLarge_1__6, L3ResultsLarge_1__5, 
         L3ResultsLarge_1__4, L3ResultsLarge_1__3, L3ResultsLarge_1__2, 
         L3ResultsLarge_1__1, L3ResultsLarge_1__0, L3ResultsLarge_2__16, 
         L3ResultsLarge_2__15, L3ResultsLarge_2__14, L3ResultsLarge_2__13, 
         L3ResultsLarge_2__12, L3ResultsLarge_2__11, L3ResultsLarge_2__10, 
         L3ResultsLarge_2__9, L3ResultsLarge_2__8, L3ResultsLarge_2__7, 
         L3ResultsLarge_2__6, L3ResultsLarge_2__5, L3ResultsLarge_2__4, 
         L3ResultsLarge_2__3, L3ResultsLarge_2__2, L3ResultsLarge_2__1, 
         L3ResultsLarge_2__0, L4ResultsLarge_0__16, L4ResultsLarge_0__15, 
         L4ResultsLarge_0__14, L4ResultsLarge_0__13, L4ResultsLarge_0__12, 
         L4ResultsLarge_0__11, L4ResultsLarge_0__10, L4ResultsLarge_0__9, 
         L4ResultsLarge_0__8, L4ResultsLarge_0__7, L4ResultsLarge_0__6, 
         L4ResultsLarge_0__5, L4ResultsLarge_0__4, L4ResultsLarge_0__3, 
         L4ResultsLarge_0__2, L4ResultsLarge_0__1, L4ResultsLarge_0__0, 
         L5FirstOperands_1__16, L5FirstOperands_1__15, L5FirstOperands_1__14, 
         L5FirstOperands_1__13, L5FirstOperands_1__12, L5FirstOperands_1__11, 
         L5FirstOperands_1__10, L5FirstOperands_1__9, L5FirstOperands_1__8, 
         L5FirstOperands_1__7, L5FirstOperands_1__6, L5FirstOperands_1__5, 
         L5FirstOperands_1__4, L5FirstOperands_1__3, L5FirstOperands_1__2, 
         L5FirstOperands_1__1, L5FirstOperands_1__0, 
         L1_0_L2_0_G1_MINI_ALU_OperationResult_15, 
         L1_0_L2_0_G1_MINI_ALU_OperationResult_14, 
         L1_0_L2_0_G1_MINI_ALU_OperationResult_13, 
         L1_0_L2_0_G1_MINI_ALU_OperationResult_12, 
         L1_0_L2_0_G1_MINI_ALU_OperationResult_11, 
         L1_0_L2_0_G1_MINI_ALU_OperationResult_10, 
         L1_0_L2_0_G1_MINI_ALU_OperationResult_9, 
         L1_0_L2_0_G1_MINI_ALU_OperationResult_8, 
         L1_0_L2_0_G1_MINI_ALU_OperationResult_7, 
         L1_0_L2_0_G1_MINI_ALU_OperationResult_6, 
         L1_0_L2_0_G1_MINI_ALU_OperationResult_5, 
         L1_0_L2_0_G1_MINI_ALU_OperationResult_4, 
         L1_0_L2_0_G1_MINI_ALU_OperationResult_3, 
         L1_0_L2_0_G1_MINI_ALU_OperationResult_2, 
         L1_0_L2_0_G1_MINI_ALU_OperationResult_1, 
         L1_0_L2_0_G1_MINI_ALU_OperationResult_0, 
         L1_0_L2_0_G1_MINI_ALU_BoothXORCheck, 
         L1_0_L2_0_G1_MINI_ALU_BoothOperand_16, 
         L1_0_L2_0_G1_MINI_ALU_BoothOperand_15, 
         L1_0_L2_0_G1_MINI_ALU_BoothOperand_14, 
         L1_0_L2_0_G1_MINI_ALU_BoothOperand_13, 
         L1_0_L2_0_G1_MINI_ALU_BoothOperand_12, 
         L1_0_L2_0_G1_MINI_ALU_BoothOperand_11, 
         L1_0_L2_0_G1_MINI_ALU_BoothOperand_10, 
         L1_0_L2_0_G1_MINI_ALU_BoothOperand_9, L1_0_L2_0_G1_MINI_ALU_BoothP_16, 
         L1_0_L2_0_G1_MINI_ALU_BoothP_15, L1_0_L2_0_G1_MINI_ALU_BoothP_14, 
         L1_0_L2_0_G1_MINI_ALU_BoothP_13, L1_0_L2_0_G1_MINI_ALU_BoothP_12, 
         L1_0_L2_0_G1_MINI_ALU_BoothP_11, L1_0_L2_0_G1_MINI_ALU_BoothP_10, 
         L1_0_L2_0_G1_MINI_ALU_BoothP_9, L1_0_L2_0_G1_MINI_ALU_BoothP_8, 
         L1_0_L2_0_G1_MINI_ALU_BoothP_7, L1_0_L2_0_G1_MINI_ALU_BoothP_6, 
         L1_0_L2_0_G1_MINI_ALU_BoothP_5, L1_0_L2_0_G1_MINI_ALU_BoothP_4, 
         L1_0_L2_0_G1_MINI_ALU_BoothP_3, L1_0_L2_0_G1_MINI_ALU_BoothP_2, 
         L1_0_L2_0_G1_MINI_ALU_BoothP_1, L1_0_L2_0_G1_MINI_ALU_BoothP_0, 
         L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_15, 
         L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_14, 
         L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_13, 
         L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_12, 
         L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_11, 
         L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_10, 
         L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_9, 
         L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_8, 
         L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_7, 
         L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_6, 
         L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_5, 
         L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_4, 
         L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_3, 
         L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_2, 
         L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_1, 
         L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_0, 
         L1_0_L2_1_G1_MINI_ALU_OperationResult_15, 
         L1_0_L2_1_G1_MINI_ALU_OperationResult_14, 
         L1_0_L2_1_G1_MINI_ALU_OperationResult_13, 
         L1_0_L2_1_G1_MINI_ALU_OperationResult_12, 
         L1_0_L2_1_G1_MINI_ALU_OperationResult_11, 
         L1_0_L2_1_G1_MINI_ALU_OperationResult_10, 
         L1_0_L2_1_G1_MINI_ALU_OperationResult_9, 
         L1_0_L2_1_G1_MINI_ALU_OperationResult_8, 
         L1_0_L2_1_G1_MINI_ALU_OperationResult_7, 
         L1_0_L2_1_G1_MINI_ALU_OperationResult_6, 
         L1_0_L2_1_G1_MINI_ALU_OperationResult_5, 
         L1_0_L2_1_G1_MINI_ALU_OperationResult_4, 
         L1_0_L2_1_G1_MINI_ALU_OperationResult_3, 
         L1_0_L2_1_G1_MINI_ALU_OperationResult_2, 
         L1_0_L2_1_G1_MINI_ALU_OperationResult_1, 
         L1_0_L2_1_G1_MINI_ALU_OperationResult_0, 
         L1_0_L2_1_G1_MINI_ALU_BoothXORCheck, 
         L1_0_L2_1_G1_MINI_ALU_BoothOperand_16, 
         L1_0_L2_1_G1_MINI_ALU_BoothOperand_15, 
         L1_0_L2_1_G1_MINI_ALU_BoothOperand_14, 
         L1_0_L2_1_G1_MINI_ALU_BoothOperand_13, 
         L1_0_L2_1_G1_MINI_ALU_BoothOperand_12, 
         L1_0_L2_1_G1_MINI_ALU_BoothOperand_11, 
         L1_0_L2_1_G1_MINI_ALU_BoothOperand_10, 
         L1_0_L2_1_G1_MINI_ALU_BoothOperand_9, L1_0_L2_1_G1_MINI_ALU_BoothP_16, 
         L1_0_L2_1_G1_MINI_ALU_BoothP_15, L1_0_L2_1_G1_MINI_ALU_BoothP_14, 
         L1_0_L2_1_G1_MINI_ALU_BoothP_13, L1_0_L2_1_G1_MINI_ALU_BoothP_12, 
         L1_0_L2_1_G1_MINI_ALU_BoothP_11, L1_0_L2_1_G1_MINI_ALU_BoothP_10, 
         L1_0_L2_1_G1_MINI_ALU_BoothP_9, L1_0_L2_1_G1_MINI_ALU_BoothP_8, 
         L1_0_L2_1_G1_MINI_ALU_BoothP_7, L1_0_L2_1_G1_MINI_ALU_BoothP_6, 
         L1_0_L2_1_G1_MINI_ALU_BoothP_5, L1_0_L2_1_G1_MINI_ALU_BoothP_4, 
         L1_0_L2_1_G1_MINI_ALU_BoothP_3, L1_0_L2_1_G1_MINI_ALU_BoothP_2, 
         L1_0_L2_1_G1_MINI_ALU_BoothP_1, L1_0_L2_1_G1_MINI_ALU_BoothP_0, 
         L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_15, 
         L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_14, 
         L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_13, 
         L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_12, 
         L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_11, 
         L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_10, 
         L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_9, 
         L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_8, 
         L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_7, 
         L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_6, 
         L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_5, 
         L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_4, 
         L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_3, 
         L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_2, 
         L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_1, 
         L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_0, 
         L1_0_L2_2_G1_MINI_ALU_OperationResult_15, 
         L1_0_L2_2_G1_MINI_ALU_OperationResult_14, 
         L1_0_L2_2_G1_MINI_ALU_OperationResult_13, 
         L1_0_L2_2_G1_MINI_ALU_OperationResult_12, 
         L1_0_L2_2_G1_MINI_ALU_OperationResult_11, 
         L1_0_L2_2_G1_MINI_ALU_OperationResult_10, 
         L1_0_L2_2_G1_MINI_ALU_OperationResult_9, 
         L1_0_L2_2_G1_MINI_ALU_OperationResult_8, 
         L1_0_L2_2_G1_MINI_ALU_OperationResult_7, 
         L1_0_L2_2_G1_MINI_ALU_OperationResult_6, 
         L1_0_L2_2_G1_MINI_ALU_OperationResult_5, 
         L1_0_L2_2_G1_MINI_ALU_OperationResult_4, 
         L1_0_L2_2_G1_MINI_ALU_OperationResult_3, 
         L1_0_L2_2_G1_MINI_ALU_OperationResult_2, 
         L1_0_L2_2_G1_MINI_ALU_OperationResult_1, 
         L1_0_L2_2_G1_MINI_ALU_OperationResult_0, 
         L1_0_L2_2_G1_MINI_ALU_BoothXORCheck, 
         L1_0_L2_2_G1_MINI_ALU_BoothOperand_16, 
         L1_0_L2_2_G1_MINI_ALU_BoothOperand_15, 
         L1_0_L2_2_G1_MINI_ALU_BoothOperand_14, 
         L1_0_L2_2_G1_MINI_ALU_BoothOperand_13, 
         L1_0_L2_2_G1_MINI_ALU_BoothOperand_12, 
         L1_0_L2_2_G1_MINI_ALU_BoothOperand_11, 
         L1_0_L2_2_G1_MINI_ALU_BoothOperand_10, 
         L1_0_L2_2_G1_MINI_ALU_BoothOperand_9, L1_0_L2_2_G1_MINI_ALU_BoothP_16, 
         L1_0_L2_2_G1_MINI_ALU_BoothP_15, L1_0_L2_2_G1_MINI_ALU_BoothP_14, 
         L1_0_L2_2_G1_MINI_ALU_BoothP_13, L1_0_L2_2_G1_MINI_ALU_BoothP_12, 
         L1_0_L2_2_G1_MINI_ALU_BoothP_11, L1_0_L2_2_G1_MINI_ALU_BoothP_10, 
         L1_0_L2_2_G1_MINI_ALU_BoothP_9, L1_0_L2_2_G1_MINI_ALU_BoothP_8, 
         L1_0_L2_2_G1_MINI_ALU_BoothP_7, L1_0_L2_2_G1_MINI_ALU_BoothP_6, 
         L1_0_L2_2_G1_MINI_ALU_BoothP_5, L1_0_L2_2_G1_MINI_ALU_BoothP_4, 
         L1_0_L2_2_G1_MINI_ALU_BoothP_3, L1_0_L2_2_G1_MINI_ALU_BoothP_2, 
         L1_0_L2_2_G1_MINI_ALU_BoothP_1, L1_0_L2_2_G1_MINI_ALU_BoothP_0, 
         L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_15, 
         L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_14, 
         L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_13, 
         L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_12, 
         L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_11, 
         L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_10, 
         L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_9, 
         L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_8, 
         L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_7, 
         L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_6, 
         L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_5, 
         L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_4, 
         L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_3, 
         L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_2, 
         L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_1, 
         L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_0, 
         L1_0_L2_3_G1_MINI_ALU_OperationResult_15, 
         L1_0_L2_3_G1_MINI_ALU_OperationResult_14, 
         L1_0_L2_3_G1_MINI_ALU_OperationResult_13, 
         L1_0_L2_3_G1_MINI_ALU_OperationResult_12, 
         L1_0_L2_3_G1_MINI_ALU_OperationResult_11, 
         L1_0_L2_3_G1_MINI_ALU_OperationResult_10, 
         L1_0_L2_3_G1_MINI_ALU_OperationResult_9, 
         L1_0_L2_3_G1_MINI_ALU_OperationResult_8, 
         L1_0_L2_3_G1_MINI_ALU_OperationResult_7, 
         L1_0_L2_3_G1_MINI_ALU_OperationResult_6, 
         L1_0_L2_3_G1_MINI_ALU_OperationResult_5, 
         L1_0_L2_3_G1_MINI_ALU_OperationResult_4, 
         L1_0_L2_3_G1_MINI_ALU_OperationResult_3, 
         L1_0_L2_3_G1_MINI_ALU_OperationResult_2, 
         L1_0_L2_3_G1_MINI_ALU_OperationResult_1, 
         L1_0_L2_3_G1_MINI_ALU_OperationResult_0, 
         L1_0_L2_3_G1_MINI_ALU_BoothXORCheck, 
         L1_0_L2_3_G1_MINI_ALU_BoothOperand_16, 
         L1_0_L2_3_G1_MINI_ALU_BoothOperand_15, 
         L1_0_L2_3_G1_MINI_ALU_BoothOperand_14, 
         L1_0_L2_3_G1_MINI_ALU_BoothOperand_13, 
         L1_0_L2_3_G1_MINI_ALU_BoothOperand_12, 
         L1_0_L2_3_G1_MINI_ALU_BoothOperand_11, 
         L1_0_L2_3_G1_MINI_ALU_BoothOperand_10, 
         L1_0_L2_3_G1_MINI_ALU_BoothOperand_9, L1_0_L2_3_G1_MINI_ALU_BoothP_16, 
         L1_0_L2_3_G1_MINI_ALU_BoothP_15, L1_0_L2_3_G1_MINI_ALU_BoothP_14, 
         L1_0_L2_3_G1_MINI_ALU_BoothP_13, L1_0_L2_3_G1_MINI_ALU_BoothP_12, 
         L1_0_L2_3_G1_MINI_ALU_BoothP_11, L1_0_L2_3_G1_MINI_ALU_BoothP_10, 
         L1_0_L2_3_G1_MINI_ALU_BoothP_9, L1_0_L2_3_G1_MINI_ALU_BoothP_8, 
         L1_0_L2_3_G1_MINI_ALU_BoothP_7, L1_0_L2_3_G1_MINI_ALU_BoothP_6, 
         L1_0_L2_3_G1_MINI_ALU_BoothP_5, L1_0_L2_3_G1_MINI_ALU_BoothP_4, 
         L1_0_L2_3_G1_MINI_ALU_BoothP_3, L1_0_L2_3_G1_MINI_ALU_BoothP_2, 
         L1_0_L2_3_G1_MINI_ALU_BoothP_1, L1_0_L2_3_G1_MINI_ALU_BoothP_0, 
         L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_15, 
         L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_14, 
         L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_13, 
         L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_12, 
         L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_11, 
         L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_10, 
         L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_9, 
         L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_8, 
         L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_7, 
         L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_6, 
         L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_5, 
         L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_4, 
         L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_3, 
         L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_2, 
         L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_1, 
         L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_0, 
         L1_0_L2_4_G1_MINI_ALU_OperationResult_15, 
         L1_0_L2_4_G1_MINI_ALU_OperationResult_14, 
         L1_0_L2_4_G1_MINI_ALU_OperationResult_13, 
         L1_0_L2_4_G1_MINI_ALU_OperationResult_12, 
         L1_0_L2_4_G1_MINI_ALU_OperationResult_11, 
         L1_0_L2_4_G1_MINI_ALU_OperationResult_10, 
         L1_0_L2_4_G1_MINI_ALU_OperationResult_9, 
         L1_0_L2_4_G1_MINI_ALU_OperationResult_8, 
         L1_0_L2_4_G1_MINI_ALU_OperationResult_7, 
         L1_0_L2_4_G1_MINI_ALU_OperationResult_6, 
         L1_0_L2_4_G1_MINI_ALU_OperationResult_5, 
         L1_0_L2_4_G1_MINI_ALU_OperationResult_4, 
         L1_0_L2_4_G1_MINI_ALU_OperationResult_3, 
         L1_0_L2_4_G1_MINI_ALU_OperationResult_2, 
         L1_0_L2_4_G1_MINI_ALU_OperationResult_1, 
         L1_0_L2_4_G1_MINI_ALU_OperationResult_0, 
         L1_0_L2_4_G1_MINI_ALU_BoothXORCheck, 
         L1_0_L2_4_G1_MINI_ALU_BoothOperand_16, 
         L1_0_L2_4_G1_MINI_ALU_BoothOperand_15, 
         L1_0_L2_4_G1_MINI_ALU_BoothOperand_14, 
         L1_0_L2_4_G1_MINI_ALU_BoothOperand_13, 
         L1_0_L2_4_G1_MINI_ALU_BoothOperand_12, 
         L1_0_L2_4_G1_MINI_ALU_BoothOperand_11, 
         L1_0_L2_4_G1_MINI_ALU_BoothOperand_10, 
         L1_0_L2_4_G1_MINI_ALU_BoothOperand_9, L1_0_L2_4_G1_MINI_ALU_BoothP_16, 
         L1_0_L2_4_G1_MINI_ALU_BoothP_15, L1_0_L2_4_G1_MINI_ALU_BoothP_14, 
         L1_0_L2_4_G1_MINI_ALU_BoothP_13, L1_0_L2_4_G1_MINI_ALU_BoothP_12, 
         L1_0_L2_4_G1_MINI_ALU_BoothP_11, L1_0_L2_4_G1_MINI_ALU_BoothP_10, 
         L1_0_L2_4_G1_MINI_ALU_BoothP_9, L1_0_L2_4_G1_MINI_ALU_BoothP_8, 
         L1_0_L2_4_G1_MINI_ALU_BoothP_7, L1_0_L2_4_G1_MINI_ALU_BoothP_6, 
         L1_0_L2_4_G1_MINI_ALU_BoothP_5, L1_0_L2_4_G1_MINI_ALU_BoothP_4, 
         L1_0_L2_4_G1_MINI_ALU_BoothP_3, L1_0_L2_4_G1_MINI_ALU_BoothP_2, 
         L1_0_L2_4_G1_MINI_ALU_BoothP_1, L1_0_L2_4_G1_MINI_ALU_BoothP_0, 
         L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_15, 
         L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_14, 
         L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_13, 
         L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_12, 
         L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_11, 
         L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_10, 
         L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_9, 
         L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_8, 
         L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_7, 
         L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_6, 
         L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_5, 
         L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_4, 
         L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_3, 
         L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_2, 
         L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_1, 
         L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_0, 
         L1_1_L2_0_G1_MINI_ALU_OperationResult_15, 
         L1_1_L2_0_G1_MINI_ALU_OperationResult_14, 
         L1_1_L2_0_G1_MINI_ALU_OperationResult_13, 
         L1_1_L2_0_G1_MINI_ALU_OperationResult_12, 
         L1_1_L2_0_G1_MINI_ALU_OperationResult_11, 
         L1_1_L2_0_G1_MINI_ALU_OperationResult_10, 
         L1_1_L2_0_G1_MINI_ALU_OperationResult_9, 
         L1_1_L2_0_G1_MINI_ALU_OperationResult_8, 
         L1_1_L2_0_G1_MINI_ALU_OperationResult_7, 
         L1_1_L2_0_G1_MINI_ALU_OperationResult_6, 
         L1_1_L2_0_G1_MINI_ALU_OperationResult_5, 
         L1_1_L2_0_G1_MINI_ALU_OperationResult_4, 
         L1_1_L2_0_G1_MINI_ALU_OperationResult_3, 
         L1_1_L2_0_G1_MINI_ALU_OperationResult_2, 
         L1_1_L2_0_G1_MINI_ALU_OperationResult_1, 
         L1_1_L2_0_G1_MINI_ALU_OperationResult_0, 
         L1_1_L2_0_G1_MINI_ALU_BoothXORCheck, 
         L1_1_L2_0_G1_MINI_ALU_BoothOperand_16, 
         L1_1_L2_0_G1_MINI_ALU_BoothOperand_15, 
         L1_1_L2_0_G1_MINI_ALU_BoothOperand_14, 
         L1_1_L2_0_G1_MINI_ALU_BoothOperand_13, 
         L1_1_L2_0_G1_MINI_ALU_BoothOperand_12, 
         L1_1_L2_0_G1_MINI_ALU_BoothOperand_11, 
         L1_1_L2_0_G1_MINI_ALU_BoothOperand_10, 
         L1_1_L2_0_G1_MINI_ALU_BoothOperand_9, L1_1_L2_0_G1_MINI_ALU_BoothP_16, 
         L1_1_L2_0_G1_MINI_ALU_BoothP_15, L1_1_L2_0_G1_MINI_ALU_BoothP_14, 
         L1_1_L2_0_G1_MINI_ALU_BoothP_13, L1_1_L2_0_G1_MINI_ALU_BoothP_12, 
         L1_1_L2_0_G1_MINI_ALU_BoothP_11, L1_1_L2_0_G1_MINI_ALU_BoothP_10, 
         L1_1_L2_0_G1_MINI_ALU_BoothP_9, L1_1_L2_0_G1_MINI_ALU_BoothP_8, 
         L1_1_L2_0_G1_MINI_ALU_BoothP_7, L1_1_L2_0_G1_MINI_ALU_BoothP_6, 
         L1_1_L2_0_G1_MINI_ALU_BoothP_5, L1_1_L2_0_G1_MINI_ALU_BoothP_4, 
         L1_1_L2_0_G1_MINI_ALU_BoothP_3, L1_1_L2_0_G1_MINI_ALU_BoothP_2, 
         L1_1_L2_0_G1_MINI_ALU_BoothP_1, L1_1_L2_0_G1_MINI_ALU_BoothP_0, 
         L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_15, 
         L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_14, 
         L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_13, 
         L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_12, 
         L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_11, 
         L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_10, 
         L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_9, 
         L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_8, 
         L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_7, 
         L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_6, 
         L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_5, 
         L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_4, 
         L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_3, 
         L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_2, 
         L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_1, 
         L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_0, 
         L1_1_L2_1_G1_MINI_ALU_OperationResult_15, 
         L1_1_L2_1_G1_MINI_ALU_OperationResult_14, 
         L1_1_L2_1_G1_MINI_ALU_OperationResult_13, 
         L1_1_L2_1_G1_MINI_ALU_OperationResult_12, 
         L1_1_L2_1_G1_MINI_ALU_OperationResult_11, 
         L1_1_L2_1_G1_MINI_ALU_OperationResult_10, 
         L1_1_L2_1_G1_MINI_ALU_OperationResult_9, 
         L1_1_L2_1_G1_MINI_ALU_OperationResult_8, 
         L1_1_L2_1_G1_MINI_ALU_OperationResult_7, 
         L1_1_L2_1_G1_MINI_ALU_OperationResult_6, 
         L1_1_L2_1_G1_MINI_ALU_OperationResult_5, 
         L1_1_L2_1_G1_MINI_ALU_OperationResult_4, 
         L1_1_L2_1_G1_MINI_ALU_OperationResult_3, 
         L1_1_L2_1_G1_MINI_ALU_OperationResult_2, 
         L1_1_L2_1_G1_MINI_ALU_OperationResult_1, 
         L1_1_L2_1_G1_MINI_ALU_OperationResult_0, 
         L1_1_L2_1_G1_MINI_ALU_BoothXORCheck, 
         L1_1_L2_1_G1_MINI_ALU_BoothOperand_16, 
         L1_1_L2_1_G1_MINI_ALU_BoothOperand_15, 
         L1_1_L2_1_G1_MINI_ALU_BoothOperand_14, 
         L1_1_L2_1_G1_MINI_ALU_BoothOperand_13, 
         L1_1_L2_1_G1_MINI_ALU_BoothOperand_12, 
         L1_1_L2_1_G1_MINI_ALU_BoothOperand_11, 
         L1_1_L2_1_G1_MINI_ALU_BoothOperand_10, 
         L1_1_L2_1_G1_MINI_ALU_BoothOperand_9, L1_1_L2_1_G1_MINI_ALU_BoothP_16, 
         L1_1_L2_1_G1_MINI_ALU_BoothP_15, L1_1_L2_1_G1_MINI_ALU_BoothP_14, 
         L1_1_L2_1_G1_MINI_ALU_BoothP_13, L1_1_L2_1_G1_MINI_ALU_BoothP_12, 
         L1_1_L2_1_G1_MINI_ALU_BoothP_11, L1_1_L2_1_G1_MINI_ALU_BoothP_10, 
         L1_1_L2_1_G1_MINI_ALU_BoothP_9, L1_1_L2_1_G1_MINI_ALU_BoothP_8, 
         L1_1_L2_1_G1_MINI_ALU_BoothP_7, L1_1_L2_1_G1_MINI_ALU_BoothP_6, 
         L1_1_L2_1_G1_MINI_ALU_BoothP_5, L1_1_L2_1_G1_MINI_ALU_BoothP_4, 
         L1_1_L2_1_G1_MINI_ALU_BoothP_3, L1_1_L2_1_G1_MINI_ALU_BoothP_2, 
         L1_1_L2_1_G1_MINI_ALU_BoothP_1, L1_1_L2_1_G1_MINI_ALU_BoothP_0, 
         L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_15, 
         L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_14, 
         L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_13, 
         L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_12, 
         L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_11, 
         L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_10, 
         L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_9, 
         L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_8, 
         L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_7, 
         L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_6, 
         L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_5, 
         L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_4, 
         L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_3, 
         L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_2, 
         L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_1, 
         L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_0, 
         L1_1_L2_2_G1_MINI_ALU_OperationResult_15, 
         L1_1_L2_2_G1_MINI_ALU_OperationResult_14, 
         L1_1_L2_2_G1_MINI_ALU_OperationResult_13, 
         L1_1_L2_2_G1_MINI_ALU_OperationResult_12, 
         L1_1_L2_2_G1_MINI_ALU_OperationResult_11, 
         L1_1_L2_2_G1_MINI_ALU_OperationResult_10, 
         L1_1_L2_2_G1_MINI_ALU_OperationResult_9, 
         L1_1_L2_2_G1_MINI_ALU_OperationResult_8, 
         L1_1_L2_2_G1_MINI_ALU_OperationResult_7, 
         L1_1_L2_2_G1_MINI_ALU_OperationResult_6, 
         L1_1_L2_2_G1_MINI_ALU_OperationResult_5, 
         L1_1_L2_2_G1_MINI_ALU_OperationResult_4, 
         L1_1_L2_2_G1_MINI_ALU_OperationResult_3, 
         L1_1_L2_2_G1_MINI_ALU_OperationResult_2, 
         L1_1_L2_2_G1_MINI_ALU_OperationResult_1, 
         L1_1_L2_2_G1_MINI_ALU_OperationResult_0, 
         L1_1_L2_2_G1_MINI_ALU_BoothXORCheck, 
         L1_1_L2_2_G1_MINI_ALU_BoothOperand_16, 
         L1_1_L2_2_G1_MINI_ALU_BoothOperand_15, 
         L1_1_L2_2_G1_MINI_ALU_BoothOperand_14, 
         L1_1_L2_2_G1_MINI_ALU_BoothOperand_13, 
         L1_1_L2_2_G1_MINI_ALU_BoothOperand_12, 
         L1_1_L2_2_G1_MINI_ALU_BoothOperand_11, 
         L1_1_L2_2_G1_MINI_ALU_BoothOperand_10, 
         L1_1_L2_2_G1_MINI_ALU_BoothOperand_9, L1_1_L2_2_G1_MINI_ALU_BoothP_16, 
         L1_1_L2_2_G1_MINI_ALU_BoothP_15, L1_1_L2_2_G1_MINI_ALU_BoothP_14, 
         L1_1_L2_2_G1_MINI_ALU_BoothP_13, L1_1_L2_2_G1_MINI_ALU_BoothP_12, 
         L1_1_L2_2_G1_MINI_ALU_BoothP_11, L1_1_L2_2_G1_MINI_ALU_BoothP_10, 
         L1_1_L2_2_G1_MINI_ALU_BoothP_9, L1_1_L2_2_G1_MINI_ALU_BoothP_8, 
         L1_1_L2_2_G1_MINI_ALU_BoothP_7, L1_1_L2_2_G1_MINI_ALU_BoothP_6, 
         L1_1_L2_2_G1_MINI_ALU_BoothP_5, L1_1_L2_2_G1_MINI_ALU_BoothP_4, 
         L1_1_L2_2_G1_MINI_ALU_BoothP_3, L1_1_L2_2_G1_MINI_ALU_BoothP_2, 
         L1_1_L2_2_G1_MINI_ALU_BoothP_1, L1_1_L2_2_G1_MINI_ALU_BoothP_0, 
         L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_15, 
         L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_14, 
         L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_13, 
         L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_12, 
         L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_11, 
         L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_10, 
         L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_9, 
         L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_8, 
         L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_7, 
         L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_6, 
         L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_5, 
         L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_4, 
         L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_3, 
         L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_2, 
         L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_1, 
         L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_0, 
         L1_1_L2_3_G1_MINI_ALU_OperationResult_15, 
         L1_1_L2_3_G1_MINI_ALU_OperationResult_14, 
         L1_1_L2_3_G1_MINI_ALU_OperationResult_13, 
         L1_1_L2_3_G1_MINI_ALU_OperationResult_12, 
         L1_1_L2_3_G1_MINI_ALU_OperationResult_11, 
         L1_1_L2_3_G1_MINI_ALU_OperationResult_10, 
         L1_1_L2_3_G1_MINI_ALU_OperationResult_9, 
         L1_1_L2_3_G1_MINI_ALU_OperationResult_8, 
         L1_1_L2_3_G1_MINI_ALU_OperationResult_7, 
         L1_1_L2_3_G1_MINI_ALU_OperationResult_6, 
         L1_1_L2_3_G1_MINI_ALU_OperationResult_5, 
         L1_1_L2_3_G1_MINI_ALU_OperationResult_4, 
         L1_1_L2_3_G1_MINI_ALU_OperationResult_3, 
         L1_1_L2_3_G1_MINI_ALU_OperationResult_2, 
         L1_1_L2_3_G1_MINI_ALU_OperationResult_1, 
         L1_1_L2_3_G1_MINI_ALU_OperationResult_0, 
         L1_1_L2_3_G1_MINI_ALU_BoothXORCheck, 
         L1_1_L2_3_G1_MINI_ALU_BoothOperand_16, 
         L1_1_L2_3_G1_MINI_ALU_BoothOperand_15, 
         L1_1_L2_3_G1_MINI_ALU_BoothOperand_14, 
         L1_1_L2_3_G1_MINI_ALU_BoothOperand_13, 
         L1_1_L2_3_G1_MINI_ALU_BoothOperand_12, 
         L1_1_L2_3_G1_MINI_ALU_BoothOperand_11, 
         L1_1_L2_3_G1_MINI_ALU_BoothOperand_10, 
         L1_1_L2_3_G1_MINI_ALU_BoothOperand_9, L1_1_L2_3_G1_MINI_ALU_BoothP_16, 
         L1_1_L2_3_G1_MINI_ALU_BoothP_15, L1_1_L2_3_G1_MINI_ALU_BoothP_14, 
         L1_1_L2_3_G1_MINI_ALU_BoothP_13, L1_1_L2_3_G1_MINI_ALU_BoothP_12, 
         L1_1_L2_3_G1_MINI_ALU_BoothP_11, L1_1_L2_3_G1_MINI_ALU_BoothP_10, 
         L1_1_L2_3_G1_MINI_ALU_BoothP_9, L1_1_L2_3_G1_MINI_ALU_BoothP_8, 
         L1_1_L2_3_G1_MINI_ALU_BoothP_7, L1_1_L2_3_G1_MINI_ALU_BoothP_6, 
         L1_1_L2_3_G1_MINI_ALU_BoothP_5, L1_1_L2_3_G1_MINI_ALU_BoothP_4, 
         L1_1_L2_3_G1_MINI_ALU_BoothP_3, L1_1_L2_3_G1_MINI_ALU_BoothP_2, 
         L1_1_L2_3_G1_MINI_ALU_BoothP_1, L1_1_L2_3_G1_MINI_ALU_BoothP_0, 
         L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_15, 
         L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_14, 
         L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_13, 
         L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_12, 
         L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_11, 
         L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_10, 
         L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_9, 
         L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_8, 
         L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_7, 
         L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_6, 
         L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_5, 
         L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_4, 
         L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_3, 
         L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_2, 
         L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_1, 
         L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_0, 
         L1_1_L2_4_G1_MINI_ALU_OperationResult_15, 
         L1_1_L2_4_G1_MINI_ALU_OperationResult_14, 
         L1_1_L2_4_G1_MINI_ALU_OperationResult_13, 
         L1_1_L2_4_G1_MINI_ALU_OperationResult_12, 
         L1_1_L2_4_G1_MINI_ALU_OperationResult_11, 
         L1_1_L2_4_G1_MINI_ALU_OperationResult_10, 
         L1_1_L2_4_G1_MINI_ALU_OperationResult_9, 
         L1_1_L2_4_G1_MINI_ALU_OperationResult_8, 
         L1_1_L2_4_G1_MINI_ALU_OperationResult_7, 
         L1_1_L2_4_G1_MINI_ALU_OperationResult_6, 
         L1_1_L2_4_G1_MINI_ALU_OperationResult_5, 
         L1_1_L2_4_G1_MINI_ALU_OperationResult_4, 
         L1_1_L2_4_G1_MINI_ALU_OperationResult_3, 
         L1_1_L2_4_G1_MINI_ALU_OperationResult_2, 
         L1_1_L2_4_G1_MINI_ALU_OperationResult_1, 
         L1_1_L2_4_G1_MINI_ALU_OperationResult_0, 
         L1_1_L2_4_G1_MINI_ALU_BoothXORCheck, 
         L1_1_L2_4_G1_MINI_ALU_BoothOperand_16, 
         L1_1_L2_4_G1_MINI_ALU_BoothOperand_15, 
         L1_1_L2_4_G1_MINI_ALU_BoothOperand_14, 
         L1_1_L2_4_G1_MINI_ALU_BoothOperand_13, 
         L1_1_L2_4_G1_MINI_ALU_BoothOperand_12, 
         L1_1_L2_4_G1_MINI_ALU_BoothOperand_11, 
         L1_1_L2_4_G1_MINI_ALU_BoothOperand_10, 
         L1_1_L2_4_G1_MINI_ALU_BoothOperand_9, L1_1_L2_4_G1_MINI_ALU_BoothP_16, 
         L1_1_L2_4_G1_MINI_ALU_BoothP_15, L1_1_L2_4_G1_MINI_ALU_BoothP_14, 
         L1_1_L2_4_G1_MINI_ALU_BoothP_13, L1_1_L2_4_G1_MINI_ALU_BoothP_12, 
         L1_1_L2_4_G1_MINI_ALU_BoothP_11, L1_1_L2_4_G1_MINI_ALU_BoothP_10, 
         L1_1_L2_4_G1_MINI_ALU_BoothP_9, L1_1_L2_4_G1_MINI_ALU_BoothP_8, 
         L1_1_L2_4_G1_MINI_ALU_BoothP_7, L1_1_L2_4_G1_MINI_ALU_BoothP_6, 
         L1_1_L2_4_G1_MINI_ALU_BoothP_5, L1_1_L2_4_G1_MINI_ALU_BoothP_4, 
         L1_1_L2_4_G1_MINI_ALU_BoothP_3, L1_1_L2_4_G1_MINI_ALU_BoothP_2, 
         L1_1_L2_4_G1_MINI_ALU_BoothP_1, L1_1_L2_4_G1_MINI_ALU_BoothP_0, 
         L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_15, 
         L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_14, 
         L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_13, 
         L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_12, 
         L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_11, 
         L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_10, 
         L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_9, 
         L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_8, 
         L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_7, 
         L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_6, 
         L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_5, 
         L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_4, 
         L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_3, 
         L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_2, 
         L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_1, 
         L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_0, 
         L1_2_L2_0_G1_MINI_ALU_OperationResult_15, 
         L1_2_L2_0_G1_MINI_ALU_OperationResult_14, 
         L1_2_L2_0_G1_MINI_ALU_OperationResult_13, 
         L1_2_L2_0_G1_MINI_ALU_OperationResult_12, 
         L1_2_L2_0_G1_MINI_ALU_OperationResult_11, 
         L1_2_L2_0_G1_MINI_ALU_OperationResult_10, 
         L1_2_L2_0_G1_MINI_ALU_OperationResult_9, 
         L1_2_L2_0_G1_MINI_ALU_OperationResult_8, 
         L1_2_L2_0_G1_MINI_ALU_OperationResult_7, 
         L1_2_L2_0_G1_MINI_ALU_OperationResult_6, 
         L1_2_L2_0_G1_MINI_ALU_OperationResult_5, 
         L1_2_L2_0_G1_MINI_ALU_OperationResult_4, 
         L1_2_L2_0_G1_MINI_ALU_OperationResult_3, 
         L1_2_L2_0_G1_MINI_ALU_OperationResult_2, 
         L1_2_L2_0_G1_MINI_ALU_OperationResult_1, 
         L1_2_L2_0_G1_MINI_ALU_OperationResult_0, 
         L1_2_L2_0_G1_MINI_ALU_BoothXORCheck, 
         L1_2_L2_0_G1_MINI_ALU_BoothOperand_16, 
         L1_2_L2_0_G1_MINI_ALU_BoothOperand_15, 
         L1_2_L2_0_G1_MINI_ALU_BoothOperand_14, 
         L1_2_L2_0_G1_MINI_ALU_BoothOperand_13, 
         L1_2_L2_0_G1_MINI_ALU_BoothOperand_12, 
         L1_2_L2_0_G1_MINI_ALU_BoothOperand_11, 
         L1_2_L2_0_G1_MINI_ALU_BoothOperand_10, 
         L1_2_L2_0_G1_MINI_ALU_BoothOperand_9, L1_2_L2_0_G1_MINI_ALU_BoothP_16, 
         L1_2_L2_0_G1_MINI_ALU_BoothP_15, L1_2_L2_0_G1_MINI_ALU_BoothP_14, 
         L1_2_L2_0_G1_MINI_ALU_BoothP_13, L1_2_L2_0_G1_MINI_ALU_BoothP_12, 
         L1_2_L2_0_G1_MINI_ALU_BoothP_11, L1_2_L2_0_G1_MINI_ALU_BoothP_10, 
         L1_2_L2_0_G1_MINI_ALU_BoothP_9, L1_2_L2_0_G1_MINI_ALU_BoothP_8, 
         L1_2_L2_0_G1_MINI_ALU_BoothP_7, L1_2_L2_0_G1_MINI_ALU_BoothP_6, 
         L1_2_L2_0_G1_MINI_ALU_BoothP_5, L1_2_L2_0_G1_MINI_ALU_BoothP_4, 
         L1_2_L2_0_G1_MINI_ALU_BoothP_3, L1_2_L2_0_G1_MINI_ALU_BoothP_2, 
         L1_2_L2_0_G1_MINI_ALU_BoothP_1, L1_2_L2_0_G1_MINI_ALU_BoothP_0, 
         L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_15, 
         L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_14, 
         L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_13, 
         L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_12, 
         L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_11, 
         L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_10, 
         L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_9, 
         L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_8, 
         L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_7, 
         L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_6, 
         L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_5, 
         L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_4, 
         L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_3, 
         L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_2, 
         L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_1, 
         L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_0, 
         L1_2_L2_1_G1_MINI_ALU_OperationResult_15, 
         L1_2_L2_1_G1_MINI_ALU_OperationResult_14, 
         L1_2_L2_1_G1_MINI_ALU_OperationResult_13, 
         L1_2_L2_1_G1_MINI_ALU_OperationResult_12, 
         L1_2_L2_1_G1_MINI_ALU_OperationResult_11, 
         L1_2_L2_1_G1_MINI_ALU_OperationResult_10, 
         L1_2_L2_1_G1_MINI_ALU_OperationResult_9, 
         L1_2_L2_1_G1_MINI_ALU_OperationResult_8, 
         L1_2_L2_1_G1_MINI_ALU_OperationResult_7, 
         L1_2_L2_1_G1_MINI_ALU_OperationResult_6, 
         L1_2_L2_1_G1_MINI_ALU_OperationResult_5, 
         L1_2_L2_1_G1_MINI_ALU_OperationResult_4, 
         L1_2_L2_1_G1_MINI_ALU_OperationResult_3, 
         L1_2_L2_1_G1_MINI_ALU_OperationResult_2, 
         L1_2_L2_1_G1_MINI_ALU_OperationResult_1, 
         L1_2_L2_1_G1_MINI_ALU_OperationResult_0, 
         L1_2_L2_1_G1_MINI_ALU_BoothXORCheck, 
         L1_2_L2_1_G1_MINI_ALU_BoothOperand_16, 
         L1_2_L2_1_G1_MINI_ALU_BoothOperand_15, 
         L1_2_L2_1_G1_MINI_ALU_BoothOperand_14, 
         L1_2_L2_1_G1_MINI_ALU_BoothOperand_13, 
         L1_2_L2_1_G1_MINI_ALU_BoothOperand_12, 
         L1_2_L2_1_G1_MINI_ALU_BoothOperand_11, 
         L1_2_L2_1_G1_MINI_ALU_BoothOperand_10, 
         L1_2_L2_1_G1_MINI_ALU_BoothOperand_9, L1_2_L2_1_G1_MINI_ALU_BoothP_16, 
         L1_2_L2_1_G1_MINI_ALU_BoothP_15, L1_2_L2_1_G1_MINI_ALU_BoothP_14, 
         L1_2_L2_1_G1_MINI_ALU_BoothP_13, L1_2_L2_1_G1_MINI_ALU_BoothP_12, 
         L1_2_L2_1_G1_MINI_ALU_BoothP_11, L1_2_L2_1_G1_MINI_ALU_BoothP_10, 
         L1_2_L2_1_G1_MINI_ALU_BoothP_9, L1_2_L2_1_G1_MINI_ALU_BoothP_8, 
         L1_2_L2_1_G1_MINI_ALU_BoothP_7, L1_2_L2_1_G1_MINI_ALU_BoothP_6, 
         L1_2_L2_1_G1_MINI_ALU_BoothP_5, L1_2_L2_1_G1_MINI_ALU_BoothP_4, 
         L1_2_L2_1_G1_MINI_ALU_BoothP_3, L1_2_L2_1_G1_MINI_ALU_BoothP_2, 
         L1_2_L2_1_G1_MINI_ALU_BoothP_1, L1_2_L2_1_G1_MINI_ALU_BoothP_0, 
         L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_15, 
         L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_14, 
         L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_13, 
         L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_12, 
         L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_11, 
         L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_10, 
         L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_9, 
         L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_8, 
         L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_7, 
         L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_6, 
         L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_5, 
         L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_4, 
         L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_3, 
         L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_2, 
         L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_1, 
         L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_0, 
         L1_2_L2_2_G1_MINI_ALU_BoothXORCheck, 
         L1_2_L2_2_G1_MINI_ALU_BoothOperand_16, 
         L1_2_L2_2_G1_MINI_ALU_BoothOperand_15, 
         L1_2_L2_2_G1_MINI_ALU_BoothOperand_14, 
         L1_2_L2_2_G1_MINI_ALU_BoothOperand_13, 
         L1_2_L2_2_G1_MINI_ALU_BoothOperand_12, 
         L1_2_L2_2_G1_MINI_ALU_BoothOperand_11, 
         L1_2_L2_2_G1_MINI_ALU_BoothOperand_10, 
         L1_2_L2_2_G1_MINI_ALU_BoothOperand_9, L1_2_L2_2_G1_MINI_ALU_BoothP_16, 
         L1_2_L2_2_G1_MINI_ALU_BoothP_15, L1_2_L2_2_G1_MINI_ALU_BoothP_14, 
         L1_2_L2_2_G1_MINI_ALU_BoothP_13, L1_2_L2_2_G1_MINI_ALU_BoothP_12, 
         L1_2_L2_2_G1_MINI_ALU_BoothP_11, L1_2_L2_2_G1_MINI_ALU_BoothP_10, 
         L1_2_L2_2_G1_MINI_ALU_BoothP_9, L1_2_L2_2_G1_MINI_ALU_BoothP_8, 
         L1_2_L2_2_G1_MINI_ALU_BoothP_7, L1_2_L2_2_G1_MINI_ALU_BoothP_6, 
         L1_2_L2_2_G1_MINI_ALU_BoothP_5, L1_2_L2_2_G1_MINI_ALU_BoothP_4, 
         L1_2_L2_2_G1_MINI_ALU_BoothP_3, L1_2_L2_2_G1_MINI_ALU_BoothP_2, 
         L1_2_L2_2_G1_MINI_ALU_BoothP_1, 
         L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_15, 
         L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_14, 
         L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_13, 
         L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_12, 
         L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_11, 
         L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_10, 
         L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_9, 
         L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_8, 
         L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_7, 
         L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_6, 
         L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_5, 
         L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_4, 
         L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_3, 
         L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_2, 
         L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_1, 
         L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_0, 
         L1_2_L2_3_G2_MINI_ALU_BoothXORCheck, 
         L1_2_L2_3_G2_MINI_ALU_BoothOperand_16, 
         L1_2_L2_3_G2_MINI_ALU_BoothOperand_15, 
         L1_2_L2_3_G2_MINI_ALU_BoothOperand_14, 
         L1_2_L2_3_G2_MINI_ALU_BoothOperand_13, 
         L1_2_L2_3_G2_MINI_ALU_BoothOperand_12, 
         L1_2_L2_3_G2_MINI_ALU_BoothOperand_11, 
         L1_2_L2_3_G2_MINI_ALU_BoothOperand_10, 
         L1_2_L2_3_G2_MINI_ALU_BoothOperand_9, L1_2_L2_3_G2_MINI_ALU_BoothP_16, 
         L1_2_L2_3_G2_MINI_ALU_BoothP_15, L1_2_L2_3_G2_MINI_ALU_BoothP_14, 
         L1_2_L2_3_G2_MINI_ALU_BoothP_13, L1_2_L2_3_G2_MINI_ALU_BoothP_12, 
         L1_2_L2_3_G2_MINI_ALU_BoothP_11, L1_2_L2_3_G2_MINI_ALU_BoothP_10, 
         L1_2_L2_3_G2_MINI_ALU_BoothP_9, L1_2_L2_3_G2_MINI_ALU_BoothP_8, 
         L1_2_L2_3_G2_MINI_ALU_BoothP_7, L1_2_L2_3_G2_MINI_ALU_BoothP_6, 
         L1_2_L2_3_G2_MINI_ALU_BoothP_5, L1_2_L2_3_G2_MINI_ALU_BoothP_4, 
         L1_2_L2_3_G2_MINI_ALU_BoothP_3, L1_2_L2_3_G2_MINI_ALU_BoothP_2, 
         L1_2_L2_3_G2_MINI_ALU_BoothP_1, L1_2_L2_3_G2_MINI_ALU_BoothP_0, 
         L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_15, 
         L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_14, 
         L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_13, 
         L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_12, 
         L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_11, 
         L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_10, 
         L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_9, 
         L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_8, 
         L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_7, 
         L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_6, 
         L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_5, 
         L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_4, 
         L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_3, 
         L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_2, 
         L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_1, 
         L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_0, 
         L1_2_L2_4_G2_MINI_ALU_BoothXORCheck, 
         L1_2_L2_4_G2_MINI_ALU_BoothOperand_16, 
         L1_2_L2_4_G2_MINI_ALU_BoothOperand_15, 
         L1_2_L2_4_G2_MINI_ALU_BoothOperand_14, 
         L1_2_L2_4_G2_MINI_ALU_BoothOperand_13, 
         L1_2_L2_4_G2_MINI_ALU_BoothOperand_12, 
         L1_2_L2_4_G2_MINI_ALU_BoothOperand_11, 
         L1_2_L2_4_G2_MINI_ALU_BoothOperand_10, 
         L1_2_L2_4_G2_MINI_ALU_BoothOperand_9, L1_2_L2_4_G2_MINI_ALU_BoothP_16, 
         L1_2_L2_4_G2_MINI_ALU_BoothP_15, L1_2_L2_4_G2_MINI_ALU_BoothP_14, 
         L1_2_L2_4_G2_MINI_ALU_BoothP_13, L1_2_L2_4_G2_MINI_ALU_BoothP_12, 
         L1_2_L2_4_G2_MINI_ALU_BoothP_11, L1_2_L2_4_G2_MINI_ALU_BoothP_10, 
         L1_2_L2_4_G2_MINI_ALU_BoothP_9, L1_2_L2_4_G2_MINI_ALU_BoothP_8, 
         L1_2_L2_4_G2_MINI_ALU_BoothP_7, L1_2_L2_4_G2_MINI_ALU_BoothP_6, 
         L1_2_L2_4_G2_MINI_ALU_BoothP_5, L1_2_L2_4_G2_MINI_ALU_BoothP_4, 
         L1_2_L2_4_G2_MINI_ALU_BoothP_3, L1_2_L2_4_G2_MINI_ALU_BoothP_2, 
         L1_2_L2_4_G2_MINI_ALU_BoothP_1, L1_2_L2_4_G2_MINI_ALU_BoothP_0, 
         L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_15, 
         L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_14, 
         L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_13, 
         L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_12, 
         L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_11, 
         L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_10, 
         L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_9, 
         L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_8, 
         L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_7, 
         L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_6, 
         L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_5, 
         L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_4, 
         L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_3, 
         L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_2, 
         L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_1, 
         L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_0, 
         L1_3_L2_0_G2_MINI_ALU_BoothXORCheck, 
         L1_3_L2_0_G2_MINI_ALU_BoothOperand_16, 
         L1_3_L2_0_G2_MINI_ALU_BoothOperand_15, 
         L1_3_L2_0_G2_MINI_ALU_BoothOperand_14, 
         L1_3_L2_0_G2_MINI_ALU_BoothOperand_13, 
         L1_3_L2_0_G2_MINI_ALU_BoothOperand_12, 
         L1_3_L2_0_G2_MINI_ALU_BoothOperand_11, 
         L1_3_L2_0_G2_MINI_ALU_BoothOperand_10, 
         L1_3_L2_0_G2_MINI_ALU_BoothOperand_9, L1_3_L2_0_G2_MINI_ALU_BoothP_16, 
         L1_3_L2_0_G2_MINI_ALU_BoothP_15, L1_3_L2_0_G2_MINI_ALU_BoothP_14, 
         L1_3_L2_0_G2_MINI_ALU_BoothP_13, L1_3_L2_0_G2_MINI_ALU_BoothP_12, 
         L1_3_L2_0_G2_MINI_ALU_BoothP_11, L1_3_L2_0_G2_MINI_ALU_BoothP_10, 
         L1_3_L2_0_G2_MINI_ALU_BoothP_9, L1_3_L2_0_G2_MINI_ALU_BoothP_8, 
         L1_3_L2_0_G2_MINI_ALU_BoothP_7, L1_3_L2_0_G2_MINI_ALU_BoothP_6, 
         L1_3_L2_0_G2_MINI_ALU_BoothP_5, L1_3_L2_0_G2_MINI_ALU_BoothP_4, 
         L1_3_L2_0_G2_MINI_ALU_BoothP_3, L1_3_L2_0_G2_MINI_ALU_BoothP_2, 
         L1_3_L2_0_G2_MINI_ALU_BoothP_1, L1_3_L2_0_G2_MINI_ALU_BoothP_0, 
         L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_15, 
         L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_14, 
         L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_13, 
         L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_12, 
         L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_11, 
         L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_10, 
         L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_9, 
         L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_8, 
         L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_7, 
         L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_6, 
         L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_5, 
         L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_4, 
         L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_3, 
         L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_2, 
         L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_1, 
         L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_0, 
         L1_3_L2_1_G2_MINI_ALU_BoothXORCheck, 
         L1_3_L2_1_G2_MINI_ALU_BoothOperand_16, 
         L1_3_L2_1_G2_MINI_ALU_BoothOperand_15, 
         L1_3_L2_1_G2_MINI_ALU_BoothOperand_14, 
         L1_3_L2_1_G2_MINI_ALU_BoothOperand_13, 
         L1_3_L2_1_G2_MINI_ALU_BoothOperand_12, 
         L1_3_L2_1_G2_MINI_ALU_BoothOperand_11, 
         L1_3_L2_1_G2_MINI_ALU_BoothOperand_10, 
         L1_3_L2_1_G2_MINI_ALU_BoothOperand_9, L1_3_L2_1_G2_MINI_ALU_BoothP_16, 
         L1_3_L2_1_G2_MINI_ALU_BoothP_15, L1_3_L2_1_G2_MINI_ALU_BoothP_14, 
         L1_3_L2_1_G2_MINI_ALU_BoothP_13, L1_3_L2_1_G2_MINI_ALU_BoothP_12, 
         L1_3_L2_1_G2_MINI_ALU_BoothP_11, L1_3_L2_1_G2_MINI_ALU_BoothP_10, 
         L1_3_L2_1_G2_MINI_ALU_BoothP_9, L1_3_L2_1_G2_MINI_ALU_BoothP_8, 
         L1_3_L2_1_G2_MINI_ALU_BoothP_7, L1_3_L2_1_G2_MINI_ALU_BoothP_6, 
         L1_3_L2_1_G2_MINI_ALU_BoothP_5, L1_3_L2_1_G2_MINI_ALU_BoothP_4, 
         L1_3_L2_1_G2_MINI_ALU_BoothP_3, L1_3_L2_1_G2_MINI_ALU_BoothP_2, 
         L1_3_L2_1_G2_MINI_ALU_BoothP_1, L1_3_L2_1_G2_MINI_ALU_BoothP_0, 
         L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_15, 
         L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_14, 
         L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_13, 
         L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_12, 
         L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_11, 
         L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_10, 
         L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_9, 
         L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_8, 
         L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_7, 
         L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_6, 
         L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_5, 
         L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_4, 
         L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_3, 
         L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_2, 
         L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_1, 
         L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_0, 
         L1_3_L2_2_G2_MINI_ALU_BoothXORCheck, 
         L1_3_L2_2_G2_MINI_ALU_BoothOperand_16, 
         L1_3_L2_2_G2_MINI_ALU_BoothOperand_15, 
         L1_3_L2_2_G2_MINI_ALU_BoothOperand_14, 
         L1_3_L2_2_G2_MINI_ALU_BoothOperand_13, 
         L1_3_L2_2_G2_MINI_ALU_BoothOperand_12, 
         L1_3_L2_2_G2_MINI_ALU_BoothOperand_11, 
         L1_3_L2_2_G2_MINI_ALU_BoothOperand_10, 
         L1_3_L2_2_G2_MINI_ALU_BoothOperand_9, L1_3_L2_2_G2_MINI_ALU_BoothP_16, 
         L1_3_L2_2_G2_MINI_ALU_BoothP_15, L1_3_L2_2_G2_MINI_ALU_BoothP_14, 
         L1_3_L2_2_G2_MINI_ALU_BoothP_13, L1_3_L2_2_G2_MINI_ALU_BoothP_12, 
         L1_3_L2_2_G2_MINI_ALU_BoothP_11, L1_3_L2_2_G2_MINI_ALU_BoothP_10, 
         L1_3_L2_2_G2_MINI_ALU_BoothP_9, L1_3_L2_2_G2_MINI_ALU_BoothP_8, 
         L1_3_L2_2_G2_MINI_ALU_BoothP_7, L1_3_L2_2_G2_MINI_ALU_BoothP_6, 
         L1_3_L2_2_G2_MINI_ALU_BoothP_5, L1_3_L2_2_G2_MINI_ALU_BoothP_4, 
         L1_3_L2_2_G2_MINI_ALU_BoothP_3, L1_3_L2_2_G2_MINI_ALU_BoothP_2, 
         L1_3_L2_2_G2_MINI_ALU_BoothP_1, L1_3_L2_2_G2_MINI_ALU_BoothP_0, 
         L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_15, 
         L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_14, 
         L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_13, 
         L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_12, 
         L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_11, 
         L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_10, 
         L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_9, 
         L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_8, 
         L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_7, 
         L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_6, 
         L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_5, 
         L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_4, 
         L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_3, 
         L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_2, 
         L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_1, 
         L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_0, 
         L1_3_L2_3_G2_MINI_ALU_BoothXORCheck, 
         L1_3_L2_3_G2_MINI_ALU_BoothOperand_16, 
         L1_3_L2_3_G2_MINI_ALU_BoothOperand_15, 
         L1_3_L2_3_G2_MINI_ALU_BoothOperand_14, 
         L1_3_L2_3_G2_MINI_ALU_BoothOperand_13, 
         L1_3_L2_3_G2_MINI_ALU_BoothOperand_12, 
         L1_3_L2_3_G2_MINI_ALU_BoothOperand_11, 
         L1_3_L2_3_G2_MINI_ALU_BoothOperand_10, 
         L1_3_L2_3_G2_MINI_ALU_BoothOperand_9, L1_3_L2_3_G2_MINI_ALU_BoothP_16, 
         L1_3_L2_3_G2_MINI_ALU_BoothP_15, L1_3_L2_3_G2_MINI_ALU_BoothP_14, 
         L1_3_L2_3_G2_MINI_ALU_BoothP_13, L1_3_L2_3_G2_MINI_ALU_BoothP_12, 
         L1_3_L2_3_G2_MINI_ALU_BoothP_11, L1_3_L2_3_G2_MINI_ALU_BoothP_10, 
         L1_3_L2_3_G2_MINI_ALU_BoothP_9, L1_3_L2_3_G2_MINI_ALU_BoothP_8, 
         L1_3_L2_3_G2_MINI_ALU_BoothP_7, L1_3_L2_3_G2_MINI_ALU_BoothP_6, 
         L1_3_L2_3_G2_MINI_ALU_BoothP_5, L1_3_L2_3_G2_MINI_ALU_BoothP_4, 
         L1_3_L2_3_G2_MINI_ALU_BoothP_3, L1_3_L2_3_G2_MINI_ALU_BoothP_2, 
         L1_3_L2_3_G2_MINI_ALU_BoothP_1, L1_3_L2_3_G2_MINI_ALU_BoothP_0, 
         L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_15, 
         L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_14, 
         L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_13, 
         L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_12, 
         L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_11, 
         L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_10, 
         L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_9, 
         L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_8, 
         L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_7, 
         L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_6, 
         L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_5, 
         L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_4, 
         L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_3, 
         L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_2, 
         L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_1, 
         L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_0, 
         L1_3_L2_4_G3_MINI_ALU_BoothXORCheck, 
         L1_3_L2_4_G3_MINI_ALU_BoothOperand_16, 
         L1_3_L2_4_G3_MINI_ALU_BoothOperand_15, 
         L1_3_L2_4_G3_MINI_ALU_BoothOperand_14, 
         L1_3_L2_4_G3_MINI_ALU_BoothOperand_13, 
         L1_3_L2_4_G3_MINI_ALU_BoothOperand_12, 
         L1_3_L2_4_G3_MINI_ALU_BoothOperand_11, 
         L1_3_L2_4_G3_MINI_ALU_BoothOperand_10, 
         L1_3_L2_4_G3_MINI_ALU_BoothOperand_9, L1_3_L2_4_G3_MINI_ALU_BoothP_16, 
         L1_3_L2_4_G3_MINI_ALU_BoothP_15, L1_3_L2_4_G3_MINI_ALU_BoothP_14, 
         L1_3_L2_4_G3_MINI_ALU_BoothP_13, L1_3_L2_4_G3_MINI_ALU_BoothP_12, 
         L1_3_L2_4_G3_MINI_ALU_BoothP_11, L1_3_L2_4_G3_MINI_ALU_BoothP_10, 
         L1_3_L2_4_G3_MINI_ALU_BoothP_9, L1_3_L2_4_G3_MINI_ALU_BoothP_8, 
         L1_3_L2_4_G3_MINI_ALU_BoothP_7, L1_3_L2_4_G3_MINI_ALU_BoothP_6, 
         L1_3_L2_4_G3_MINI_ALU_BoothP_5, L1_3_L2_4_G3_MINI_ALU_BoothP_4, 
         L1_3_L2_4_G3_MINI_ALU_BoothP_3, L1_3_L2_4_G3_MINI_ALU_BoothP_2, 
         L1_3_L2_4_G3_MINI_ALU_BoothP_1, L1_3_L2_4_G3_MINI_ALU_BoothP_0, 
         L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_15, 
         L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_14, 
         L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_13, 
         L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_12, 
         L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_11, 
         L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_10, 
         L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_9, 
         L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_8, 
         L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_7, 
         L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_6, 
         L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_5, 
         L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_4, 
         L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_3, 
         L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_2, 
         L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_1, 
         L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_0, 
         L1_4_L2_0_G3_MINI_ALU_BoothXORCheck, 
         L1_4_L2_0_G3_MINI_ALU_BoothOperand_16, 
         L1_4_L2_0_G3_MINI_ALU_BoothOperand_15, 
         L1_4_L2_0_G3_MINI_ALU_BoothOperand_14, 
         L1_4_L2_0_G3_MINI_ALU_BoothOperand_13, 
         L1_4_L2_0_G3_MINI_ALU_BoothOperand_12, 
         L1_4_L2_0_G3_MINI_ALU_BoothOperand_11, 
         L1_4_L2_0_G3_MINI_ALU_BoothOperand_10, 
         L1_4_L2_0_G3_MINI_ALU_BoothOperand_9, L1_4_L2_0_G3_MINI_ALU_BoothP_16, 
         L1_4_L2_0_G3_MINI_ALU_BoothP_15, L1_4_L2_0_G3_MINI_ALU_BoothP_14, 
         L1_4_L2_0_G3_MINI_ALU_BoothP_13, L1_4_L2_0_G3_MINI_ALU_BoothP_12, 
         L1_4_L2_0_G3_MINI_ALU_BoothP_11, L1_4_L2_0_G3_MINI_ALU_BoothP_10, 
         L1_4_L2_0_G3_MINI_ALU_BoothP_9, L1_4_L2_0_G3_MINI_ALU_BoothP_8, 
         L1_4_L2_0_G3_MINI_ALU_BoothP_7, L1_4_L2_0_G3_MINI_ALU_BoothP_6, 
         L1_4_L2_0_G3_MINI_ALU_BoothP_5, L1_4_L2_0_G3_MINI_ALU_BoothP_4, 
         L1_4_L2_0_G3_MINI_ALU_BoothP_3, L1_4_L2_0_G3_MINI_ALU_BoothP_2, 
         L1_4_L2_0_G3_MINI_ALU_BoothP_1, L1_4_L2_0_G3_MINI_ALU_BoothP_0, 
         L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_15, 
         L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_14, 
         L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_13, 
         L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_12, 
         L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_11, 
         L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_10, 
         L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_9, 
         L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_8, 
         L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_7, 
         L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_6, 
         L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_5, 
         L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_4, 
         L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_3, 
         L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_2, 
         L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_1, 
         L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_0, 
         L1_4_L2_1_G3_MINI_ALU_BoothXORCheck, 
         L1_4_L2_1_G3_MINI_ALU_BoothOperand_16, 
         L1_4_L2_1_G3_MINI_ALU_BoothOperand_15, 
         L1_4_L2_1_G3_MINI_ALU_BoothOperand_14, 
         L1_4_L2_1_G3_MINI_ALU_BoothOperand_13, 
         L1_4_L2_1_G3_MINI_ALU_BoothOperand_12, 
         L1_4_L2_1_G3_MINI_ALU_BoothOperand_11, 
         L1_4_L2_1_G3_MINI_ALU_BoothOperand_10, 
         L1_4_L2_1_G3_MINI_ALU_BoothOperand_9, L1_4_L2_1_G3_MINI_ALU_BoothP_16, 
         L1_4_L2_1_G3_MINI_ALU_BoothP_15, L1_4_L2_1_G3_MINI_ALU_BoothP_14, 
         L1_4_L2_1_G3_MINI_ALU_BoothP_13, L1_4_L2_1_G3_MINI_ALU_BoothP_12, 
         L1_4_L2_1_G3_MINI_ALU_BoothP_11, L1_4_L2_1_G3_MINI_ALU_BoothP_10, 
         L1_4_L2_1_G3_MINI_ALU_BoothP_9, L1_4_L2_1_G3_MINI_ALU_BoothP_8, 
         L1_4_L2_1_G3_MINI_ALU_BoothP_7, L1_4_L2_1_G3_MINI_ALU_BoothP_6, 
         L1_4_L2_1_G3_MINI_ALU_BoothP_5, L1_4_L2_1_G3_MINI_ALU_BoothP_4, 
         L1_4_L2_1_G3_MINI_ALU_BoothP_3, L1_4_L2_1_G3_MINI_ALU_BoothP_2, 
         L1_4_L2_1_G3_MINI_ALU_BoothP_1, L1_4_L2_1_G3_MINI_ALU_BoothP_0, 
         L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_15, 
         L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_14, 
         L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_13, 
         L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_12, 
         L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_11, 
         L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_10, 
         L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_9, 
         L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_8, 
         L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_7, 
         L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_6, 
         L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_5, 
         L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_4, 
         L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_3, 
         L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_2, 
         L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_1, 
         L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_0, 
         L1_4_L2_2_G4_MINI_ALU_BoothXORCheck, 
         L1_4_L2_2_G4_MINI_ALU_BoothOperand_16, 
         L1_4_L2_2_G4_MINI_ALU_BoothOperand_15, 
         L1_4_L2_2_G4_MINI_ALU_BoothOperand_14, 
         L1_4_L2_2_G4_MINI_ALU_BoothOperand_13, 
         L1_4_L2_2_G4_MINI_ALU_BoothOperand_12, 
         L1_4_L2_2_G4_MINI_ALU_BoothOperand_11, 
         L1_4_L2_2_G4_MINI_ALU_BoothOperand_10, 
         L1_4_L2_2_G4_MINI_ALU_BoothOperand_9, L1_4_L2_2_G4_MINI_ALU_BoothP_16, 
         L1_4_L2_2_G4_MINI_ALU_BoothP_15, L1_4_L2_2_G4_MINI_ALU_BoothP_14, 
         L1_4_L2_2_G4_MINI_ALU_BoothP_13, L1_4_L2_2_G4_MINI_ALU_BoothP_12, 
         L1_4_L2_2_G4_MINI_ALU_BoothP_11, L1_4_L2_2_G4_MINI_ALU_BoothP_10, 
         L1_4_L2_2_G4_MINI_ALU_BoothP_9, L1_4_L2_2_G4_MINI_ALU_BoothP_8, 
         L1_4_L2_2_G4_MINI_ALU_BoothP_7, L1_4_L2_2_G4_MINI_ALU_BoothP_6, 
         L1_4_L2_2_G4_MINI_ALU_BoothP_5, L1_4_L2_2_G4_MINI_ALU_BoothP_4, 
         L1_4_L2_2_G4_MINI_ALU_BoothP_3, L1_4_L2_2_G4_MINI_ALU_BoothP_2, 
         L1_4_L2_2_G4_MINI_ALU_BoothP_1, L1_4_L2_2_G4_MINI_ALU_BoothP_0, 
         L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_15, 
         L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_14, 
         L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_13, 
         L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_12, 
         L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_11, 
         L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_10, 
         L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_9, 
         L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_8, 
         L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_7, 
         L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_6, 
         L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_5, 
         L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_4, 
         L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_3, 
         L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_2, 
         L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_1, 
         L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_0, 
         L1_4_L2_3_G5_MINI_ALU_BoothXORCheck, 
         L1_4_L2_3_G5_MINI_ALU_BoothOperand_16, 
         L1_4_L2_3_G5_MINI_ALU_BoothOperand_15, 
         L1_4_L2_3_G5_MINI_ALU_BoothOperand_14, 
         L1_4_L2_3_G5_MINI_ALU_BoothOperand_13, 
         L1_4_L2_3_G5_MINI_ALU_BoothOperand_12, 
         L1_4_L2_3_G5_MINI_ALU_BoothOperand_11, 
         L1_4_L2_3_G5_MINI_ALU_BoothOperand_10, 
         L1_4_L2_3_G5_MINI_ALU_BoothOperand_9, L1_4_L2_3_G5_MINI_ALU_BoothP_16, 
         L1_4_L2_3_G5_MINI_ALU_BoothP_15, L1_4_L2_3_G5_MINI_ALU_BoothP_14, 
         L1_4_L2_3_G5_MINI_ALU_BoothP_13, L1_4_L2_3_G5_MINI_ALU_BoothP_12, 
         L1_4_L2_3_G5_MINI_ALU_BoothP_11, L1_4_L2_3_G5_MINI_ALU_BoothP_10, 
         L1_4_L2_3_G5_MINI_ALU_BoothP_9, L1_4_L2_3_G5_MINI_ALU_BoothP_8, 
         L1_4_L2_3_G5_MINI_ALU_BoothP_7, L1_4_L2_3_G5_MINI_ALU_BoothP_6, 
         L1_4_L2_3_G5_MINI_ALU_BoothP_5, L1_4_L2_3_G5_MINI_ALU_BoothP_4, 
         L1_4_L2_3_G5_MINI_ALU_BoothP_3, L1_4_L2_3_G5_MINI_ALU_BoothP_2, 
         L1_4_L2_3_G5_MINI_ALU_BoothP_1, L1_4_L2_3_G5_MINI_ALU_BoothP_0, 
         L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_15, 
         L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_14, 
         L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_13, 
         L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_12, 
         L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_11, 
         L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_10, 
         L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_9, 
         L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_8, 
         L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_7, 
         L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_6, 
         L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_5, 
         L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_4, 
         L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_3, 
         L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_2, 
         L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_1, 
         L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_0, 
         L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_7, 
         L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_6, 
         L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_5, 
         L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_4, 
         L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_3, 
         L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_2, 
         L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_1, 
         L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_0, 
         L1_4_L2_4_G5_MINI_ALU_OperationResult_15, 
         L1_4_L2_4_G5_MINI_ALU_OperationResult_14, 
         L1_4_L2_4_G5_MINI_ALU_OperationResult_13, 
         L1_4_L2_4_G5_MINI_ALU_OperationResult_12, 
         L1_4_L2_4_G5_MINI_ALU_OperationResult_11, 
         L1_4_L2_4_G5_MINI_ALU_OperationResult_10, 
         L1_4_L2_4_G5_MINI_ALU_OperationResult_9, 
         L1_4_L2_4_G5_MINI_ALU_OperationResult_8, 
         L1_4_L2_4_G5_MINI_ALU_OperationResult_7, 
         L1_4_L2_4_G5_MINI_ALU_OperationResult_6, 
         L1_4_L2_4_G5_MINI_ALU_OperationResult_5, 
         L1_4_L2_4_G5_MINI_ALU_OperationResult_4, 
         L1_4_L2_4_G5_MINI_ALU_OperationResult_3, 
         L1_4_L2_4_G5_MINI_ALU_OperationResult_2, 
         L1_4_L2_4_G5_MINI_ALU_OperationResult_1, 
         L1_4_L2_4_G5_MINI_ALU_OperationResult_0, 
         L1_4_L2_4_G5_MINI_ALU_BoothXORCheck, 
         L1_4_L2_4_G5_MINI_ALU_BoothOperand_16, 
         L1_4_L2_4_G5_MINI_ALU_BoothOperand_15, 
         L1_4_L2_4_G5_MINI_ALU_BoothOperand_14, 
         L1_4_L2_4_G5_MINI_ALU_BoothOperand_13, 
         L1_4_L2_4_G5_MINI_ALU_BoothOperand_12, 
         L1_4_L2_4_G5_MINI_ALU_BoothOperand_11, 
         L1_4_L2_4_G5_MINI_ALU_BoothOperand_10, 
         L1_4_L2_4_G5_MINI_ALU_BoothOperand_9, L1_4_L2_4_G5_MINI_ALU_BoothP_16, 
         L1_4_L2_4_G5_MINI_ALU_BoothP_15, L1_4_L2_4_G5_MINI_ALU_BoothP_14, 
         L1_4_L2_4_G5_MINI_ALU_BoothP_13, L1_4_L2_4_G5_MINI_ALU_BoothP_12, 
         L1_4_L2_4_G5_MINI_ALU_BoothP_11, L1_4_L2_4_G5_MINI_ALU_BoothP_10, 
         L1_4_L2_4_G5_MINI_ALU_BoothP_9, L1_4_L2_4_G5_MINI_ALU_BoothP_8, 
         L1_4_L2_4_G5_MINI_ALU_BoothP_7, L1_4_L2_4_G5_MINI_ALU_BoothP_6, 
         L1_4_L2_4_G5_MINI_ALU_BoothP_5, L1_4_L2_4_G5_MINI_ALU_BoothP_4, 
         L1_4_L2_4_G5_MINI_ALU_BoothP_3, L1_4_L2_4_G5_MINI_ALU_BoothP_2, 
         L1_4_L2_4_G5_MINI_ALU_BoothP_1, L1_4_L2_4_G5_MINI_ALU_BoothP_0, 
         L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_15, 
         L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_14, 
         L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_13, 
         L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_12, 
         L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_11, 
         L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_10, 
         L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_9, 
         L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_8, 
         L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_7, 
         L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_6, 
         L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_5, 
         L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_4, 
         L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_3, 
         L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_2, 
         L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_1, 
         L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_0, L1FirstOperands_12__16, nx22, 
         CounterOut_0, NOT__145383, nx1032, NOT_CounterOut_0, nx1036, 
         CounterOut_3, CounterOut_2, CounterOut_1, nx1046, nx1058, nx1066, 
         nx2853, nx2865, nx2869, nx2873, nx3230, nx3233, nx3235, nx3239, nx3241, 
         nx3244, nx3246, nx3270, nx3272, nx3274, nx3276, nx3278, nx3280, nx3282, 
         nx3284, nx3286, nx3292;
    wire [903:0] \$dummy ;




    booth_adder_17 L1_0_L2_0_G1_MINI_ALU_BOOTH_ADDER (.AdderFirstOperand ({
                   L1FirstOperands_12__16,L1FirstOperands_0__15,
                   L1FirstOperands_0__14,L1FirstOperands_0__13,
                   L1FirstOperands_0__12,L1FirstOperands_0__11,
                   L1FirstOperands_0__10,L1FirstOperands_0__9,
                   L1FirstOperands_0__8,L1FirstOperands_0__7,
                   L1FirstOperands_0__6,L1FirstOperands_0__5,
                   L1FirstOperands_0__4,L1FirstOperands_0__3,
                   L1FirstOperands_0__2,L1FirstOperands_0__1,
                   L1FirstOperands_0__0}), .AdderSecondOperand ({
                   L1FirstOperands_12__16,
                   L1_0_L2_0_G1_MINI_ALU_OperationResult_15,
                   L1_0_L2_0_G1_MINI_ALU_OperationResult_14,
                   L1_0_L2_0_G1_MINI_ALU_OperationResult_13,
                   L1_0_L2_0_G1_MINI_ALU_OperationResult_12,
                   L1_0_L2_0_G1_MINI_ALU_OperationResult_11,
                   L1_0_L2_0_G1_MINI_ALU_OperationResult_10,
                   L1_0_L2_0_G1_MINI_ALU_OperationResult_9,
                   L1_0_L2_0_G1_MINI_ALU_OperationResult_8,
                   L1_0_L2_0_G1_MINI_ALU_OperationResult_7,
                   L1_0_L2_0_G1_MINI_ALU_OperationResult_6,
                   L1_0_L2_0_G1_MINI_ALU_OperationResult_5,
                   L1_0_L2_0_G1_MINI_ALU_OperationResult_4,
                   L1_0_L2_0_G1_MINI_ALU_OperationResult_3,
                   L1_0_L2_0_G1_MINI_ALU_OperationResult_2,
                   L1_0_L2_0_G1_MINI_ALU_OperationResult_1,
                   L1_0_L2_0_G1_MINI_ALU_OperationResult_0}), .BoothOperand ({
                   L1_0_L2_0_G1_MINI_ALU_BoothOperand_16,
                   L1_0_L2_0_G1_MINI_ALU_BoothOperand_15,
                   L1_0_L2_0_G1_MINI_ALU_BoothOperand_14,
                   L1_0_L2_0_G1_MINI_ALU_BoothOperand_13,
                   L1_0_L2_0_G1_MINI_ALU_BoothOperand_12,
                   L1_0_L2_0_G1_MINI_ALU_BoothOperand_11,
                   L1_0_L2_0_G1_MINI_ALU_BoothOperand_10,
                   L1_0_L2_0_G1_MINI_ALU_BoothOperand_9,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16}), .BoothP ({
                   L1_0_L2_0_G1_MINI_ALU_BoothP_16,
                   L1_0_L2_0_G1_MINI_ALU_BoothP_15,
                   L1_0_L2_0_G1_MINI_ALU_BoothP_14,
                   L1_0_L2_0_G1_MINI_ALU_BoothP_13,
                   L1_0_L2_0_G1_MINI_ALU_BoothP_12,
                   L1_0_L2_0_G1_MINI_ALU_BoothP_11,
                   L1_0_L2_0_G1_MINI_ALU_BoothP_10,
                   L1_0_L2_0_G1_MINI_ALU_BoothP_9,L1_0_L2_0_G1_MINI_ALU_BoothP_8
                   ,L1_0_L2_0_G1_MINI_ALU_BoothP_7,
                   L1_0_L2_0_G1_MINI_ALU_BoothP_6,L1_0_L2_0_G1_MINI_ALU_BoothP_5
                   ,L1_0_L2_0_G1_MINI_ALU_BoothP_4,
                   L1_0_L2_0_G1_MINI_ALU_BoothP_3,L1_0_L2_0_G1_MINI_ALU_BoothP_2
                   ,L1_0_L2_0_G1_MINI_ALU_BoothP_1,
                   L1_0_L2_0_G1_MINI_ALU_BoothP_0}), .SelOperand (nx3282), .Operation (
                   L1_0_L2_0_G1_MINI_ALU_BoothXORCheck), .AdderResult ({
                   L1ResultsLarge_0__16,L1ResultsLarge_0__15,
                   L1ResultsLarge_0__14,L1ResultsLarge_0__13,
                   L1ResultsLarge_0__12,L1ResultsLarge_0__11,
                   L1ResultsLarge_0__10,L1ResultsLarge_0__9,L1ResultsLarge_0__8,
                   L1ResultsLarge_0__7,L1ResultsLarge_0__6,L1ResultsLarge_0__5,
                   L1ResultsLarge_0__4,L1ResultsLarge_0__3,L1ResultsLarge_0__2,
                   L1ResultsLarge_0__1,L1ResultsLarge_0__0}), .AdderBoothResult (
                   {\$dummy [0],L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_15,
                   L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_14,
                   L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_13,
                   L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_12,
                   L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_11,
                   L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_10,
                   L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_9,
                   L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_8,
                   L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_7,
                   L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_6,
                   L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_5,
                   L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_4,
                   L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_3,
                   L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_2,
                   L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_1,
                   L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_0})) ;
    booth_unit_17 L1_0_L2_0_G1_MINI_ALU_BOOTH_UNIT (.CLK (CLK), .RST (RST), .Start (
                  Start), .Instr (Instr), .LoopingAndResultNotReady (nx3272), .Filter (
                  {FilterDin_0__0__7,FilterDin_0__0__6,FilterDin_0__0__5,
                  FilterDin_0__0__4,FilterDin_0__0__3,FilterDin_0__0__2,
                  FilterDin_0__0__1,FilterDin_0__0__0}), .Window ({
                  WindowDin_0__0__7,WindowDin_0__0__6,WindowDin_0__0__5,
                  WindowDin_0__0__4,WindowDin_0__0__3,WindowDin_0__0__2,
                  WindowDin_0__0__1,WindowDin_0__0__0}), .AdderBoothResult ({
                  L1FirstOperands_12__16,
                  L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_15,
                  L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_14,
                  L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_13,
                  L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_12,
                  L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_11,
                  L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_10,
                  L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_9,
                  L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_8,
                  L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_7,
                  L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_6,
                  L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_5,
                  L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_4,
                  L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_3,
                  L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_2,
                  L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_1,
                  L1_0_L2_0_G1_MINI_ALU_AdderBoothResult_0}), .BoothXORCheck (
                  L1_0_L2_0_G1_MINI_ALU_BoothXORCheck), .BoothResult ({
                  \$dummy [1],\$dummy [2],\$dummy [3],\$dummy [4],\$dummy [5],
                  \$dummy [6],\$dummy [7],\$dummy [8]}), .BoothAddingOperand ({
                  L1_0_L2_0_G1_MINI_ALU_BoothOperand_16,
                  L1_0_L2_0_G1_MINI_ALU_BoothOperand_15,
                  L1_0_L2_0_G1_MINI_ALU_BoothOperand_14,
                  L1_0_L2_0_G1_MINI_ALU_BoothOperand_13,
                  L1_0_L2_0_G1_MINI_ALU_BoothOperand_12,
                  L1_0_L2_0_G1_MINI_ALU_BoothOperand_11,
                  L1_0_L2_0_G1_MINI_ALU_BoothOperand_10,
                  L1_0_L2_0_G1_MINI_ALU_BoothOperand_9,\$dummy [9],\$dummy [10],
                  \$dummy [11],\$dummy [12],\$dummy [13],\$dummy [14],
                  \$dummy [15],\$dummy [16],\$dummy [17]}), .BoothP ({
                  L1_0_L2_0_G1_MINI_ALU_BoothP_16,
                  L1_0_L2_0_G1_MINI_ALU_BoothP_15,
                  L1_0_L2_0_G1_MINI_ALU_BoothP_14,
                  L1_0_L2_0_G1_MINI_ALU_BoothP_13,
                  L1_0_L2_0_G1_MINI_ALU_BoothP_12,
                  L1_0_L2_0_G1_MINI_ALU_BoothP_11,
                  L1_0_L2_0_G1_MINI_ALU_BoothP_10,L1_0_L2_0_G1_MINI_ALU_BoothP_9
                  ,L1_0_L2_0_G1_MINI_ALU_BoothP_8,L1_0_L2_0_G1_MINI_ALU_BoothP_7
                  ,L1_0_L2_0_G1_MINI_ALU_BoothP_6,L1_0_L2_0_G1_MINI_ALU_BoothP_5
                  ,L1_0_L2_0_G1_MINI_ALU_BoothP_4,L1_0_L2_0_G1_MINI_ALU_BoothP_3
                  ,L1_0_L2_0_G1_MINI_ALU_BoothP_2,L1_0_L2_0_G1_MINI_ALU_BoothP_1
                  ,L1_0_L2_0_G1_MINI_ALU_BoothP_0}), .LargeWindowShifted ({
                  \$dummy [18],\$dummy [19],\$dummy [20],\$dummy [21],
                  \$dummy [22],\$dummy [23],\$dummy [24],\$dummy [25],
                  \$dummy [26],\$dummy [27],\$dummy [28],\$dummy [29],
                  \$dummy [30],\$dummy [31],\$dummy [32],\$dummy [33],
                  \$dummy [34]})) ;
    booth_adder_17 L1_0_L2_1_G1_MINI_ALU_BOOTH_ADDER (.AdderFirstOperand ({
                   L1FirstOperands_12__16,L1FirstOperands_0__15,
                   L1FirstOperands_0__14,L1FirstOperands_0__13,
                   L1FirstOperands_0__12,L1FirstOperands_0__11,
                   L1FirstOperands_0__10,L1FirstOperands_0__9,
                   L1FirstOperands_0__8,L1FirstOperands_0__7,
                   L1FirstOperands_0__6,L1FirstOperands_0__5,
                   L1FirstOperands_0__4,L1FirstOperands_0__3,
                   L1FirstOperands_0__2,L1FirstOperands_0__1,
                   L1FirstOperands_0__0}), .AdderSecondOperand ({
                   L1FirstOperands_12__16,
                   L1_0_L2_1_G1_MINI_ALU_OperationResult_15,
                   L1_0_L2_1_G1_MINI_ALU_OperationResult_14,
                   L1_0_L2_1_G1_MINI_ALU_OperationResult_13,
                   L1_0_L2_1_G1_MINI_ALU_OperationResult_12,
                   L1_0_L2_1_G1_MINI_ALU_OperationResult_11,
                   L1_0_L2_1_G1_MINI_ALU_OperationResult_10,
                   L1_0_L2_1_G1_MINI_ALU_OperationResult_9,
                   L1_0_L2_1_G1_MINI_ALU_OperationResult_8,
                   L1_0_L2_1_G1_MINI_ALU_OperationResult_7,
                   L1_0_L2_1_G1_MINI_ALU_OperationResult_6,
                   L1_0_L2_1_G1_MINI_ALU_OperationResult_5,
                   L1_0_L2_1_G1_MINI_ALU_OperationResult_4,
                   L1_0_L2_1_G1_MINI_ALU_OperationResult_3,
                   L1_0_L2_1_G1_MINI_ALU_OperationResult_2,
                   L1_0_L2_1_G1_MINI_ALU_OperationResult_1,
                   L1_0_L2_1_G1_MINI_ALU_OperationResult_0}), .BoothOperand ({
                   L1_0_L2_1_G1_MINI_ALU_BoothOperand_16,
                   L1_0_L2_1_G1_MINI_ALU_BoothOperand_15,
                   L1_0_L2_1_G1_MINI_ALU_BoothOperand_14,
                   L1_0_L2_1_G1_MINI_ALU_BoothOperand_13,
                   L1_0_L2_1_G1_MINI_ALU_BoothOperand_12,
                   L1_0_L2_1_G1_MINI_ALU_BoothOperand_11,
                   L1_0_L2_1_G1_MINI_ALU_BoothOperand_10,
                   L1_0_L2_1_G1_MINI_ALU_BoothOperand_9,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16}), .BoothP ({
                   L1_0_L2_1_G1_MINI_ALU_BoothP_16,
                   L1_0_L2_1_G1_MINI_ALU_BoothP_15,
                   L1_0_L2_1_G1_MINI_ALU_BoothP_14,
                   L1_0_L2_1_G1_MINI_ALU_BoothP_13,
                   L1_0_L2_1_G1_MINI_ALU_BoothP_12,
                   L1_0_L2_1_G1_MINI_ALU_BoothP_11,
                   L1_0_L2_1_G1_MINI_ALU_BoothP_10,
                   L1_0_L2_1_G1_MINI_ALU_BoothP_9,L1_0_L2_1_G1_MINI_ALU_BoothP_8
                   ,L1_0_L2_1_G1_MINI_ALU_BoothP_7,
                   L1_0_L2_1_G1_MINI_ALU_BoothP_6,L1_0_L2_1_G1_MINI_ALU_BoothP_5
                   ,L1_0_L2_1_G1_MINI_ALU_BoothP_4,
                   L1_0_L2_1_G1_MINI_ALU_BoothP_3,L1_0_L2_1_G1_MINI_ALU_BoothP_2
                   ,L1_0_L2_1_G1_MINI_ALU_BoothP_1,
                   L1_0_L2_1_G1_MINI_ALU_BoothP_0}), .SelOperand (nx3282), .Operation (
                   L1_0_L2_1_G1_MINI_ALU_BoothXORCheck), .AdderResult ({
                   L1ResultsLarge_1__16,L1ResultsLarge_1__15,
                   L1ResultsLarge_1__14,L1ResultsLarge_1__13,
                   L1ResultsLarge_1__12,L1ResultsLarge_1__11,
                   L1ResultsLarge_1__10,L1ResultsLarge_1__9,L1ResultsLarge_1__8,
                   L1ResultsLarge_1__7,L1ResultsLarge_1__6,L1ResultsLarge_1__5,
                   L1ResultsLarge_1__4,L1ResultsLarge_1__3,L1ResultsLarge_1__2,
                   L1ResultsLarge_1__1,L1ResultsLarge_1__0}), .AdderBoothResult (
                   {\$dummy [35],L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_15,
                   L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_14,
                   L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_13,
                   L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_12,
                   L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_11,
                   L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_10,
                   L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_9,
                   L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_8,
                   L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_7,
                   L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_6,
                   L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_5,
                   L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_4,
                   L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_3,
                   L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_2,
                   L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_1,
                   L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_0})) ;
    booth_unit_17 L1_0_L2_1_G1_MINI_ALU_BOOTH_UNIT (.CLK (CLK), .RST (RST), .Start (
                  Start), .Instr (Instr), .LoopingAndResultNotReady (nx3272), .Filter (
                  {FilterDin_0__1__7,FilterDin_0__1__6,FilterDin_0__1__5,
                  FilterDin_0__1__4,FilterDin_0__1__3,FilterDin_0__1__2,
                  FilterDin_0__1__1,FilterDin_0__1__0}), .Window ({
                  WindowDin_0__1__7,WindowDin_0__1__6,WindowDin_0__1__5,
                  WindowDin_0__1__4,WindowDin_0__1__3,WindowDin_0__1__2,
                  WindowDin_0__1__1,WindowDin_0__1__0}), .AdderBoothResult ({
                  L1FirstOperands_12__16,
                  L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_15,
                  L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_14,
                  L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_13,
                  L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_12,
                  L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_11,
                  L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_10,
                  L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_9,
                  L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_8,
                  L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_7,
                  L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_6,
                  L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_5,
                  L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_4,
                  L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_3,
                  L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_2,
                  L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_1,
                  L1_0_L2_1_G1_MINI_ALU_AdderBoothResult_0}), .BoothXORCheck (
                  L1_0_L2_1_G1_MINI_ALU_BoothXORCheck), .BoothResult ({
                  \$dummy [36],\$dummy [37],\$dummy [38],\$dummy [39],
                  \$dummy [40],\$dummy [41],\$dummy [42],\$dummy [43]}), .BoothAddingOperand (
                  {L1_0_L2_1_G1_MINI_ALU_BoothOperand_16,
                  L1_0_L2_1_G1_MINI_ALU_BoothOperand_15,
                  L1_0_L2_1_G1_MINI_ALU_BoothOperand_14,
                  L1_0_L2_1_G1_MINI_ALU_BoothOperand_13,
                  L1_0_L2_1_G1_MINI_ALU_BoothOperand_12,
                  L1_0_L2_1_G1_MINI_ALU_BoothOperand_11,
                  L1_0_L2_1_G1_MINI_ALU_BoothOperand_10,
                  L1_0_L2_1_G1_MINI_ALU_BoothOperand_9,\$dummy [44],\$dummy [45]
                  ,\$dummy [46],\$dummy [47],\$dummy [48],\$dummy [49],
                  \$dummy [50],\$dummy [51],\$dummy [52]}), .BoothP ({
                  L1_0_L2_1_G1_MINI_ALU_BoothP_16,
                  L1_0_L2_1_G1_MINI_ALU_BoothP_15,
                  L1_0_L2_1_G1_MINI_ALU_BoothP_14,
                  L1_0_L2_1_G1_MINI_ALU_BoothP_13,
                  L1_0_L2_1_G1_MINI_ALU_BoothP_12,
                  L1_0_L2_1_G1_MINI_ALU_BoothP_11,
                  L1_0_L2_1_G1_MINI_ALU_BoothP_10,L1_0_L2_1_G1_MINI_ALU_BoothP_9
                  ,L1_0_L2_1_G1_MINI_ALU_BoothP_8,L1_0_L2_1_G1_MINI_ALU_BoothP_7
                  ,L1_0_L2_1_G1_MINI_ALU_BoothP_6,L1_0_L2_1_G1_MINI_ALU_BoothP_5
                  ,L1_0_L2_1_G1_MINI_ALU_BoothP_4,L1_0_L2_1_G1_MINI_ALU_BoothP_3
                  ,L1_0_L2_1_G1_MINI_ALU_BoothP_2,L1_0_L2_1_G1_MINI_ALU_BoothP_1
                  ,L1_0_L2_1_G1_MINI_ALU_BoothP_0}), .LargeWindowShifted ({
                  \$dummy [53],\$dummy [54],\$dummy [55],\$dummy [56],
                  \$dummy [57],\$dummy [58],\$dummy [59],\$dummy [60],
                  \$dummy [61],\$dummy [62],\$dummy [63],\$dummy [64],
                  \$dummy [65],\$dummy [66],\$dummy [67],\$dummy [68],
                  \$dummy [69]})) ;
    booth_adder_17 L1_0_L2_2_G1_MINI_ALU_BOOTH_ADDER (.AdderFirstOperand ({
                   L1FirstOperands_12__16,L1FirstOperands_2__15,
                   L1FirstOperands_2__14,L1FirstOperands_2__13,
                   L1FirstOperands_2__12,L1FirstOperands_2__11,
                   L1FirstOperands_2__10,L1FirstOperands_2__9,
                   L1FirstOperands_2__8,L1FirstOperands_2__7,
                   L1FirstOperands_2__6,L1FirstOperands_2__5,
                   L1FirstOperands_2__4,L1FirstOperands_2__3,
                   L1FirstOperands_2__2,L1FirstOperands_2__1,
                   L1FirstOperands_2__0}), .AdderSecondOperand ({
                   L1FirstOperands_12__16,
                   L1_0_L2_2_G1_MINI_ALU_OperationResult_15,
                   L1_0_L2_2_G1_MINI_ALU_OperationResult_14,
                   L1_0_L2_2_G1_MINI_ALU_OperationResult_13,
                   L1_0_L2_2_G1_MINI_ALU_OperationResult_12,
                   L1_0_L2_2_G1_MINI_ALU_OperationResult_11,
                   L1_0_L2_2_G1_MINI_ALU_OperationResult_10,
                   L1_0_L2_2_G1_MINI_ALU_OperationResult_9,
                   L1_0_L2_2_G1_MINI_ALU_OperationResult_8,
                   L1_0_L2_2_G1_MINI_ALU_OperationResult_7,
                   L1_0_L2_2_G1_MINI_ALU_OperationResult_6,
                   L1_0_L2_2_G1_MINI_ALU_OperationResult_5,
                   L1_0_L2_2_G1_MINI_ALU_OperationResult_4,
                   L1_0_L2_2_G1_MINI_ALU_OperationResult_3,
                   L1_0_L2_2_G1_MINI_ALU_OperationResult_2,
                   L1_0_L2_2_G1_MINI_ALU_OperationResult_1,
                   L1_0_L2_2_G1_MINI_ALU_OperationResult_0}), .BoothOperand ({
                   L1_0_L2_2_G1_MINI_ALU_BoothOperand_16,
                   L1_0_L2_2_G1_MINI_ALU_BoothOperand_15,
                   L1_0_L2_2_G1_MINI_ALU_BoothOperand_14,
                   L1_0_L2_2_G1_MINI_ALU_BoothOperand_13,
                   L1_0_L2_2_G1_MINI_ALU_BoothOperand_12,
                   L1_0_L2_2_G1_MINI_ALU_BoothOperand_11,
                   L1_0_L2_2_G1_MINI_ALU_BoothOperand_10,
                   L1_0_L2_2_G1_MINI_ALU_BoothOperand_9,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16}), .BoothP ({
                   L1_0_L2_2_G1_MINI_ALU_BoothP_16,
                   L1_0_L2_2_G1_MINI_ALU_BoothP_15,
                   L1_0_L2_2_G1_MINI_ALU_BoothP_14,
                   L1_0_L2_2_G1_MINI_ALU_BoothP_13,
                   L1_0_L2_2_G1_MINI_ALU_BoothP_12,
                   L1_0_L2_2_G1_MINI_ALU_BoothP_11,
                   L1_0_L2_2_G1_MINI_ALU_BoothP_10,
                   L1_0_L2_2_G1_MINI_ALU_BoothP_9,L1_0_L2_2_G1_MINI_ALU_BoothP_8
                   ,L1_0_L2_2_G1_MINI_ALU_BoothP_7,
                   L1_0_L2_2_G1_MINI_ALU_BoothP_6,L1_0_L2_2_G1_MINI_ALU_BoothP_5
                   ,L1_0_L2_2_G1_MINI_ALU_BoothP_4,
                   L1_0_L2_2_G1_MINI_ALU_BoothP_3,L1_0_L2_2_G1_MINI_ALU_BoothP_2
                   ,L1_0_L2_2_G1_MINI_ALU_BoothP_1,
                   L1_0_L2_2_G1_MINI_ALU_BoothP_0}), .SelOperand (nx3280), .Operation (
                   L1_0_L2_2_G1_MINI_ALU_BoothXORCheck), .AdderResult ({
                   L1ResultsLarge_2__16,L1ResultsLarge_2__15,
                   L1ResultsLarge_2__14,L1ResultsLarge_2__13,
                   L1ResultsLarge_2__12,L1ResultsLarge_2__11,
                   L1ResultsLarge_2__10,L1ResultsLarge_2__9,L1ResultsLarge_2__8,
                   L1ResultsLarge_2__7,L1ResultsLarge_2__6,L1ResultsLarge_2__5,
                   L1ResultsLarge_2__4,L1ResultsLarge_2__3,L1ResultsLarge_2__2,
                   L1ResultsLarge_2__1,L1ResultsLarge_2__0}), .AdderBoothResult (
                   {\$dummy [70],L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_15,
                   L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_14,
                   L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_13,
                   L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_12,
                   L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_11,
                   L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_10,
                   L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_9,
                   L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_8,
                   L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_7,
                   L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_6,
                   L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_5,
                   L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_4,
                   L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_3,
                   L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_2,
                   L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_1,
                   L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_0})) ;
    booth_unit_17 L1_0_L2_2_G1_MINI_ALU_BOOTH_UNIT (.CLK (CLK), .RST (RST), .Start (
                  Start), .Instr (Instr), .LoopingAndResultNotReady (nx3272), .Filter (
                  {FilterDin_0__2__7,FilterDin_0__2__6,FilterDin_0__2__5,
                  FilterDin_0__2__4,FilterDin_0__2__3,FilterDin_0__2__2,
                  FilterDin_0__2__1,FilterDin_0__2__0}), .Window ({
                  WindowDin_0__2__7,WindowDin_0__2__6,WindowDin_0__2__5,
                  WindowDin_0__2__4,WindowDin_0__2__3,WindowDin_0__2__2,
                  WindowDin_0__2__1,WindowDin_0__2__0}), .AdderBoothResult ({
                  L1FirstOperands_12__16,
                  L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_15,
                  L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_14,
                  L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_13,
                  L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_12,
                  L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_11,
                  L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_10,
                  L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_9,
                  L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_8,
                  L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_7,
                  L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_6,
                  L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_5,
                  L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_4,
                  L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_3,
                  L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_2,
                  L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_1,
                  L1_0_L2_2_G1_MINI_ALU_AdderBoothResult_0}), .BoothXORCheck (
                  L1_0_L2_2_G1_MINI_ALU_BoothXORCheck), .BoothResult ({
                  \$dummy [71],\$dummy [72],\$dummy [73],\$dummy [74],
                  \$dummy [75],\$dummy [76],\$dummy [77],\$dummy [78]}), .BoothAddingOperand (
                  {L1_0_L2_2_G1_MINI_ALU_BoothOperand_16,
                  L1_0_L2_2_G1_MINI_ALU_BoothOperand_15,
                  L1_0_L2_2_G1_MINI_ALU_BoothOperand_14,
                  L1_0_L2_2_G1_MINI_ALU_BoothOperand_13,
                  L1_0_L2_2_G1_MINI_ALU_BoothOperand_12,
                  L1_0_L2_2_G1_MINI_ALU_BoothOperand_11,
                  L1_0_L2_2_G1_MINI_ALU_BoothOperand_10,
                  L1_0_L2_2_G1_MINI_ALU_BoothOperand_9,\$dummy [79],\$dummy [80]
                  ,\$dummy [81],\$dummy [82],\$dummy [83],\$dummy [84],
                  \$dummy [85],\$dummy [86],\$dummy [87]}), .BoothP ({
                  L1_0_L2_2_G1_MINI_ALU_BoothP_16,
                  L1_0_L2_2_G1_MINI_ALU_BoothP_15,
                  L1_0_L2_2_G1_MINI_ALU_BoothP_14,
                  L1_0_L2_2_G1_MINI_ALU_BoothP_13,
                  L1_0_L2_2_G1_MINI_ALU_BoothP_12,
                  L1_0_L2_2_G1_MINI_ALU_BoothP_11,
                  L1_0_L2_2_G1_MINI_ALU_BoothP_10,L1_0_L2_2_G1_MINI_ALU_BoothP_9
                  ,L1_0_L2_2_G1_MINI_ALU_BoothP_8,L1_0_L2_2_G1_MINI_ALU_BoothP_7
                  ,L1_0_L2_2_G1_MINI_ALU_BoothP_6,L1_0_L2_2_G1_MINI_ALU_BoothP_5
                  ,L1_0_L2_2_G1_MINI_ALU_BoothP_4,L1_0_L2_2_G1_MINI_ALU_BoothP_3
                  ,L1_0_L2_2_G1_MINI_ALU_BoothP_2,L1_0_L2_2_G1_MINI_ALU_BoothP_1
                  ,L1_0_L2_2_G1_MINI_ALU_BoothP_0}), .LargeWindowShifted ({
                  \$dummy [88],\$dummy [89],\$dummy [90],\$dummy [91],
                  \$dummy [92],\$dummy [93],\$dummy [94],\$dummy [95],
                  \$dummy [96],\$dummy [97],\$dummy [98],\$dummy [99],
                  \$dummy [100],\$dummy [101],\$dummy [102],\$dummy [103],
                  \$dummy [104]})) ;
    booth_adder_17 L1_0_L2_3_G1_MINI_ALU_BOOTH_ADDER (.AdderFirstOperand ({
                   L1FirstOperands_12__16,L1FirstOperands_3__15,
                   L1FirstOperands_3__14,L1FirstOperands_3__13,
                   L1FirstOperands_3__12,L1FirstOperands_3__11,
                   L1FirstOperands_3__10,L1FirstOperands_3__9,
                   L1FirstOperands_3__8,L1FirstOperands_3__7,
                   L1FirstOperands_3__6,L1FirstOperands_3__5,
                   L1FirstOperands_3__4,L1FirstOperands_3__3,
                   L1FirstOperands_3__2,L1FirstOperands_3__1,
                   L1FirstOperands_3__0}), .AdderSecondOperand ({
                   L1FirstOperands_12__16,
                   L1_0_L2_3_G1_MINI_ALU_OperationResult_15,
                   L1_0_L2_3_G1_MINI_ALU_OperationResult_14,
                   L1_0_L2_3_G1_MINI_ALU_OperationResult_13,
                   L1_0_L2_3_G1_MINI_ALU_OperationResult_12,
                   L1_0_L2_3_G1_MINI_ALU_OperationResult_11,
                   L1_0_L2_3_G1_MINI_ALU_OperationResult_10,
                   L1_0_L2_3_G1_MINI_ALU_OperationResult_9,
                   L1_0_L2_3_G1_MINI_ALU_OperationResult_8,
                   L1_0_L2_3_G1_MINI_ALU_OperationResult_7,
                   L1_0_L2_3_G1_MINI_ALU_OperationResult_6,
                   L1_0_L2_3_G1_MINI_ALU_OperationResult_5,
                   L1_0_L2_3_G1_MINI_ALU_OperationResult_4,
                   L1_0_L2_3_G1_MINI_ALU_OperationResult_3,
                   L1_0_L2_3_G1_MINI_ALU_OperationResult_2,
                   L1_0_L2_3_G1_MINI_ALU_OperationResult_1,
                   L1_0_L2_3_G1_MINI_ALU_OperationResult_0}), .BoothOperand ({
                   L1_0_L2_3_G1_MINI_ALU_BoothOperand_16,
                   L1_0_L2_3_G1_MINI_ALU_BoothOperand_15,
                   L1_0_L2_3_G1_MINI_ALU_BoothOperand_14,
                   L1_0_L2_3_G1_MINI_ALU_BoothOperand_13,
                   L1_0_L2_3_G1_MINI_ALU_BoothOperand_12,
                   L1_0_L2_3_G1_MINI_ALU_BoothOperand_11,
                   L1_0_L2_3_G1_MINI_ALU_BoothOperand_10,
                   L1_0_L2_3_G1_MINI_ALU_BoothOperand_9,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16}), .BoothP ({
                   L1_0_L2_3_G1_MINI_ALU_BoothP_16,
                   L1_0_L2_3_G1_MINI_ALU_BoothP_15,
                   L1_0_L2_3_G1_MINI_ALU_BoothP_14,
                   L1_0_L2_3_G1_MINI_ALU_BoothP_13,
                   L1_0_L2_3_G1_MINI_ALU_BoothP_12,
                   L1_0_L2_3_G1_MINI_ALU_BoothP_11,
                   L1_0_L2_3_G1_MINI_ALU_BoothP_10,
                   L1_0_L2_3_G1_MINI_ALU_BoothP_9,L1_0_L2_3_G1_MINI_ALU_BoothP_8
                   ,L1_0_L2_3_G1_MINI_ALU_BoothP_7,
                   L1_0_L2_3_G1_MINI_ALU_BoothP_6,L1_0_L2_3_G1_MINI_ALU_BoothP_5
                   ,L1_0_L2_3_G1_MINI_ALU_BoothP_4,
                   L1_0_L2_3_G1_MINI_ALU_BoothP_3,L1_0_L2_3_G1_MINI_ALU_BoothP_2
                   ,L1_0_L2_3_G1_MINI_ALU_BoothP_1,
                   L1_0_L2_3_G1_MINI_ALU_BoothP_0}), .SelOperand (nx3280), .Operation (
                   L1_0_L2_3_G1_MINI_ALU_BoothXORCheck), .AdderResult ({
                   L1ResultsLarge_3__16,L1ResultsLarge_3__15,
                   L1ResultsLarge_3__14,L1ResultsLarge_3__13,
                   L1ResultsLarge_3__12,L1ResultsLarge_3__11,
                   L1ResultsLarge_3__10,L1ResultsLarge_3__9,L1ResultsLarge_3__8,
                   L1ResultsLarge_3__7,L1ResultsLarge_3__6,L1ResultsLarge_3__5,
                   L1ResultsLarge_3__4,L1ResultsLarge_3__3,L1ResultsLarge_3__2,
                   L1ResultsLarge_3__1,L1ResultsLarge_3__0}), .AdderBoothResult (
                   {\$dummy [105],L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_15,
                   L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_14,
                   L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_13,
                   L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_12,
                   L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_11,
                   L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_10,
                   L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_9,
                   L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_8,
                   L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_7,
                   L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_6,
                   L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_5,
                   L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_4,
                   L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_3,
                   L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_2,
                   L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_1,
                   L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_0})) ;
    booth_unit_17 L1_0_L2_3_G1_MINI_ALU_BOOTH_UNIT (.CLK (CLK), .RST (RST), .Start (
                  Start), .Instr (Instr), .LoopingAndResultNotReady (nx3272), .Filter (
                  {FilterDin_0__3__7,FilterDin_0__3__6,FilterDin_0__3__5,
                  FilterDin_0__3__4,FilterDin_0__3__3,FilterDin_0__3__2,
                  FilterDin_0__3__1,FilterDin_0__3__0}), .Window ({
                  WindowDin_0__3__7,WindowDin_0__3__6,WindowDin_0__3__5,
                  WindowDin_0__3__4,WindowDin_0__3__3,WindowDin_0__3__2,
                  WindowDin_0__3__1,WindowDin_0__3__0}), .AdderBoothResult ({
                  L1FirstOperands_12__16,
                  L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_15,
                  L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_14,
                  L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_13,
                  L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_12,
                  L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_11,
                  L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_10,
                  L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_9,
                  L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_8,
                  L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_7,
                  L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_6,
                  L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_5,
                  L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_4,
                  L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_3,
                  L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_2,
                  L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_1,
                  L1_0_L2_3_G1_MINI_ALU_AdderBoothResult_0}), .BoothXORCheck (
                  L1_0_L2_3_G1_MINI_ALU_BoothXORCheck), .BoothResult ({
                  \$dummy [106],\$dummy [107],\$dummy [108],\$dummy [109],
                  \$dummy [110],\$dummy [111],\$dummy [112],\$dummy [113]}), .BoothAddingOperand (
                  {L1_0_L2_3_G1_MINI_ALU_BoothOperand_16,
                  L1_0_L2_3_G1_MINI_ALU_BoothOperand_15,
                  L1_0_L2_3_G1_MINI_ALU_BoothOperand_14,
                  L1_0_L2_3_G1_MINI_ALU_BoothOperand_13,
                  L1_0_L2_3_G1_MINI_ALU_BoothOperand_12,
                  L1_0_L2_3_G1_MINI_ALU_BoothOperand_11,
                  L1_0_L2_3_G1_MINI_ALU_BoothOperand_10,
                  L1_0_L2_3_G1_MINI_ALU_BoothOperand_9,\$dummy [114],
                  \$dummy [115],\$dummy [116],\$dummy [117],\$dummy [118],
                  \$dummy [119],\$dummy [120],\$dummy [121],\$dummy [122]}), .BoothP (
                  {L1_0_L2_3_G1_MINI_ALU_BoothP_16,
                  L1_0_L2_3_G1_MINI_ALU_BoothP_15,
                  L1_0_L2_3_G1_MINI_ALU_BoothP_14,
                  L1_0_L2_3_G1_MINI_ALU_BoothP_13,
                  L1_0_L2_3_G1_MINI_ALU_BoothP_12,
                  L1_0_L2_3_G1_MINI_ALU_BoothP_11,
                  L1_0_L2_3_G1_MINI_ALU_BoothP_10,L1_0_L2_3_G1_MINI_ALU_BoothP_9
                  ,L1_0_L2_3_G1_MINI_ALU_BoothP_8,L1_0_L2_3_G1_MINI_ALU_BoothP_7
                  ,L1_0_L2_3_G1_MINI_ALU_BoothP_6,L1_0_L2_3_G1_MINI_ALU_BoothP_5
                  ,L1_0_L2_3_G1_MINI_ALU_BoothP_4,L1_0_L2_3_G1_MINI_ALU_BoothP_3
                  ,L1_0_L2_3_G1_MINI_ALU_BoothP_2,L1_0_L2_3_G1_MINI_ALU_BoothP_1
                  ,L1_0_L2_3_G1_MINI_ALU_BoothP_0}), .LargeWindowShifted ({
                  \$dummy [123],\$dummy [124],\$dummy [125],\$dummy [126],
                  \$dummy [127],\$dummy [128],\$dummy [129],\$dummy [130],
                  \$dummy [131],\$dummy [132],\$dummy [133],\$dummy [134],
                  \$dummy [135],\$dummy [136],\$dummy [137],\$dummy [138],
                  \$dummy [139]})) ;
    booth_adder_17 L1_0_L2_4_G1_MINI_ALU_BOOTH_ADDER (.AdderFirstOperand ({
                   L1FirstOperands_12__16,L1FirstOperands_4__15,
                   L1FirstOperands_4__14,L1FirstOperands_4__13,
                   L1FirstOperands_4__12,L1FirstOperands_4__11,
                   L1FirstOperands_4__10,L1FirstOperands_4__9,
                   L1FirstOperands_4__8,L1FirstOperands_4__7,
                   L1FirstOperands_4__6,L1FirstOperands_4__5,
                   L1FirstOperands_4__4,L1FirstOperands_4__3,
                   L1FirstOperands_4__2,L1FirstOperands_4__1,
                   L1FirstOperands_4__0}), .AdderSecondOperand ({
                   L1FirstOperands_12__16,
                   L1_0_L2_4_G1_MINI_ALU_OperationResult_15,
                   L1_0_L2_4_G1_MINI_ALU_OperationResult_14,
                   L1_0_L2_4_G1_MINI_ALU_OperationResult_13,
                   L1_0_L2_4_G1_MINI_ALU_OperationResult_12,
                   L1_0_L2_4_G1_MINI_ALU_OperationResult_11,
                   L1_0_L2_4_G1_MINI_ALU_OperationResult_10,
                   L1_0_L2_4_G1_MINI_ALU_OperationResult_9,
                   L1_0_L2_4_G1_MINI_ALU_OperationResult_8,
                   L1_0_L2_4_G1_MINI_ALU_OperationResult_7,
                   L1_0_L2_4_G1_MINI_ALU_OperationResult_6,
                   L1_0_L2_4_G1_MINI_ALU_OperationResult_5,
                   L1_0_L2_4_G1_MINI_ALU_OperationResult_4,
                   L1_0_L2_4_G1_MINI_ALU_OperationResult_3,
                   L1_0_L2_4_G1_MINI_ALU_OperationResult_2,
                   L1_0_L2_4_G1_MINI_ALU_OperationResult_1,
                   L1_0_L2_4_G1_MINI_ALU_OperationResult_0}), .BoothOperand ({
                   L1_0_L2_4_G1_MINI_ALU_BoothOperand_16,
                   L1_0_L2_4_G1_MINI_ALU_BoothOperand_15,
                   L1_0_L2_4_G1_MINI_ALU_BoothOperand_14,
                   L1_0_L2_4_G1_MINI_ALU_BoothOperand_13,
                   L1_0_L2_4_G1_MINI_ALU_BoothOperand_12,
                   L1_0_L2_4_G1_MINI_ALU_BoothOperand_11,
                   L1_0_L2_4_G1_MINI_ALU_BoothOperand_10,
                   L1_0_L2_4_G1_MINI_ALU_BoothOperand_9,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16}), .BoothP ({
                   L1_0_L2_4_G1_MINI_ALU_BoothP_16,
                   L1_0_L2_4_G1_MINI_ALU_BoothP_15,
                   L1_0_L2_4_G1_MINI_ALU_BoothP_14,
                   L1_0_L2_4_G1_MINI_ALU_BoothP_13,
                   L1_0_L2_4_G1_MINI_ALU_BoothP_12,
                   L1_0_L2_4_G1_MINI_ALU_BoothP_11,
                   L1_0_L2_4_G1_MINI_ALU_BoothP_10,
                   L1_0_L2_4_G1_MINI_ALU_BoothP_9,L1_0_L2_4_G1_MINI_ALU_BoothP_8
                   ,L1_0_L2_4_G1_MINI_ALU_BoothP_7,
                   L1_0_L2_4_G1_MINI_ALU_BoothP_6,L1_0_L2_4_G1_MINI_ALU_BoothP_5
                   ,L1_0_L2_4_G1_MINI_ALU_BoothP_4,
                   L1_0_L2_4_G1_MINI_ALU_BoothP_3,L1_0_L2_4_G1_MINI_ALU_BoothP_2
                   ,L1_0_L2_4_G1_MINI_ALU_BoothP_1,
                   L1_0_L2_4_G1_MINI_ALU_BoothP_0}), .SelOperand (nx3280), .Operation (
                   L1_0_L2_4_G1_MINI_ALU_BoothXORCheck), .AdderResult ({
                   L1ResultsLarge_4__16,L1ResultsLarge_4__15,
                   L1ResultsLarge_4__14,L1ResultsLarge_4__13,
                   L1ResultsLarge_4__12,L1ResultsLarge_4__11,
                   L1ResultsLarge_4__10,L1ResultsLarge_4__9,L1ResultsLarge_4__8,
                   L1ResultsLarge_4__7,L1ResultsLarge_4__6,L1ResultsLarge_4__5,
                   L1ResultsLarge_4__4,L1ResultsLarge_4__3,L1ResultsLarge_4__2,
                   L1ResultsLarge_4__1,L1ResultsLarge_4__0}), .AdderBoothResult (
                   {\$dummy [140],L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_15,
                   L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_14,
                   L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_13,
                   L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_12,
                   L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_11,
                   L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_10,
                   L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_9,
                   L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_8,
                   L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_7,
                   L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_6,
                   L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_5,
                   L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_4,
                   L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_3,
                   L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_2,
                   L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_1,
                   L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_0})) ;
    booth_unit_17 L1_0_L2_4_G1_MINI_ALU_BOOTH_UNIT (.CLK (CLK), .RST (RST), .Start (
                  Start), .Instr (Instr), .LoopingAndResultNotReady (nx3272), .Filter (
                  {FilterDin_0__4__7,FilterDin_0__4__6,FilterDin_0__4__5,
                  FilterDin_0__4__4,FilterDin_0__4__3,FilterDin_0__4__2,
                  FilterDin_0__4__1,FilterDin_0__4__0}), .Window ({
                  WindowDin_0__4__7,WindowDin_0__4__6,WindowDin_0__4__5,
                  WindowDin_0__4__4,WindowDin_0__4__3,WindowDin_0__4__2,
                  WindowDin_0__4__1,WindowDin_0__4__0}), .AdderBoothResult ({
                  L1FirstOperands_12__16,
                  L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_15,
                  L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_14,
                  L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_13,
                  L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_12,
                  L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_11,
                  L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_10,
                  L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_9,
                  L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_8,
                  L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_7,
                  L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_6,
                  L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_5,
                  L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_4,
                  L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_3,
                  L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_2,
                  L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_1,
                  L1_0_L2_4_G1_MINI_ALU_AdderBoothResult_0}), .BoothXORCheck (
                  L1_0_L2_4_G1_MINI_ALU_BoothXORCheck), .BoothResult ({
                  \$dummy [141],\$dummy [142],\$dummy [143],\$dummy [144],
                  \$dummy [145],\$dummy [146],\$dummy [147],\$dummy [148]}), .BoothAddingOperand (
                  {L1_0_L2_4_G1_MINI_ALU_BoothOperand_16,
                  L1_0_L2_4_G1_MINI_ALU_BoothOperand_15,
                  L1_0_L2_4_G1_MINI_ALU_BoothOperand_14,
                  L1_0_L2_4_G1_MINI_ALU_BoothOperand_13,
                  L1_0_L2_4_G1_MINI_ALU_BoothOperand_12,
                  L1_0_L2_4_G1_MINI_ALU_BoothOperand_11,
                  L1_0_L2_4_G1_MINI_ALU_BoothOperand_10,
                  L1_0_L2_4_G1_MINI_ALU_BoothOperand_9,\$dummy [149],
                  \$dummy [150],\$dummy [151],\$dummy [152],\$dummy [153],
                  \$dummy [154],\$dummy [155],\$dummy [156],\$dummy [157]}), .BoothP (
                  {L1_0_L2_4_G1_MINI_ALU_BoothP_16,
                  L1_0_L2_4_G1_MINI_ALU_BoothP_15,
                  L1_0_L2_4_G1_MINI_ALU_BoothP_14,
                  L1_0_L2_4_G1_MINI_ALU_BoothP_13,
                  L1_0_L2_4_G1_MINI_ALU_BoothP_12,
                  L1_0_L2_4_G1_MINI_ALU_BoothP_11,
                  L1_0_L2_4_G1_MINI_ALU_BoothP_10,L1_0_L2_4_G1_MINI_ALU_BoothP_9
                  ,L1_0_L2_4_G1_MINI_ALU_BoothP_8,L1_0_L2_4_G1_MINI_ALU_BoothP_7
                  ,L1_0_L2_4_G1_MINI_ALU_BoothP_6,L1_0_L2_4_G1_MINI_ALU_BoothP_5
                  ,L1_0_L2_4_G1_MINI_ALU_BoothP_4,L1_0_L2_4_G1_MINI_ALU_BoothP_3
                  ,L1_0_L2_4_G1_MINI_ALU_BoothP_2,L1_0_L2_4_G1_MINI_ALU_BoothP_1
                  ,L1_0_L2_4_G1_MINI_ALU_BoothP_0}), .LargeWindowShifted ({
                  \$dummy [158],\$dummy [159],\$dummy [160],\$dummy [161],
                  \$dummy [162],\$dummy [163],\$dummy [164],\$dummy [165],
                  \$dummy [166],\$dummy [167],\$dummy [168],\$dummy [169],
                  \$dummy [170],\$dummy [171],\$dummy [172],\$dummy [173],
                  \$dummy [174]})) ;
    booth_adder_17 L1_1_L2_0_G1_MINI_ALU_BOOTH_ADDER (.AdderFirstOperand ({
                   L1FirstOperands_12__16,L1FirstOperands_2__15,
                   L1FirstOperands_2__14,L1FirstOperands_2__13,
                   L1FirstOperands_2__12,L1FirstOperands_2__11,
                   L1FirstOperands_2__10,L1FirstOperands_2__9,
                   L1FirstOperands_2__8,L1FirstOperands_2__7,
                   L1FirstOperands_2__6,L1FirstOperands_2__5,
                   L1FirstOperands_2__4,L1FirstOperands_2__3,
                   L1FirstOperands_2__2,L1FirstOperands_2__1,
                   L1FirstOperands_2__0}), .AdderSecondOperand ({
                   L1FirstOperands_12__16,
                   L1_1_L2_0_G1_MINI_ALU_OperationResult_15,
                   L1_1_L2_0_G1_MINI_ALU_OperationResult_14,
                   L1_1_L2_0_G1_MINI_ALU_OperationResult_13,
                   L1_1_L2_0_G1_MINI_ALU_OperationResult_12,
                   L1_1_L2_0_G1_MINI_ALU_OperationResult_11,
                   L1_1_L2_0_G1_MINI_ALU_OperationResult_10,
                   L1_1_L2_0_G1_MINI_ALU_OperationResult_9,
                   L1_1_L2_0_G1_MINI_ALU_OperationResult_8,
                   L1_1_L2_0_G1_MINI_ALU_OperationResult_7,
                   L1_1_L2_0_G1_MINI_ALU_OperationResult_6,
                   L1_1_L2_0_G1_MINI_ALU_OperationResult_5,
                   L1_1_L2_0_G1_MINI_ALU_OperationResult_4,
                   L1_1_L2_0_G1_MINI_ALU_OperationResult_3,
                   L1_1_L2_0_G1_MINI_ALU_OperationResult_2,
                   L1_1_L2_0_G1_MINI_ALU_OperationResult_1,
                   L1_1_L2_0_G1_MINI_ALU_OperationResult_0}), .BoothOperand ({
                   L1_1_L2_0_G1_MINI_ALU_BoothOperand_16,
                   L1_1_L2_0_G1_MINI_ALU_BoothOperand_15,
                   L1_1_L2_0_G1_MINI_ALU_BoothOperand_14,
                   L1_1_L2_0_G1_MINI_ALU_BoothOperand_13,
                   L1_1_L2_0_G1_MINI_ALU_BoothOperand_12,
                   L1_1_L2_0_G1_MINI_ALU_BoothOperand_11,
                   L1_1_L2_0_G1_MINI_ALU_BoothOperand_10,
                   L1_1_L2_0_G1_MINI_ALU_BoothOperand_9,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16}), .BoothP ({
                   L1_1_L2_0_G1_MINI_ALU_BoothP_16,
                   L1_1_L2_0_G1_MINI_ALU_BoothP_15,
                   L1_1_L2_0_G1_MINI_ALU_BoothP_14,
                   L1_1_L2_0_G1_MINI_ALU_BoothP_13,
                   L1_1_L2_0_G1_MINI_ALU_BoothP_12,
                   L1_1_L2_0_G1_MINI_ALU_BoothP_11,
                   L1_1_L2_0_G1_MINI_ALU_BoothP_10,
                   L1_1_L2_0_G1_MINI_ALU_BoothP_9,L1_1_L2_0_G1_MINI_ALU_BoothP_8
                   ,L1_1_L2_0_G1_MINI_ALU_BoothP_7,
                   L1_1_L2_0_G1_MINI_ALU_BoothP_6,L1_1_L2_0_G1_MINI_ALU_BoothP_5
                   ,L1_1_L2_0_G1_MINI_ALU_BoothP_4,
                   L1_1_L2_0_G1_MINI_ALU_BoothP_3,L1_1_L2_0_G1_MINI_ALU_BoothP_2
                   ,L1_1_L2_0_G1_MINI_ALU_BoothP_1,
                   L1_1_L2_0_G1_MINI_ALU_BoothP_0}), .SelOperand (nx3280), .Operation (
                   L1_1_L2_0_G1_MINI_ALU_BoothXORCheck), .AdderResult ({
                   L1ResultsLarge_5__16,L1ResultsLarge_5__15,
                   L1ResultsLarge_5__14,L1ResultsLarge_5__13,
                   L1ResultsLarge_5__12,L1ResultsLarge_5__11,
                   L1ResultsLarge_5__10,L1ResultsLarge_5__9,L1ResultsLarge_5__8,
                   L1ResultsLarge_5__7,L1ResultsLarge_5__6,L1ResultsLarge_5__5,
                   L1ResultsLarge_5__4,L1ResultsLarge_5__3,L1ResultsLarge_5__2,
                   L1ResultsLarge_5__1,L1ResultsLarge_5__0}), .AdderBoothResult (
                   {\$dummy [175],L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_15,
                   L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_14,
                   L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_13,
                   L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_12,
                   L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_11,
                   L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_10,
                   L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_9,
                   L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_8,
                   L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_7,
                   L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_6,
                   L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_5,
                   L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_4,
                   L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_3,
                   L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_2,
                   L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_1,
                   L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_0})) ;
    booth_unit_17 L1_1_L2_0_G1_MINI_ALU_BOOTH_UNIT (.CLK (CLK), .RST (RST), .Start (
                  Start), .Instr (Instr), .LoopingAndResultNotReady (nx3272), .Filter (
                  {FilterDin_1__0__7,FilterDin_1__0__6,FilterDin_1__0__5,
                  FilterDin_1__0__4,FilterDin_1__0__3,FilterDin_1__0__2,
                  FilterDin_1__0__1,FilterDin_1__0__0}), .Window ({
                  WindowDin_1__0__7,WindowDin_1__0__6,WindowDin_1__0__5,
                  WindowDin_1__0__4,WindowDin_1__0__3,WindowDin_1__0__2,
                  WindowDin_1__0__1,WindowDin_1__0__0}), .AdderBoothResult ({
                  L1FirstOperands_12__16,
                  L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_15,
                  L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_14,
                  L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_13,
                  L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_12,
                  L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_11,
                  L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_10,
                  L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_9,
                  L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_8,
                  L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_7,
                  L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_6,
                  L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_5,
                  L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_4,
                  L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_3,
                  L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_2,
                  L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_1,
                  L1_1_L2_0_G1_MINI_ALU_AdderBoothResult_0}), .BoothXORCheck (
                  L1_1_L2_0_G1_MINI_ALU_BoothXORCheck), .BoothResult ({
                  \$dummy [176],\$dummy [177],\$dummy [178],\$dummy [179],
                  \$dummy [180],\$dummy [181],\$dummy [182],\$dummy [183]}), .BoothAddingOperand (
                  {L1_1_L2_0_G1_MINI_ALU_BoothOperand_16,
                  L1_1_L2_0_G1_MINI_ALU_BoothOperand_15,
                  L1_1_L2_0_G1_MINI_ALU_BoothOperand_14,
                  L1_1_L2_0_G1_MINI_ALU_BoothOperand_13,
                  L1_1_L2_0_G1_MINI_ALU_BoothOperand_12,
                  L1_1_L2_0_G1_MINI_ALU_BoothOperand_11,
                  L1_1_L2_0_G1_MINI_ALU_BoothOperand_10,
                  L1_1_L2_0_G1_MINI_ALU_BoothOperand_9,\$dummy [184],
                  \$dummy [185],\$dummy [186],\$dummy [187],\$dummy [188],
                  \$dummy [189],\$dummy [190],\$dummy [191],\$dummy [192]}), .BoothP (
                  {L1_1_L2_0_G1_MINI_ALU_BoothP_16,
                  L1_1_L2_0_G1_MINI_ALU_BoothP_15,
                  L1_1_L2_0_G1_MINI_ALU_BoothP_14,
                  L1_1_L2_0_G1_MINI_ALU_BoothP_13,
                  L1_1_L2_0_G1_MINI_ALU_BoothP_12,
                  L1_1_L2_0_G1_MINI_ALU_BoothP_11,
                  L1_1_L2_0_G1_MINI_ALU_BoothP_10,L1_1_L2_0_G1_MINI_ALU_BoothP_9
                  ,L1_1_L2_0_G1_MINI_ALU_BoothP_8,L1_1_L2_0_G1_MINI_ALU_BoothP_7
                  ,L1_1_L2_0_G1_MINI_ALU_BoothP_6,L1_1_L2_0_G1_MINI_ALU_BoothP_5
                  ,L1_1_L2_0_G1_MINI_ALU_BoothP_4,L1_1_L2_0_G1_MINI_ALU_BoothP_3
                  ,L1_1_L2_0_G1_MINI_ALU_BoothP_2,L1_1_L2_0_G1_MINI_ALU_BoothP_1
                  ,L1_1_L2_0_G1_MINI_ALU_BoothP_0}), .LargeWindowShifted ({
                  \$dummy [193],\$dummy [194],\$dummy [195],\$dummy [196],
                  \$dummy [197],\$dummy [198],\$dummy [199],\$dummy [200],
                  \$dummy [201],\$dummy [202],\$dummy [203],\$dummy [204],
                  \$dummy [205],\$dummy [206],\$dummy [207],\$dummy [208],
                  \$dummy [209]})) ;
    booth_adder_17 L1_1_L2_1_G1_MINI_ALU_BOOTH_ADDER (.AdderFirstOperand ({
                   L1FirstOperands_12__16,L1FirstOperands_6__15,
                   L1FirstOperands_6__14,L1FirstOperands_6__13,
                   L1FirstOperands_6__12,L1FirstOperands_6__11,
                   L1FirstOperands_6__10,L1FirstOperands_6__9,
                   L1FirstOperands_6__8,L1FirstOperands_6__7,
                   L1FirstOperands_6__6,L1FirstOperands_6__5,
                   L1FirstOperands_6__4,L1FirstOperands_6__3,
                   L1FirstOperands_6__2,L1FirstOperands_6__1,
                   L1FirstOperands_6__0}), .AdderSecondOperand ({
                   L1FirstOperands_12__16,
                   L1_1_L2_1_G1_MINI_ALU_OperationResult_15,
                   L1_1_L2_1_G1_MINI_ALU_OperationResult_14,
                   L1_1_L2_1_G1_MINI_ALU_OperationResult_13,
                   L1_1_L2_1_G1_MINI_ALU_OperationResult_12,
                   L1_1_L2_1_G1_MINI_ALU_OperationResult_11,
                   L1_1_L2_1_G1_MINI_ALU_OperationResult_10,
                   L1_1_L2_1_G1_MINI_ALU_OperationResult_9,
                   L1_1_L2_1_G1_MINI_ALU_OperationResult_8,
                   L1_1_L2_1_G1_MINI_ALU_OperationResult_7,
                   L1_1_L2_1_G1_MINI_ALU_OperationResult_6,
                   L1_1_L2_1_G1_MINI_ALU_OperationResult_5,
                   L1_1_L2_1_G1_MINI_ALU_OperationResult_4,
                   L1_1_L2_1_G1_MINI_ALU_OperationResult_3,
                   L1_1_L2_1_G1_MINI_ALU_OperationResult_2,
                   L1_1_L2_1_G1_MINI_ALU_OperationResult_1,
                   L1_1_L2_1_G1_MINI_ALU_OperationResult_0}), .BoothOperand ({
                   L1_1_L2_1_G1_MINI_ALU_BoothOperand_16,
                   L1_1_L2_1_G1_MINI_ALU_BoothOperand_15,
                   L1_1_L2_1_G1_MINI_ALU_BoothOperand_14,
                   L1_1_L2_1_G1_MINI_ALU_BoothOperand_13,
                   L1_1_L2_1_G1_MINI_ALU_BoothOperand_12,
                   L1_1_L2_1_G1_MINI_ALU_BoothOperand_11,
                   L1_1_L2_1_G1_MINI_ALU_BoothOperand_10,
                   L1_1_L2_1_G1_MINI_ALU_BoothOperand_9,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16}), .BoothP ({
                   L1_1_L2_1_G1_MINI_ALU_BoothP_16,
                   L1_1_L2_1_G1_MINI_ALU_BoothP_15,
                   L1_1_L2_1_G1_MINI_ALU_BoothP_14,
                   L1_1_L2_1_G1_MINI_ALU_BoothP_13,
                   L1_1_L2_1_G1_MINI_ALU_BoothP_12,
                   L1_1_L2_1_G1_MINI_ALU_BoothP_11,
                   L1_1_L2_1_G1_MINI_ALU_BoothP_10,
                   L1_1_L2_1_G1_MINI_ALU_BoothP_9,L1_1_L2_1_G1_MINI_ALU_BoothP_8
                   ,L1_1_L2_1_G1_MINI_ALU_BoothP_7,
                   L1_1_L2_1_G1_MINI_ALU_BoothP_6,L1_1_L2_1_G1_MINI_ALU_BoothP_5
                   ,L1_1_L2_1_G1_MINI_ALU_BoothP_4,
                   L1_1_L2_1_G1_MINI_ALU_BoothP_3,L1_1_L2_1_G1_MINI_ALU_BoothP_2
                   ,L1_1_L2_1_G1_MINI_ALU_BoothP_1,
                   L1_1_L2_1_G1_MINI_ALU_BoothP_0}), .SelOperand (nx3280), .Operation (
                   L1_1_L2_1_G1_MINI_ALU_BoothXORCheck), .AdderResult ({
                   L1ResultsLarge_6__16,L1ResultsLarge_6__15,
                   L1ResultsLarge_6__14,L1ResultsLarge_6__13,
                   L1ResultsLarge_6__12,L1ResultsLarge_6__11,
                   L1ResultsLarge_6__10,L1ResultsLarge_6__9,L1ResultsLarge_6__8,
                   L1ResultsLarge_6__7,L1ResultsLarge_6__6,L1ResultsLarge_6__5,
                   L1ResultsLarge_6__4,L1ResultsLarge_6__3,L1ResultsLarge_6__2,
                   L1ResultsLarge_6__1,L1ResultsLarge_6__0}), .AdderBoothResult (
                   {\$dummy [210],L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_15,
                   L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_14,
                   L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_13,
                   L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_12,
                   L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_11,
                   L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_10,
                   L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_9,
                   L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_8,
                   L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_7,
                   L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_6,
                   L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_5,
                   L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_4,
                   L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_3,
                   L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_2,
                   L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_1,
                   L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_0})) ;
    booth_unit_17 L1_1_L2_1_G1_MINI_ALU_BOOTH_UNIT (.CLK (CLK), .RST (RST), .Start (
                  Start), .Instr (Instr), .LoopingAndResultNotReady (nx3272), .Filter (
                  {FilterDin_1__1__7,FilterDin_1__1__6,FilterDin_1__1__5,
                  FilterDin_1__1__4,FilterDin_1__1__3,FilterDin_1__1__2,
                  FilterDin_1__1__1,FilterDin_1__1__0}), .Window ({
                  WindowDin_1__1__7,WindowDin_1__1__6,WindowDin_1__1__5,
                  WindowDin_1__1__4,WindowDin_1__1__3,WindowDin_1__1__2,
                  WindowDin_1__1__1,WindowDin_1__1__0}), .AdderBoothResult ({
                  L1FirstOperands_12__16,
                  L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_15,
                  L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_14,
                  L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_13,
                  L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_12,
                  L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_11,
                  L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_10,
                  L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_9,
                  L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_8,
                  L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_7,
                  L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_6,
                  L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_5,
                  L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_4,
                  L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_3,
                  L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_2,
                  L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_1,
                  L1_1_L2_1_G1_MINI_ALU_AdderBoothResult_0}), .BoothXORCheck (
                  L1_1_L2_1_G1_MINI_ALU_BoothXORCheck), .BoothResult ({
                  \$dummy [211],\$dummy [212],\$dummy [213],\$dummy [214],
                  \$dummy [215],\$dummy [216],\$dummy [217],\$dummy [218]}), .BoothAddingOperand (
                  {L1_1_L2_1_G1_MINI_ALU_BoothOperand_16,
                  L1_1_L2_1_G1_MINI_ALU_BoothOperand_15,
                  L1_1_L2_1_G1_MINI_ALU_BoothOperand_14,
                  L1_1_L2_1_G1_MINI_ALU_BoothOperand_13,
                  L1_1_L2_1_G1_MINI_ALU_BoothOperand_12,
                  L1_1_L2_1_G1_MINI_ALU_BoothOperand_11,
                  L1_1_L2_1_G1_MINI_ALU_BoothOperand_10,
                  L1_1_L2_1_G1_MINI_ALU_BoothOperand_9,\$dummy [219],
                  \$dummy [220],\$dummy [221],\$dummy [222],\$dummy [223],
                  \$dummy [224],\$dummy [225],\$dummy [226],\$dummy [227]}), .BoothP (
                  {L1_1_L2_1_G1_MINI_ALU_BoothP_16,
                  L1_1_L2_1_G1_MINI_ALU_BoothP_15,
                  L1_1_L2_1_G1_MINI_ALU_BoothP_14,
                  L1_1_L2_1_G1_MINI_ALU_BoothP_13,
                  L1_1_L2_1_G1_MINI_ALU_BoothP_12,
                  L1_1_L2_1_G1_MINI_ALU_BoothP_11,
                  L1_1_L2_1_G1_MINI_ALU_BoothP_10,L1_1_L2_1_G1_MINI_ALU_BoothP_9
                  ,L1_1_L2_1_G1_MINI_ALU_BoothP_8,L1_1_L2_1_G1_MINI_ALU_BoothP_7
                  ,L1_1_L2_1_G1_MINI_ALU_BoothP_6,L1_1_L2_1_G1_MINI_ALU_BoothP_5
                  ,L1_1_L2_1_G1_MINI_ALU_BoothP_4,L1_1_L2_1_G1_MINI_ALU_BoothP_3
                  ,L1_1_L2_1_G1_MINI_ALU_BoothP_2,L1_1_L2_1_G1_MINI_ALU_BoothP_1
                  ,L1_1_L2_1_G1_MINI_ALU_BoothP_0}), .LargeWindowShifted ({
                  \$dummy [228],\$dummy [229],\$dummy [230],\$dummy [231],
                  \$dummy [232],\$dummy [233],\$dummy [234],\$dummy [235],
                  \$dummy [236],\$dummy [237],\$dummy [238],\$dummy [239],
                  \$dummy [240],\$dummy [241],\$dummy [242],\$dummy [243],
                  \$dummy [244]})) ;
    booth_adder_17 L1_1_L2_2_G1_MINI_ALU_BOOTH_ADDER (.AdderFirstOperand ({
                   L1FirstOperands_12__16,L1FirstOperands_7__15,
                   L1FirstOperands_7__14,L1FirstOperands_7__13,
                   L1FirstOperands_7__12,L1FirstOperands_7__11,
                   L1FirstOperands_7__10,L1FirstOperands_7__9,
                   L1FirstOperands_7__8,L1FirstOperands_7__7,
                   L1FirstOperands_7__6,L1FirstOperands_7__5,
                   L1FirstOperands_7__4,L1FirstOperands_7__3,
                   L1FirstOperands_7__2,L1FirstOperands_7__1,
                   L1FirstOperands_7__0}), .AdderSecondOperand ({
                   L1FirstOperands_12__16,
                   L1_1_L2_2_G1_MINI_ALU_OperationResult_15,
                   L1_1_L2_2_G1_MINI_ALU_OperationResult_14,
                   L1_1_L2_2_G1_MINI_ALU_OperationResult_13,
                   L1_1_L2_2_G1_MINI_ALU_OperationResult_12,
                   L1_1_L2_2_G1_MINI_ALU_OperationResult_11,
                   L1_1_L2_2_G1_MINI_ALU_OperationResult_10,
                   L1_1_L2_2_G1_MINI_ALU_OperationResult_9,
                   L1_1_L2_2_G1_MINI_ALU_OperationResult_8,
                   L1_1_L2_2_G1_MINI_ALU_OperationResult_7,
                   L1_1_L2_2_G1_MINI_ALU_OperationResult_6,
                   L1_1_L2_2_G1_MINI_ALU_OperationResult_5,
                   L1_1_L2_2_G1_MINI_ALU_OperationResult_4,
                   L1_1_L2_2_G1_MINI_ALU_OperationResult_3,
                   L1_1_L2_2_G1_MINI_ALU_OperationResult_2,
                   L1_1_L2_2_G1_MINI_ALU_OperationResult_1,
                   L1_1_L2_2_G1_MINI_ALU_OperationResult_0}), .BoothOperand ({
                   L1_1_L2_2_G1_MINI_ALU_BoothOperand_16,
                   L1_1_L2_2_G1_MINI_ALU_BoothOperand_15,
                   L1_1_L2_2_G1_MINI_ALU_BoothOperand_14,
                   L1_1_L2_2_G1_MINI_ALU_BoothOperand_13,
                   L1_1_L2_2_G1_MINI_ALU_BoothOperand_12,
                   L1_1_L2_2_G1_MINI_ALU_BoothOperand_11,
                   L1_1_L2_2_G1_MINI_ALU_BoothOperand_10,
                   L1_1_L2_2_G1_MINI_ALU_BoothOperand_9,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16}), .BoothP ({
                   L1_1_L2_2_G1_MINI_ALU_BoothP_16,
                   L1_1_L2_2_G1_MINI_ALU_BoothP_15,
                   L1_1_L2_2_G1_MINI_ALU_BoothP_14,
                   L1_1_L2_2_G1_MINI_ALU_BoothP_13,
                   L1_1_L2_2_G1_MINI_ALU_BoothP_12,
                   L1_1_L2_2_G1_MINI_ALU_BoothP_11,
                   L1_1_L2_2_G1_MINI_ALU_BoothP_10,
                   L1_1_L2_2_G1_MINI_ALU_BoothP_9,L1_1_L2_2_G1_MINI_ALU_BoothP_8
                   ,L1_1_L2_2_G1_MINI_ALU_BoothP_7,
                   L1_1_L2_2_G1_MINI_ALU_BoothP_6,L1_1_L2_2_G1_MINI_ALU_BoothP_5
                   ,L1_1_L2_2_G1_MINI_ALU_BoothP_4,
                   L1_1_L2_2_G1_MINI_ALU_BoothP_3,L1_1_L2_2_G1_MINI_ALU_BoothP_2
                   ,L1_1_L2_2_G1_MINI_ALU_BoothP_1,
                   L1_1_L2_2_G1_MINI_ALU_BoothP_0}), .SelOperand (nx3280), .Operation (
                   L1_1_L2_2_G1_MINI_ALU_BoothXORCheck), .AdderResult ({
                   L1ResultsLarge_7__16,L1ResultsLarge_7__15,
                   L1ResultsLarge_7__14,L1ResultsLarge_7__13,
                   L1ResultsLarge_7__12,L1ResultsLarge_7__11,
                   L1ResultsLarge_7__10,L1ResultsLarge_7__9,L1ResultsLarge_7__8,
                   L1ResultsLarge_7__7,L1ResultsLarge_7__6,L1ResultsLarge_7__5,
                   L1ResultsLarge_7__4,L1ResultsLarge_7__3,L1ResultsLarge_7__2,
                   L1ResultsLarge_7__1,L1ResultsLarge_7__0}), .AdderBoothResult (
                   {\$dummy [245],L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_15,
                   L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_14,
                   L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_13,
                   L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_12,
                   L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_11,
                   L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_10,
                   L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_9,
                   L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_8,
                   L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_7,
                   L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_6,
                   L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_5,
                   L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_4,
                   L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_3,
                   L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_2,
                   L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_1,
                   L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_0})) ;
    booth_unit_17 L1_1_L2_2_G1_MINI_ALU_BOOTH_UNIT (.CLK (CLK), .RST (RST), .Start (
                  Start), .Instr (Instr), .LoopingAndResultNotReady (nx3274), .Filter (
                  {FilterDin_1__2__7,FilterDin_1__2__6,FilterDin_1__2__5,
                  FilterDin_1__2__4,FilterDin_1__2__3,FilterDin_1__2__2,
                  FilterDin_1__2__1,FilterDin_1__2__0}), .Window ({
                  WindowDin_1__2__7,WindowDin_1__2__6,WindowDin_1__2__5,
                  WindowDin_1__2__4,WindowDin_1__2__3,WindowDin_1__2__2,
                  WindowDin_1__2__1,WindowDin_1__2__0}), .AdderBoothResult ({
                  L1FirstOperands_12__16,
                  L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_15,
                  L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_14,
                  L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_13,
                  L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_12,
                  L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_11,
                  L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_10,
                  L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_9,
                  L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_8,
                  L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_7,
                  L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_6,
                  L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_5,
                  L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_4,
                  L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_3,
                  L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_2,
                  L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_1,
                  L1_1_L2_2_G1_MINI_ALU_AdderBoothResult_0}), .BoothXORCheck (
                  L1_1_L2_2_G1_MINI_ALU_BoothXORCheck), .BoothResult ({
                  \$dummy [246],\$dummy [247],\$dummy [248],\$dummy [249],
                  \$dummy [250],\$dummy [251],\$dummy [252],\$dummy [253]}), .BoothAddingOperand (
                  {L1_1_L2_2_G1_MINI_ALU_BoothOperand_16,
                  L1_1_L2_2_G1_MINI_ALU_BoothOperand_15,
                  L1_1_L2_2_G1_MINI_ALU_BoothOperand_14,
                  L1_1_L2_2_G1_MINI_ALU_BoothOperand_13,
                  L1_1_L2_2_G1_MINI_ALU_BoothOperand_12,
                  L1_1_L2_2_G1_MINI_ALU_BoothOperand_11,
                  L1_1_L2_2_G1_MINI_ALU_BoothOperand_10,
                  L1_1_L2_2_G1_MINI_ALU_BoothOperand_9,\$dummy [254],
                  \$dummy [255],\$dummy [256],\$dummy [257],\$dummy [258],
                  \$dummy [259],\$dummy [260],\$dummy [261],\$dummy [262]}), .BoothP (
                  {L1_1_L2_2_G1_MINI_ALU_BoothP_16,
                  L1_1_L2_2_G1_MINI_ALU_BoothP_15,
                  L1_1_L2_2_G1_MINI_ALU_BoothP_14,
                  L1_1_L2_2_G1_MINI_ALU_BoothP_13,
                  L1_1_L2_2_G1_MINI_ALU_BoothP_12,
                  L1_1_L2_2_G1_MINI_ALU_BoothP_11,
                  L1_1_L2_2_G1_MINI_ALU_BoothP_10,L1_1_L2_2_G1_MINI_ALU_BoothP_9
                  ,L1_1_L2_2_G1_MINI_ALU_BoothP_8,L1_1_L2_2_G1_MINI_ALU_BoothP_7
                  ,L1_1_L2_2_G1_MINI_ALU_BoothP_6,L1_1_L2_2_G1_MINI_ALU_BoothP_5
                  ,L1_1_L2_2_G1_MINI_ALU_BoothP_4,L1_1_L2_2_G1_MINI_ALU_BoothP_3
                  ,L1_1_L2_2_G1_MINI_ALU_BoothP_2,L1_1_L2_2_G1_MINI_ALU_BoothP_1
                  ,L1_1_L2_2_G1_MINI_ALU_BoothP_0}), .LargeWindowShifted ({
                  \$dummy [263],\$dummy [264],\$dummy [265],\$dummy [266],
                  \$dummy [267],\$dummy [268],\$dummy [269],\$dummy [270],
                  \$dummy [271],\$dummy [272],\$dummy [273],\$dummy [274],
                  \$dummy [275],\$dummy [276],\$dummy [277],\$dummy [278],
                  \$dummy [279]})) ;
    booth_adder_17 L1_1_L2_3_G1_MINI_ALU_BOOTH_ADDER (.AdderFirstOperand ({
                   L1FirstOperands_12__16,L1FirstOperands_8__15,
                   L1FirstOperands_8__14,L1FirstOperands_8__13,
                   L1FirstOperands_8__12,L1FirstOperands_8__11,
                   L1FirstOperands_8__10,L1FirstOperands_8__9,
                   L1FirstOperands_8__8,L1FirstOperands_8__7,
                   L1FirstOperands_8__6,L1FirstOperands_8__5,
                   L1FirstOperands_8__4,L1FirstOperands_8__3,
                   L1FirstOperands_8__2,L1FirstOperands_8__1,
                   L1FirstOperands_8__0}), .AdderSecondOperand ({
                   L1FirstOperands_12__16,
                   L1_1_L2_3_G1_MINI_ALU_OperationResult_15,
                   L1_1_L2_3_G1_MINI_ALU_OperationResult_14,
                   L1_1_L2_3_G1_MINI_ALU_OperationResult_13,
                   L1_1_L2_3_G1_MINI_ALU_OperationResult_12,
                   L1_1_L2_3_G1_MINI_ALU_OperationResult_11,
                   L1_1_L2_3_G1_MINI_ALU_OperationResult_10,
                   L1_1_L2_3_G1_MINI_ALU_OperationResult_9,
                   L1_1_L2_3_G1_MINI_ALU_OperationResult_8,
                   L1_1_L2_3_G1_MINI_ALU_OperationResult_7,
                   L1_1_L2_3_G1_MINI_ALU_OperationResult_6,
                   L1_1_L2_3_G1_MINI_ALU_OperationResult_5,
                   L1_1_L2_3_G1_MINI_ALU_OperationResult_4,
                   L1_1_L2_3_G1_MINI_ALU_OperationResult_3,
                   L1_1_L2_3_G1_MINI_ALU_OperationResult_2,
                   L1_1_L2_3_G1_MINI_ALU_OperationResult_1,
                   L1_1_L2_3_G1_MINI_ALU_OperationResult_0}), .BoothOperand ({
                   L1_1_L2_3_G1_MINI_ALU_BoothOperand_16,
                   L1_1_L2_3_G1_MINI_ALU_BoothOperand_15,
                   L1_1_L2_3_G1_MINI_ALU_BoothOperand_14,
                   L1_1_L2_3_G1_MINI_ALU_BoothOperand_13,
                   L1_1_L2_3_G1_MINI_ALU_BoothOperand_12,
                   L1_1_L2_3_G1_MINI_ALU_BoothOperand_11,
                   L1_1_L2_3_G1_MINI_ALU_BoothOperand_10,
                   L1_1_L2_3_G1_MINI_ALU_BoothOperand_9,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16}), .BoothP ({
                   L1_1_L2_3_G1_MINI_ALU_BoothP_16,
                   L1_1_L2_3_G1_MINI_ALU_BoothP_15,
                   L1_1_L2_3_G1_MINI_ALU_BoothP_14,
                   L1_1_L2_3_G1_MINI_ALU_BoothP_13,
                   L1_1_L2_3_G1_MINI_ALU_BoothP_12,
                   L1_1_L2_3_G1_MINI_ALU_BoothP_11,
                   L1_1_L2_3_G1_MINI_ALU_BoothP_10,
                   L1_1_L2_3_G1_MINI_ALU_BoothP_9,L1_1_L2_3_G1_MINI_ALU_BoothP_8
                   ,L1_1_L2_3_G1_MINI_ALU_BoothP_7,
                   L1_1_L2_3_G1_MINI_ALU_BoothP_6,L1_1_L2_3_G1_MINI_ALU_BoothP_5
                   ,L1_1_L2_3_G1_MINI_ALU_BoothP_4,
                   L1_1_L2_3_G1_MINI_ALU_BoothP_3,L1_1_L2_3_G1_MINI_ALU_BoothP_2
                   ,L1_1_L2_3_G1_MINI_ALU_BoothP_1,
                   L1_1_L2_3_G1_MINI_ALU_BoothP_0}), .SelOperand (nx3282), .Operation (
                   L1_1_L2_3_G1_MINI_ALU_BoothXORCheck), .AdderResult ({
                   L1ResultsLarge_8__16,L1ResultsLarge_8__15,
                   L1ResultsLarge_8__14,L1ResultsLarge_8__13,
                   L1ResultsLarge_8__12,L1ResultsLarge_8__11,
                   L1ResultsLarge_8__10,L1ResultsLarge_8__9,L1ResultsLarge_8__8,
                   L1ResultsLarge_8__7,L1ResultsLarge_8__6,L1ResultsLarge_8__5,
                   L1ResultsLarge_8__4,L1ResultsLarge_8__3,L1ResultsLarge_8__2,
                   L1ResultsLarge_8__1,L1ResultsLarge_8__0}), .AdderBoothResult (
                   {\$dummy [280],L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_15,
                   L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_14,
                   L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_13,
                   L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_12,
                   L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_11,
                   L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_10,
                   L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_9,
                   L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_8,
                   L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_7,
                   L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_6,
                   L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_5,
                   L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_4,
                   L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_3,
                   L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_2,
                   L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_1,
                   L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_0})) ;
    booth_unit_17 L1_1_L2_3_G1_MINI_ALU_BOOTH_UNIT (.CLK (CLK), .RST (RST), .Start (
                  Start), .Instr (Instr), .LoopingAndResultNotReady (nx3274), .Filter (
                  {FilterDin_1__3__7,FilterDin_1__3__6,FilterDin_1__3__5,
                  FilterDin_1__3__4,FilterDin_1__3__3,FilterDin_1__3__2,
                  FilterDin_1__3__1,FilterDin_1__3__0}), .Window ({
                  WindowDin_1__3__7,WindowDin_1__3__6,WindowDin_1__3__5,
                  WindowDin_1__3__4,WindowDin_1__3__3,WindowDin_1__3__2,
                  WindowDin_1__3__1,WindowDin_1__3__0}), .AdderBoothResult ({
                  L1FirstOperands_12__16,
                  L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_15,
                  L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_14,
                  L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_13,
                  L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_12,
                  L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_11,
                  L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_10,
                  L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_9,
                  L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_8,
                  L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_7,
                  L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_6,
                  L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_5,
                  L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_4,
                  L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_3,
                  L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_2,
                  L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_1,
                  L1_1_L2_3_G1_MINI_ALU_AdderBoothResult_0}), .BoothXORCheck (
                  L1_1_L2_3_G1_MINI_ALU_BoothXORCheck), .BoothResult ({
                  \$dummy [281],\$dummy [282],\$dummy [283],\$dummy [284],
                  \$dummy [285],\$dummy [286],\$dummy [287],\$dummy [288]}), .BoothAddingOperand (
                  {L1_1_L2_3_G1_MINI_ALU_BoothOperand_16,
                  L1_1_L2_3_G1_MINI_ALU_BoothOperand_15,
                  L1_1_L2_3_G1_MINI_ALU_BoothOperand_14,
                  L1_1_L2_3_G1_MINI_ALU_BoothOperand_13,
                  L1_1_L2_3_G1_MINI_ALU_BoothOperand_12,
                  L1_1_L2_3_G1_MINI_ALU_BoothOperand_11,
                  L1_1_L2_3_G1_MINI_ALU_BoothOperand_10,
                  L1_1_L2_3_G1_MINI_ALU_BoothOperand_9,\$dummy [289],
                  \$dummy [290],\$dummy [291],\$dummy [292],\$dummy [293],
                  \$dummy [294],\$dummy [295],\$dummy [296],\$dummy [297]}), .BoothP (
                  {L1_1_L2_3_G1_MINI_ALU_BoothP_16,
                  L1_1_L2_3_G1_MINI_ALU_BoothP_15,
                  L1_1_L2_3_G1_MINI_ALU_BoothP_14,
                  L1_1_L2_3_G1_MINI_ALU_BoothP_13,
                  L1_1_L2_3_G1_MINI_ALU_BoothP_12,
                  L1_1_L2_3_G1_MINI_ALU_BoothP_11,
                  L1_1_L2_3_G1_MINI_ALU_BoothP_10,L1_1_L2_3_G1_MINI_ALU_BoothP_9
                  ,L1_1_L2_3_G1_MINI_ALU_BoothP_8,L1_1_L2_3_G1_MINI_ALU_BoothP_7
                  ,L1_1_L2_3_G1_MINI_ALU_BoothP_6,L1_1_L2_3_G1_MINI_ALU_BoothP_5
                  ,L1_1_L2_3_G1_MINI_ALU_BoothP_4,L1_1_L2_3_G1_MINI_ALU_BoothP_3
                  ,L1_1_L2_3_G1_MINI_ALU_BoothP_2,L1_1_L2_3_G1_MINI_ALU_BoothP_1
                  ,L1_1_L2_3_G1_MINI_ALU_BoothP_0}), .LargeWindowShifted ({
                  \$dummy [298],\$dummy [299],\$dummy [300],\$dummy [301],
                  \$dummy [302],\$dummy [303],\$dummy [304],\$dummy [305],
                  \$dummy [306],\$dummy [307],\$dummy [308],\$dummy [309],
                  \$dummy [310],\$dummy [311],\$dummy [312],\$dummy [313],
                  \$dummy [314]})) ;
    booth_adder_17 L1_1_L2_4_G1_MINI_ALU_BOOTH_ADDER (.AdderFirstOperand ({
                   L1FirstOperands_12__16,L1FirstOperands_4__15,
                   L1FirstOperands_4__14,L1FirstOperands_4__13,
                   L1FirstOperands_4__12,L1FirstOperands_4__11,
                   L1FirstOperands_4__10,L1FirstOperands_4__9,
                   L1FirstOperands_4__8,L1FirstOperands_4__7,
                   L1FirstOperands_4__6,L1FirstOperands_4__5,
                   L1FirstOperands_4__4,L1FirstOperands_4__3,
                   L1FirstOperands_4__2,L1FirstOperands_4__1,
                   L1FirstOperands_4__0}), .AdderSecondOperand ({
                   L1FirstOperands_12__16,
                   L1_1_L2_4_G1_MINI_ALU_OperationResult_15,
                   L1_1_L2_4_G1_MINI_ALU_OperationResult_14,
                   L1_1_L2_4_G1_MINI_ALU_OperationResult_13,
                   L1_1_L2_4_G1_MINI_ALU_OperationResult_12,
                   L1_1_L2_4_G1_MINI_ALU_OperationResult_11,
                   L1_1_L2_4_G1_MINI_ALU_OperationResult_10,
                   L1_1_L2_4_G1_MINI_ALU_OperationResult_9,
                   L1_1_L2_4_G1_MINI_ALU_OperationResult_8,
                   L1_1_L2_4_G1_MINI_ALU_OperationResult_7,
                   L1_1_L2_4_G1_MINI_ALU_OperationResult_6,
                   L1_1_L2_4_G1_MINI_ALU_OperationResult_5,
                   L1_1_L2_4_G1_MINI_ALU_OperationResult_4,
                   L1_1_L2_4_G1_MINI_ALU_OperationResult_3,
                   L1_1_L2_4_G1_MINI_ALU_OperationResult_2,
                   L1_1_L2_4_G1_MINI_ALU_OperationResult_1,
                   L1_1_L2_4_G1_MINI_ALU_OperationResult_0}), .BoothOperand ({
                   L1_1_L2_4_G1_MINI_ALU_BoothOperand_16,
                   L1_1_L2_4_G1_MINI_ALU_BoothOperand_15,
                   L1_1_L2_4_G1_MINI_ALU_BoothOperand_14,
                   L1_1_L2_4_G1_MINI_ALU_BoothOperand_13,
                   L1_1_L2_4_G1_MINI_ALU_BoothOperand_12,
                   L1_1_L2_4_G1_MINI_ALU_BoothOperand_11,
                   L1_1_L2_4_G1_MINI_ALU_BoothOperand_10,
                   L1_1_L2_4_G1_MINI_ALU_BoothOperand_9,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16}), .BoothP ({
                   L1_1_L2_4_G1_MINI_ALU_BoothP_16,
                   L1_1_L2_4_G1_MINI_ALU_BoothP_15,
                   L1_1_L2_4_G1_MINI_ALU_BoothP_14,
                   L1_1_L2_4_G1_MINI_ALU_BoothP_13,
                   L1_1_L2_4_G1_MINI_ALU_BoothP_12,
                   L1_1_L2_4_G1_MINI_ALU_BoothP_11,
                   L1_1_L2_4_G1_MINI_ALU_BoothP_10,
                   L1_1_L2_4_G1_MINI_ALU_BoothP_9,L1_1_L2_4_G1_MINI_ALU_BoothP_8
                   ,L1_1_L2_4_G1_MINI_ALU_BoothP_7,
                   L1_1_L2_4_G1_MINI_ALU_BoothP_6,L1_1_L2_4_G1_MINI_ALU_BoothP_5
                   ,L1_1_L2_4_G1_MINI_ALU_BoothP_4,
                   L1_1_L2_4_G1_MINI_ALU_BoothP_3,L1_1_L2_4_G1_MINI_ALU_BoothP_2
                   ,L1_1_L2_4_G1_MINI_ALU_BoothP_1,
                   L1_1_L2_4_G1_MINI_ALU_BoothP_0}), .SelOperand (nx3282), .Operation (
                   L1_1_L2_4_G1_MINI_ALU_BoothXORCheck), .AdderResult ({
                   L1ResultsLarge_9__16,L1ResultsLarge_9__15,
                   L1ResultsLarge_9__14,L1ResultsLarge_9__13,
                   L1ResultsLarge_9__12,L1ResultsLarge_9__11,
                   L1ResultsLarge_9__10,L1ResultsLarge_9__9,L1ResultsLarge_9__8,
                   L1ResultsLarge_9__7,L1ResultsLarge_9__6,L1ResultsLarge_9__5,
                   L1ResultsLarge_9__4,L1ResultsLarge_9__3,L1ResultsLarge_9__2,
                   L1ResultsLarge_9__1,L1ResultsLarge_9__0}), .AdderBoothResult (
                   {\$dummy [315],L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_15,
                   L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_14,
                   L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_13,
                   L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_12,
                   L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_11,
                   L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_10,
                   L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_9,
                   L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_8,
                   L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_7,
                   L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_6,
                   L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_5,
                   L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_4,
                   L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_3,
                   L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_2,
                   L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_1,
                   L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_0})) ;
    booth_unit_17 L1_1_L2_4_G1_MINI_ALU_BOOTH_UNIT (.CLK (CLK), .RST (RST), .Start (
                  Start), .Instr (Instr), .LoopingAndResultNotReady (nx3274), .Filter (
                  {FilterDin_1__4__7,FilterDin_1__4__6,FilterDin_1__4__5,
                  FilterDin_1__4__4,FilterDin_1__4__3,FilterDin_1__4__2,
                  FilterDin_1__4__1,FilterDin_1__4__0}), .Window ({
                  WindowDin_1__4__7,WindowDin_1__4__6,WindowDin_1__4__5,
                  WindowDin_1__4__4,WindowDin_1__4__3,WindowDin_1__4__2,
                  WindowDin_1__4__1,WindowDin_1__4__0}), .AdderBoothResult ({
                  L1FirstOperands_12__16,
                  L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_15,
                  L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_14,
                  L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_13,
                  L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_12,
                  L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_11,
                  L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_10,
                  L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_9,
                  L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_8,
                  L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_7,
                  L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_6,
                  L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_5,
                  L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_4,
                  L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_3,
                  L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_2,
                  L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_1,
                  L1_1_L2_4_G1_MINI_ALU_AdderBoothResult_0}), .BoothXORCheck (
                  L1_1_L2_4_G1_MINI_ALU_BoothXORCheck), .BoothResult ({
                  \$dummy [316],\$dummy [317],\$dummy [318],\$dummy [319],
                  \$dummy [320],\$dummy [321],\$dummy [322],\$dummy [323]}), .BoothAddingOperand (
                  {L1_1_L2_4_G1_MINI_ALU_BoothOperand_16,
                  L1_1_L2_4_G1_MINI_ALU_BoothOperand_15,
                  L1_1_L2_4_G1_MINI_ALU_BoothOperand_14,
                  L1_1_L2_4_G1_MINI_ALU_BoothOperand_13,
                  L1_1_L2_4_G1_MINI_ALU_BoothOperand_12,
                  L1_1_L2_4_G1_MINI_ALU_BoothOperand_11,
                  L1_1_L2_4_G1_MINI_ALU_BoothOperand_10,
                  L1_1_L2_4_G1_MINI_ALU_BoothOperand_9,\$dummy [324],
                  \$dummy [325],\$dummy [326],\$dummy [327],\$dummy [328],
                  \$dummy [329],\$dummy [330],\$dummy [331],\$dummy [332]}), .BoothP (
                  {L1_1_L2_4_G1_MINI_ALU_BoothP_16,
                  L1_1_L2_4_G1_MINI_ALU_BoothP_15,
                  L1_1_L2_4_G1_MINI_ALU_BoothP_14,
                  L1_1_L2_4_G1_MINI_ALU_BoothP_13,
                  L1_1_L2_4_G1_MINI_ALU_BoothP_12,
                  L1_1_L2_4_G1_MINI_ALU_BoothP_11,
                  L1_1_L2_4_G1_MINI_ALU_BoothP_10,L1_1_L2_4_G1_MINI_ALU_BoothP_9
                  ,L1_1_L2_4_G1_MINI_ALU_BoothP_8,L1_1_L2_4_G1_MINI_ALU_BoothP_7
                  ,L1_1_L2_4_G1_MINI_ALU_BoothP_6,L1_1_L2_4_G1_MINI_ALU_BoothP_5
                  ,L1_1_L2_4_G1_MINI_ALU_BoothP_4,L1_1_L2_4_G1_MINI_ALU_BoothP_3
                  ,L1_1_L2_4_G1_MINI_ALU_BoothP_2,L1_1_L2_4_G1_MINI_ALU_BoothP_1
                  ,L1_1_L2_4_G1_MINI_ALU_BoothP_0}), .LargeWindowShifted ({
                  \$dummy [333],\$dummy [334],\$dummy [335],\$dummy [336],
                  \$dummy [337],\$dummy [338],\$dummy [339],\$dummy [340],
                  \$dummy [341],\$dummy [342],\$dummy [343],\$dummy [344],
                  \$dummy [345],\$dummy [346],\$dummy [347],\$dummy [348],
                  \$dummy [349]})) ;
    booth_adder_17 L1_2_L2_0_G1_MINI_ALU_BOOTH_ADDER (.AdderFirstOperand ({
                   L1FirstOperands_12__16,L1FirstOperands_10__15,
                   L1FirstOperands_10__14,L1FirstOperands_10__13,
                   L1FirstOperands_10__12,L1FirstOperands_10__11,
                   L1FirstOperands_10__10,L1FirstOperands_10__9,
                   L1FirstOperands_10__8,L1FirstOperands_10__7,
                   L1FirstOperands_10__6,L1FirstOperands_10__5,
                   L1FirstOperands_10__4,L1FirstOperands_10__3,
                   L1FirstOperands_10__2,L1FirstOperands_10__1,
                   L1FirstOperands_10__0}), .AdderSecondOperand ({
                   L1FirstOperands_12__16,
                   L1_2_L2_0_G1_MINI_ALU_OperationResult_15,
                   L1_2_L2_0_G1_MINI_ALU_OperationResult_14,
                   L1_2_L2_0_G1_MINI_ALU_OperationResult_13,
                   L1_2_L2_0_G1_MINI_ALU_OperationResult_12,
                   L1_2_L2_0_G1_MINI_ALU_OperationResult_11,
                   L1_2_L2_0_G1_MINI_ALU_OperationResult_10,
                   L1_2_L2_0_G1_MINI_ALU_OperationResult_9,
                   L1_2_L2_0_G1_MINI_ALU_OperationResult_8,
                   L1_2_L2_0_G1_MINI_ALU_OperationResult_7,
                   L1_2_L2_0_G1_MINI_ALU_OperationResult_6,
                   L1_2_L2_0_G1_MINI_ALU_OperationResult_5,
                   L1_2_L2_0_G1_MINI_ALU_OperationResult_4,
                   L1_2_L2_0_G1_MINI_ALU_OperationResult_3,
                   L1_2_L2_0_G1_MINI_ALU_OperationResult_2,
                   L1_2_L2_0_G1_MINI_ALU_OperationResult_1,
                   L1_2_L2_0_G1_MINI_ALU_OperationResult_0}), .BoothOperand ({
                   L1_2_L2_0_G1_MINI_ALU_BoothOperand_16,
                   L1_2_L2_0_G1_MINI_ALU_BoothOperand_15,
                   L1_2_L2_0_G1_MINI_ALU_BoothOperand_14,
                   L1_2_L2_0_G1_MINI_ALU_BoothOperand_13,
                   L1_2_L2_0_G1_MINI_ALU_BoothOperand_12,
                   L1_2_L2_0_G1_MINI_ALU_BoothOperand_11,
                   L1_2_L2_0_G1_MINI_ALU_BoothOperand_10,
                   L1_2_L2_0_G1_MINI_ALU_BoothOperand_9,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16}), .BoothP ({
                   L1_2_L2_0_G1_MINI_ALU_BoothP_16,
                   L1_2_L2_0_G1_MINI_ALU_BoothP_15,
                   L1_2_L2_0_G1_MINI_ALU_BoothP_14,
                   L1_2_L2_0_G1_MINI_ALU_BoothP_13,
                   L1_2_L2_0_G1_MINI_ALU_BoothP_12,
                   L1_2_L2_0_G1_MINI_ALU_BoothP_11,
                   L1_2_L2_0_G1_MINI_ALU_BoothP_10,
                   L1_2_L2_0_G1_MINI_ALU_BoothP_9,L1_2_L2_0_G1_MINI_ALU_BoothP_8
                   ,L1_2_L2_0_G1_MINI_ALU_BoothP_7,
                   L1_2_L2_0_G1_MINI_ALU_BoothP_6,L1_2_L2_0_G1_MINI_ALU_BoothP_5
                   ,L1_2_L2_0_G1_MINI_ALU_BoothP_4,
                   L1_2_L2_0_G1_MINI_ALU_BoothP_3,L1_2_L2_0_G1_MINI_ALU_BoothP_2
                   ,L1_2_L2_0_G1_MINI_ALU_BoothP_1,
                   L1_2_L2_0_G1_MINI_ALU_BoothP_0}), .SelOperand (nx3282), .Operation (
                   L1_2_L2_0_G1_MINI_ALU_BoothXORCheck), .AdderResult ({
                   L1ResultsLarge_10__16,L1ResultsLarge_10__15,
                   L1ResultsLarge_10__14,L1ResultsLarge_10__13,
                   L1ResultsLarge_10__12,L1ResultsLarge_10__11,
                   L1ResultsLarge_10__10,L1ResultsLarge_10__9,
                   L1ResultsLarge_10__8,L1ResultsLarge_10__7,
                   L1ResultsLarge_10__6,L1ResultsLarge_10__5,
                   L1ResultsLarge_10__4,L1ResultsLarge_10__3,
                   L1ResultsLarge_10__2,L1ResultsLarge_10__1,
                   L1ResultsLarge_10__0}), .AdderBoothResult ({\$dummy [350],
                   L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_15,
                   L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_14,
                   L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_13,
                   L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_12,
                   L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_11,
                   L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_10,
                   L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_9,
                   L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_8,
                   L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_7,
                   L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_6,
                   L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_5,
                   L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_4,
                   L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_3,
                   L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_2,
                   L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_1,
                   L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_0})) ;
    booth_unit_17 L1_2_L2_0_G1_MINI_ALU_BOOTH_UNIT (.CLK (CLK), .RST (RST), .Start (
                  Start), .Instr (Instr), .LoopingAndResultNotReady (nx3274), .Filter (
                  {FilterDin_2__0__7,FilterDin_2__0__6,FilterDin_2__0__5,
                  FilterDin_2__0__4,FilterDin_2__0__3,FilterDin_2__0__2,
                  FilterDin_2__0__1,FilterDin_2__0__0}), .Window ({
                  WindowDin_2__0__7,WindowDin_2__0__6,WindowDin_2__0__5,
                  WindowDin_2__0__4,WindowDin_2__0__3,WindowDin_2__0__2,
                  WindowDin_2__0__1,WindowDin_2__0__0}), .AdderBoothResult ({
                  L1FirstOperands_12__16,
                  L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_15,
                  L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_14,
                  L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_13,
                  L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_12,
                  L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_11,
                  L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_10,
                  L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_9,
                  L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_8,
                  L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_7,
                  L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_6,
                  L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_5,
                  L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_4,
                  L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_3,
                  L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_2,
                  L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_1,
                  L1_2_L2_0_G1_MINI_ALU_AdderBoothResult_0}), .BoothXORCheck (
                  L1_2_L2_0_G1_MINI_ALU_BoothXORCheck), .BoothResult ({
                  \$dummy [351],\$dummy [352],\$dummy [353],\$dummy [354],
                  \$dummy [355],\$dummy [356],\$dummy [357],\$dummy [358]}), .BoothAddingOperand (
                  {L1_2_L2_0_G1_MINI_ALU_BoothOperand_16,
                  L1_2_L2_0_G1_MINI_ALU_BoothOperand_15,
                  L1_2_L2_0_G1_MINI_ALU_BoothOperand_14,
                  L1_2_L2_0_G1_MINI_ALU_BoothOperand_13,
                  L1_2_L2_0_G1_MINI_ALU_BoothOperand_12,
                  L1_2_L2_0_G1_MINI_ALU_BoothOperand_11,
                  L1_2_L2_0_G1_MINI_ALU_BoothOperand_10,
                  L1_2_L2_0_G1_MINI_ALU_BoothOperand_9,\$dummy [359],
                  \$dummy [360],\$dummy [361],\$dummy [362],\$dummy [363],
                  \$dummy [364],\$dummy [365],\$dummy [366],\$dummy [367]}), .BoothP (
                  {L1_2_L2_0_G1_MINI_ALU_BoothP_16,
                  L1_2_L2_0_G1_MINI_ALU_BoothP_15,
                  L1_2_L2_0_G1_MINI_ALU_BoothP_14,
                  L1_2_L2_0_G1_MINI_ALU_BoothP_13,
                  L1_2_L2_0_G1_MINI_ALU_BoothP_12,
                  L1_2_L2_0_G1_MINI_ALU_BoothP_11,
                  L1_2_L2_0_G1_MINI_ALU_BoothP_10,L1_2_L2_0_G1_MINI_ALU_BoothP_9
                  ,L1_2_L2_0_G1_MINI_ALU_BoothP_8,L1_2_L2_0_G1_MINI_ALU_BoothP_7
                  ,L1_2_L2_0_G1_MINI_ALU_BoothP_6,L1_2_L2_0_G1_MINI_ALU_BoothP_5
                  ,L1_2_L2_0_G1_MINI_ALU_BoothP_4,L1_2_L2_0_G1_MINI_ALU_BoothP_3
                  ,L1_2_L2_0_G1_MINI_ALU_BoothP_2,L1_2_L2_0_G1_MINI_ALU_BoothP_1
                  ,L1_2_L2_0_G1_MINI_ALU_BoothP_0}), .LargeWindowShifted ({
                  \$dummy [368],\$dummy [369],\$dummy [370],\$dummy [371],
                  \$dummy [372],\$dummy [373],\$dummy [374],\$dummy [375],
                  \$dummy [376],\$dummy [377],\$dummy [378],\$dummy [379],
                  \$dummy [380],\$dummy [381],\$dummy [382],\$dummy [383],
                  \$dummy [384]})) ;
    booth_adder_17 L1_2_L2_1_G1_MINI_ALU_BOOTH_ADDER (.AdderFirstOperand ({
                   L1FirstOperands_12__16,L1FirstOperands_11__15,
                   L1FirstOperands_11__14,L1FirstOperands_11__13,
                   L1FirstOperands_11__12,L1FirstOperands_11__11,
                   L1FirstOperands_11__10,L1FirstOperands_11__9,
                   L1FirstOperands_11__8,L1FirstOperands_11__7,
                   L1FirstOperands_11__6,L1FirstOperands_11__5,
                   L1FirstOperands_11__4,L1FirstOperands_11__3,
                   L1FirstOperands_11__2,L1FirstOperands_11__1,
                   L1FirstOperands_11__0}), .AdderSecondOperand ({
                   L1FirstOperands_12__16,
                   L1_2_L2_1_G1_MINI_ALU_OperationResult_15,
                   L1_2_L2_1_G1_MINI_ALU_OperationResult_14,
                   L1_2_L2_1_G1_MINI_ALU_OperationResult_13,
                   L1_2_L2_1_G1_MINI_ALU_OperationResult_12,
                   L1_2_L2_1_G1_MINI_ALU_OperationResult_11,
                   L1_2_L2_1_G1_MINI_ALU_OperationResult_10,
                   L1_2_L2_1_G1_MINI_ALU_OperationResult_9,
                   L1_2_L2_1_G1_MINI_ALU_OperationResult_8,
                   L1_2_L2_1_G1_MINI_ALU_OperationResult_7,
                   L1_2_L2_1_G1_MINI_ALU_OperationResult_6,
                   L1_2_L2_1_G1_MINI_ALU_OperationResult_5,
                   L1_2_L2_1_G1_MINI_ALU_OperationResult_4,
                   L1_2_L2_1_G1_MINI_ALU_OperationResult_3,
                   L1_2_L2_1_G1_MINI_ALU_OperationResult_2,
                   L1_2_L2_1_G1_MINI_ALU_OperationResult_1,
                   L1_2_L2_1_G1_MINI_ALU_OperationResult_0}), .BoothOperand ({
                   L1_2_L2_1_G1_MINI_ALU_BoothOperand_16,
                   L1_2_L2_1_G1_MINI_ALU_BoothOperand_15,
                   L1_2_L2_1_G1_MINI_ALU_BoothOperand_14,
                   L1_2_L2_1_G1_MINI_ALU_BoothOperand_13,
                   L1_2_L2_1_G1_MINI_ALU_BoothOperand_12,
                   L1_2_L2_1_G1_MINI_ALU_BoothOperand_11,
                   L1_2_L2_1_G1_MINI_ALU_BoothOperand_10,
                   L1_2_L2_1_G1_MINI_ALU_BoothOperand_9,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16,
                   L1FirstOperands_12__16,L1FirstOperands_12__16}), .BoothP ({
                   L1_2_L2_1_G1_MINI_ALU_BoothP_16,
                   L1_2_L2_1_G1_MINI_ALU_BoothP_15,
                   L1_2_L2_1_G1_MINI_ALU_BoothP_14,
                   L1_2_L2_1_G1_MINI_ALU_BoothP_13,
                   L1_2_L2_1_G1_MINI_ALU_BoothP_12,
                   L1_2_L2_1_G1_MINI_ALU_BoothP_11,
                   L1_2_L2_1_G1_MINI_ALU_BoothP_10,
                   L1_2_L2_1_G1_MINI_ALU_BoothP_9,L1_2_L2_1_G1_MINI_ALU_BoothP_8
                   ,L1_2_L2_1_G1_MINI_ALU_BoothP_7,
                   L1_2_L2_1_G1_MINI_ALU_BoothP_6,L1_2_L2_1_G1_MINI_ALU_BoothP_5
                   ,L1_2_L2_1_G1_MINI_ALU_BoothP_4,
                   L1_2_L2_1_G1_MINI_ALU_BoothP_3,L1_2_L2_1_G1_MINI_ALU_BoothP_2
                   ,L1_2_L2_1_G1_MINI_ALU_BoothP_1,
                   L1_2_L2_1_G1_MINI_ALU_BoothP_0}), .SelOperand (nx3282), .Operation (
                   L1_2_L2_1_G1_MINI_ALU_BoothXORCheck), .AdderResult ({
                   L1ResultsLarge_11__16,L1ResultsLarge_11__15,
                   L1ResultsLarge_11__14,L1ResultsLarge_11__13,
                   L1ResultsLarge_11__12,L1ResultsLarge_11__11,
                   L1ResultsLarge_11__10,L1ResultsLarge_11__9,
                   L1ResultsLarge_11__8,L1ResultsLarge_11__7,
                   L1ResultsLarge_11__6,L1ResultsLarge_11__5,
                   L1ResultsLarge_11__4,L1ResultsLarge_11__3,
                   L1ResultsLarge_11__2,L1ResultsLarge_11__1,
                   L1ResultsLarge_11__0}), .AdderBoothResult ({\$dummy [385],
                   L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_15,
                   L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_14,
                   L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_13,
                   L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_12,
                   L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_11,
                   L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_10,
                   L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_9,
                   L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_8,
                   L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_7,
                   L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_6,
                   L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_5,
                   L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_4,
                   L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_3,
                   L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_2,
                   L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_1,
                   L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_0})) ;
    booth_unit_17 L1_2_L2_1_G1_MINI_ALU_BOOTH_UNIT (.CLK (CLK), .RST (RST), .Start (
                  Start), .Instr (Instr), .LoopingAndResultNotReady (nx3274), .Filter (
                  {FilterDin_2__1__7,FilterDin_2__1__6,FilterDin_2__1__5,
                  FilterDin_2__1__4,FilterDin_2__1__3,FilterDin_2__1__2,
                  FilterDin_2__1__1,FilterDin_2__1__0}), .Window ({
                  WindowDin_2__1__7,WindowDin_2__1__6,WindowDin_2__1__5,
                  WindowDin_2__1__4,WindowDin_2__1__3,WindowDin_2__1__2,
                  WindowDin_2__1__1,WindowDin_2__1__0}), .AdderBoothResult ({
                  L1FirstOperands_12__16,
                  L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_15,
                  L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_14,
                  L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_13,
                  L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_12,
                  L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_11,
                  L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_10,
                  L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_9,
                  L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_8,
                  L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_7,
                  L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_6,
                  L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_5,
                  L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_4,
                  L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_3,
                  L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_2,
                  L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_1,
                  L1_2_L2_1_G1_MINI_ALU_AdderBoothResult_0}), .BoothXORCheck (
                  L1_2_L2_1_G1_MINI_ALU_BoothXORCheck), .BoothResult ({
                  \$dummy [386],\$dummy [387],\$dummy [388],\$dummy [389],
                  \$dummy [390],\$dummy [391],\$dummy [392],\$dummy [393]}), .BoothAddingOperand (
                  {L1_2_L2_1_G1_MINI_ALU_BoothOperand_16,
                  L1_2_L2_1_G1_MINI_ALU_BoothOperand_15,
                  L1_2_L2_1_G1_MINI_ALU_BoothOperand_14,
                  L1_2_L2_1_G1_MINI_ALU_BoothOperand_13,
                  L1_2_L2_1_G1_MINI_ALU_BoothOperand_12,
                  L1_2_L2_1_G1_MINI_ALU_BoothOperand_11,
                  L1_2_L2_1_G1_MINI_ALU_BoothOperand_10,
                  L1_2_L2_1_G1_MINI_ALU_BoothOperand_9,\$dummy [394],
                  \$dummy [395],\$dummy [396],\$dummy [397],\$dummy [398],
                  \$dummy [399],\$dummy [400],\$dummy [401],\$dummy [402]}), .BoothP (
                  {L1_2_L2_1_G1_MINI_ALU_BoothP_16,
                  L1_2_L2_1_G1_MINI_ALU_BoothP_15,
                  L1_2_L2_1_G1_MINI_ALU_BoothP_14,
                  L1_2_L2_1_G1_MINI_ALU_BoothP_13,
                  L1_2_L2_1_G1_MINI_ALU_BoothP_12,
                  L1_2_L2_1_G1_MINI_ALU_BoothP_11,
                  L1_2_L2_1_G1_MINI_ALU_BoothP_10,L1_2_L2_1_G1_MINI_ALU_BoothP_9
                  ,L1_2_L2_1_G1_MINI_ALU_BoothP_8,L1_2_L2_1_G1_MINI_ALU_BoothP_7
                  ,L1_2_L2_1_G1_MINI_ALU_BoothP_6,L1_2_L2_1_G1_MINI_ALU_BoothP_5
                  ,L1_2_L2_1_G1_MINI_ALU_BoothP_4,L1_2_L2_1_G1_MINI_ALU_BoothP_3
                  ,L1_2_L2_1_G1_MINI_ALU_BoothP_2,L1_2_L2_1_G1_MINI_ALU_BoothP_1
                  ,L1_2_L2_1_G1_MINI_ALU_BoothP_0}), .LargeWindowShifted ({
                  \$dummy [403],\$dummy [404],\$dummy [405],\$dummy [406],
                  \$dummy [407],\$dummy [408],\$dummy [409],\$dummy [410],
                  \$dummy [411],\$dummy [412],\$dummy [413],\$dummy [414],
                  \$dummy [415],\$dummy [416],\$dummy [417],\$dummy [418],
                  \$dummy [419]})) ;
    booth_adder_17_unfolded15 L1_2_L2_2_G1_MINI_ALU_BOOTH_ADDER (.AdderFirstOperand (
                              {L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16}), .AdderSecondOperand ({
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16}), .BoothOperand ({
                              L1_2_L2_2_G1_MINI_ALU_BoothOperand_16,
                              L1_2_L2_2_G1_MINI_ALU_BoothOperand_15,
                              L1_2_L2_2_G1_MINI_ALU_BoothOperand_14,
                              L1_2_L2_2_G1_MINI_ALU_BoothOperand_13,
                              L1_2_L2_2_G1_MINI_ALU_BoothOperand_12,
                              L1_2_L2_2_G1_MINI_ALU_BoothOperand_11,
                              L1_2_L2_2_G1_MINI_ALU_BoothOperand_10,
                              L1_2_L2_2_G1_MINI_ALU_BoothOperand_9,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16}), .BoothP ({
                              L1_2_L2_2_G1_MINI_ALU_BoothP_16,
                              L1_2_L2_2_G1_MINI_ALU_BoothP_15,
                              L1_2_L2_2_G1_MINI_ALU_BoothP_14,
                              L1_2_L2_2_G1_MINI_ALU_BoothP_13,
                              L1_2_L2_2_G1_MINI_ALU_BoothP_12,
                              L1_2_L2_2_G1_MINI_ALU_BoothP_11,
                              L1_2_L2_2_G1_MINI_ALU_BoothP_10,
                              L1_2_L2_2_G1_MINI_ALU_BoothP_9,
                              L1_2_L2_2_G1_MINI_ALU_BoothP_8,
                              L1_2_L2_2_G1_MINI_ALU_BoothP_7,
                              L1_2_L2_2_G1_MINI_ALU_BoothP_6,
                              L1_2_L2_2_G1_MINI_ALU_BoothP_5,
                              L1_2_L2_2_G1_MINI_ALU_BoothP_4,
                              L1_2_L2_2_G1_MINI_ALU_BoothP_3,
                              L1_2_L2_2_G1_MINI_ALU_BoothP_2,
                              L1_2_L2_2_G1_MINI_ALU_BoothP_1,
                              L1FirstOperands_12__16}), .SelOperand (nx3280), .Operation (
                              L1_2_L2_2_G1_MINI_ALU_BoothXORCheck), .AdderResult (
                              {\$dummy [420],\$dummy [421],\$dummy [422],
                              \$dummy [423],\$dummy [424],\$dummy [425],
                              \$dummy [426],\$dummy [427],\$dummy [428],
                              \$dummy [429],\$dummy [430],\$dummy [431],
                              \$dummy [432],\$dummy [433],\$dummy [434],
                              \$dummy [435],\$dummy [436]}), .AdderBoothResult (
                              {\$dummy [437],
                              L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_15,
                              L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_14,
                              L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_13,
                              L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_12,
                              L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_11,
                              L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_10,
                              L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_9,
                              L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_8,
                              L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_7,
                              L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_6,
                              L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_5,
                              L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_4,
                              L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_3,
                              L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_2,
                              L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_1,
                              L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_0})) ;
    booth_unit_17_unfolded5 L1_2_L2_2_G1_MINI_ALU_BOOTH_UNIT (.CLK (CLK), .RST (
                            RST), .Start (Start), .Instr (Instr), .LoopingAndResultNotReady (
                            nx3274), .Filter ({FilterDin_2__2__7,
                            FilterDin_2__2__6,FilterDin_2__2__5,
                            FilterDin_2__2__4,FilterDin_2__2__3,
                            FilterDin_2__2__2,FilterDin_2__2__1,
                            FilterDin_2__2__0}), .Window ({WindowDin_2__2__7,
                            WindowDin_2__2__6,WindowDin_2__2__5,
                            WindowDin_2__2__4,WindowDin_2__2__3,
                            WindowDin_2__2__2,WindowDin_2__2__1,
                            WindowDin_2__2__0}), .AdderBoothResult ({
                            L1FirstOperands_12__16,
                            L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_15,
                            L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_14,
                            L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_13,
                            L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_12,
                            L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_11,
                            L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_10,
                            L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_9,
                            L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_8,
                            L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_7,
                            L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_6,
                            L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_5,
                            L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_4,
                            L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_3,
                            L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_2,
                            L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_1,
                            L1_2_L2_2_G1_MINI_ALU_AdderBoothResult_0}), .BoothXORCheck (
                            L1_2_L2_2_G1_MINI_ALU_BoothXORCheck), .BoothResult (
                            {\$dummy [438],\$dummy [439],\$dummy [440],
                            \$dummy [441],\$dummy [442],\$dummy [443],
                            \$dummy [444],\$dummy [445]}), .BoothAddingOperand (
                            {L1_2_L2_2_G1_MINI_ALU_BoothOperand_16,
                            L1_2_L2_2_G1_MINI_ALU_BoothOperand_15,
                            L1_2_L2_2_G1_MINI_ALU_BoothOperand_14,
                            L1_2_L2_2_G1_MINI_ALU_BoothOperand_13,
                            L1_2_L2_2_G1_MINI_ALU_BoothOperand_12,
                            L1_2_L2_2_G1_MINI_ALU_BoothOperand_11,
                            L1_2_L2_2_G1_MINI_ALU_BoothOperand_10,
                            L1_2_L2_2_G1_MINI_ALU_BoothOperand_9,\$dummy [446],
                            \$dummy [447],\$dummy [448],\$dummy [449],
                            \$dummy [450],\$dummy [451],\$dummy [452],
                            \$dummy [453],\$dummy [454]}), .BoothP ({
                            L1_2_L2_2_G1_MINI_ALU_BoothP_16,
                            L1_2_L2_2_G1_MINI_ALU_BoothP_15,
                            L1_2_L2_2_G1_MINI_ALU_BoothP_14,
                            L1_2_L2_2_G1_MINI_ALU_BoothP_13,
                            L1_2_L2_2_G1_MINI_ALU_BoothP_12,
                            L1_2_L2_2_G1_MINI_ALU_BoothP_11,
                            L1_2_L2_2_G1_MINI_ALU_BoothP_10,
                            L1_2_L2_2_G1_MINI_ALU_BoothP_9,
                            L1_2_L2_2_G1_MINI_ALU_BoothP_8,
                            L1_2_L2_2_G1_MINI_ALU_BoothP_7,
                            L1_2_L2_2_G1_MINI_ALU_BoothP_6,
                            L1_2_L2_2_G1_MINI_ALU_BoothP_5,
                            L1_2_L2_2_G1_MINI_ALU_BoothP_4,
                            L1_2_L2_2_G1_MINI_ALU_BoothP_3,
                            L1_2_L2_2_G1_MINI_ALU_BoothP_2,
                            L1_2_L2_2_G1_MINI_ALU_BoothP_1,\$dummy [455]}), .LargeWindowShifted (
                            {\$dummy [456],\$dummy [457],\$dummy [458],
                            \$dummy [459],\$dummy [460],\$dummy [461],
                            \$dummy [462],\$dummy [463],\$dummy [464],
                            \$dummy [465],\$dummy [466],\$dummy [467],
                            \$dummy [468],\$dummy [469],\$dummy [470],
                            \$dummy [471],\$dummy [472]})) ;
    booth_adder_17_unfolded16 L1_2_L2_3_G2_MINI_ALU_BOOTH_ADDER (.AdderFirstOperand (
                              {L1ResultsLarge_0__16,L1ResultsLarge_0__15,
                              L1ResultsLarge_0__14,L1ResultsLarge_0__13,
                              L1ResultsLarge_0__12,L1ResultsLarge_0__11,
                              L1ResultsLarge_0__10,L1ResultsLarge_0__9,
                              L1ResultsLarge_0__8,L1ResultsLarge_0__7,
                              L1ResultsLarge_0__6,L1ResultsLarge_0__5,
                              L1ResultsLarge_0__4,L1ResultsLarge_0__3,
                              L1ResultsLarge_0__2,L1ResultsLarge_0__1,
                              L1ResultsLarge_0__0}), .AdderSecondOperand ({
                              L1ResultsLarge_1__16,L1ResultsLarge_1__15,
                              L1ResultsLarge_1__14,L1ResultsLarge_1__13,
                              L1ResultsLarge_1__12,L1ResultsLarge_1__11,
                              L1ResultsLarge_1__10,L1ResultsLarge_1__9,
                              L1ResultsLarge_1__8,L1ResultsLarge_1__7,
                              L1ResultsLarge_1__6,L1ResultsLarge_1__5,
                              L1ResultsLarge_1__4,L1ResultsLarge_1__3,
                              L1ResultsLarge_1__2,L1ResultsLarge_1__1,
                              L1ResultsLarge_1__0}), .BoothOperand ({
                              L1_2_L2_3_G2_MINI_ALU_BoothOperand_16,
                              L1_2_L2_3_G2_MINI_ALU_BoothOperand_15,
                              L1_2_L2_3_G2_MINI_ALU_BoothOperand_14,
                              L1_2_L2_3_G2_MINI_ALU_BoothOperand_13,
                              L1_2_L2_3_G2_MINI_ALU_BoothOperand_12,
                              L1_2_L2_3_G2_MINI_ALU_BoothOperand_11,
                              L1_2_L2_3_G2_MINI_ALU_BoothOperand_10,
                              L1_2_L2_3_G2_MINI_ALU_BoothOperand_9,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16}), .BoothP ({
                              L1_2_L2_3_G2_MINI_ALU_BoothP_16,
                              L1_2_L2_3_G2_MINI_ALU_BoothP_15,
                              L1_2_L2_3_G2_MINI_ALU_BoothP_14,
                              L1_2_L2_3_G2_MINI_ALU_BoothP_13,
                              L1_2_L2_3_G2_MINI_ALU_BoothP_12,
                              L1_2_L2_3_G2_MINI_ALU_BoothP_11,
                              L1_2_L2_3_G2_MINI_ALU_BoothP_10,
                              L1_2_L2_3_G2_MINI_ALU_BoothP_9,
                              L1_2_L2_3_G2_MINI_ALU_BoothP_8,
                              L1_2_L2_3_G2_MINI_ALU_BoothP_7,
                              L1_2_L2_3_G2_MINI_ALU_BoothP_6,
                              L1_2_L2_3_G2_MINI_ALU_BoothP_5,
                              L1_2_L2_3_G2_MINI_ALU_BoothP_4,
                              L1_2_L2_3_G2_MINI_ALU_BoothP_3,
                              L1_2_L2_3_G2_MINI_ALU_BoothP_2,
                              L1_2_L2_3_G2_MINI_ALU_BoothP_1,
                              L1_2_L2_3_G2_MINI_ALU_BoothP_0}), .SelOperand (
                              nx3284), .Operation (
                              L1_2_L2_3_G2_MINI_ALU_BoothXORCheck), .AdderResult (
                              {L2ResultsLarge_0__16,L2ResultsLarge_0__15,
                              L2ResultsLarge_0__14,L2ResultsLarge_0__13,
                              L2ResultsLarge_0__12,L2ResultsLarge_0__11,
                              L2ResultsLarge_0__10,L2ResultsLarge_0__9,
                              L2ResultsLarge_0__8,L2ResultsLarge_0__7,
                              L2ResultsLarge_0__6,L2ResultsLarge_0__5,
                              L2ResultsLarge_0__4,L2ResultsLarge_0__3,
                              L2ResultsLarge_0__2,L2ResultsLarge_0__1,
                              L2ResultsLarge_0__0}), .AdderBoothResult ({
                              \$dummy [473],
                              L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_15,
                              L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_14,
                              L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_13,
                              L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_12,
                              L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_11,
                              L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_10,
                              L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_9,
                              L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_8,
                              L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_7,
                              L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_6,
                              L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_5,
                              L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_4,
                              L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_3,
                              L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_2,
                              L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_1,
                              L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_0})) ;
    booth_unit_17 L1_2_L2_3_G2_MINI_ALU_BOOTH_UNIT (.CLK (CLK), .RST (RST), .Start (
                  Start), .Instr (Instr), .LoopingAndResultNotReady (nx3274), .Filter (
                  {FilterDin_2__3__7,FilterDin_2__3__6,FilterDin_2__3__5,
                  FilterDin_2__3__4,FilterDin_2__3__3,FilterDin_2__3__2,
                  FilterDin_2__3__1,FilterDin_2__3__0}), .Window ({
                  WindowDin_2__3__7,WindowDin_2__3__6,WindowDin_2__3__5,
                  WindowDin_2__3__4,WindowDin_2__3__3,WindowDin_2__3__2,
                  WindowDin_2__3__1,WindowDin_2__3__0}), .AdderBoothResult ({
                  L1FirstOperands_12__16,
                  L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_15,
                  L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_14,
                  L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_13,
                  L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_12,
                  L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_11,
                  L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_10,
                  L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_9,
                  L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_8,
                  L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_7,
                  L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_6,
                  L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_5,
                  L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_4,
                  L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_3,
                  L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_2,
                  L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_1,
                  L1_2_L2_3_G2_MINI_ALU_AdderBoothResult_0}), .BoothXORCheck (
                  L1_2_L2_3_G2_MINI_ALU_BoothXORCheck), .BoothResult ({
                  \$dummy [474],\$dummy [475],\$dummy [476],\$dummy [477],
                  \$dummy [478],\$dummy [479],\$dummy [480],\$dummy [481]}), .BoothAddingOperand (
                  {L1_2_L2_3_G2_MINI_ALU_BoothOperand_16,
                  L1_2_L2_3_G2_MINI_ALU_BoothOperand_15,
                  L1_2_L2_3_G2_MINI_ALU_BoothOperand_14,
                  L1_2_L2_3_G2_MINI_ALU_BoothOperand_13,
                  L1_2_L2_3_G2_MINI_ALU_BoothOperand_12,
                  L1_2_L2_3_G2_MINI_ALU_BoothOperand_11,
                  L1_2_L2_3_G2_MINI_ALU_BoothOperand_10,
                  L1_2_L2_3_G2_MINI_ALU_BoothOperand_9,\$dummy [482],
                  \$dummy [483],\$dummy [484],\$dummy [485],\$dummy [486],
                  \$dummy [487],\$dummy [488],\$dummy [489],\$dummy [490]}), .BoothP (
                  {L1_2_L2_3_G2_MINI_ALU_BoothP_16,
                  L1_2_L2_3_G2_MINI_ALU_BoothP_15,
                  L1_2_L2_3_G2_MINI_ALU_BoothP_14,
                  L1_2_L2_3_G2_MINI_ALU_BoothP_13,
                  L1_2_L2_3_G2_MINI_ALU_BoothP_12,
                  L1_2_L2_3_G2_MINI_ALU_BoothP_11,
                  L1_2_L2_3_G2_MINI_ALU_BoothP_10,L1_2_L2_3_G2_MINI_ALU_BoothP_9
                  ,L1_2_L2_3_G2_MINI_ALU_BoothP_8,L1_2_L2_3_G2_MINI_ALU_BoothP_7
                  ,L1_2_L2_3_G2_MINI_ALU_BoothP_6,L1_2_L2_3_G2_MINI_ALU_BoothP_5
                  ,L1_2_L2_3_G2_MINI_ALU_BoothP_4,L1_2_L2_3_G2_MINI_ALU_BoothP_3
                  ,L1_2_L2_3_G2_MINI_ALU_BoothP_2,L1_2_L2_3_G2_MINI_ALU_BoothP_1
                  ,L1_2_L2_3_G2_MINI_ALU_BoothP_0}), .LargeWindowShifted ({
                  \$dummy [491],\$dummy [492],\$dummy [493],\$dummy [494],
                  \$dummy [495],\$dummy [496],\$dummy [497],\$dummy [498],
                  \$dummy [499],\$dummy [500],\$dummy [501],\$dummy [502],
                  \$dummy [503],\$dummy [504],\$dummy [505],\$dummy [506],
                  \$dummy [507]})) ;
    booth_adder_17_unfolded16 L1_2_L2_4_G2_MINI_ALU_BOOTH_ADDER (.AdderFirstOperand (
                              {L1ResultsLarge_2__16,L1ResultsLarge_2__15,
                              L1ResultsLarge_2__14,L1ResultsLarge_2__13,
                              L1ResultsLarge_2__12,L1ResultsLarge_2__11,
                              L1ResultsLarge_2__10,L1ResultsLarge_2__9,
                              L1ResultsLarge_2__8,L1ResultsLarge_2__7,
                              L1ResultsLarge_2__6,L1ResultsLarge_2__5,
                              L1ResultsLarge_2__4,L1ResultsLarge_2__3,
                              L1ResultsLarge_2__2,L1ResultsLarge_2__1,
                              L1ResultsLarge_2__0}), .AdderSecondOperand ({
                              L1ResultsLarge_3__16,L1ResultsLarge_3__15,
                              L1ResultsLarge_3__14,L1ResultsLarge_3__13,
                              L1ResultsLarge_3__12,L1ResultsLarge_3__11,
                              L1ResultsLarge_3__10,L1ResultsLarge_3__9,
                              L1ResultsLarge_3__8,L1ResultsLarge_3__7,
                              L1ResultsLarge_3__6,L1ResultsLarge_3__5,
                              L1ResultsLarge_3__4,L1ResultsLarge_3__3,
                              L1ResultsLarge_3__2,L1ResultsLarge_3__1,
                              L1ResultsLarge_3__0}), .BoothOperand ({
                              L1_2_L2_4_G2_MINI_ALU_BoothOperand_16,
                              L1_2_L2_4_G2_MINI_ALU_BoothOperand_15,
                              L1_2_L2_4_G2_MINI_ALU_BoothOperand_14,
                              L1_2_L2_4_G2_MINI_ALU_BoothOperand_13,
                              L1_2_L2_4_G2_MINI_ALU_BoothOperand_12,
                              L1_2_L2_4_G2_MINI_ALU_BoothOperand_11,
                              L1_2_L2_4_G2_MINI_ALU_BoothOperand_10,
                              L1_2_L2_4_G2_MINI_ALU_BoothOperand_9,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16}), .BoothP ({
                              L1_2_L2_4_G2_MINI_ALU_BoothP_16,
                              L1_2_L2_4_G2_MINI_ALU_BoothP_15,
                              L1_2_L2_4_G2_MINI_ALU_BoothP_14,
                              L1_2_L2_4_G2_MINI_ALU_BoothP_13,
                              L1_2_L2_4_G2_MINI_ALU_BoothP_12,
                              L1_2_L2_4_G2_MINI_ALU_BoothP_11,
                              L1_2_L2_4_G2_MINI_ALU_BoothP_10,
                              L1_2_L2_4_G2_MINI_ALU_BoothP_9,
                              L1_2_L2_4_G2_MINI_ALU_BoothP_8,
                              L1_2_L2_4_G2_MINI_ALU_BoothP_7,
                              L1_2_L2_4_G2_MINI_ALU_BoothP_6,
                              L1_2_L2_4_G2_MINI_ALU_BoothP_5,
                              L1_2_L2_4_G2_MINI_ALU_BoothP_4,
                              L1_2_L2_4_G2_MINI_ALU_BoothP_3,
                              L1_2_L2_4_G2_MINI_ALU_BoothP_2,
                              L1_2_L2_4_G2_MINI_ALU_BoothP_1,
                              L1_2_L2_4_G2_MINI_ALU_BoothP_0}), .SelOperand (
                              nx3284), .Operation (
                              L1_2_L2_4_G2_MINI_ALU_BoothXORCheck), .AdderResult (
                              {L2ResultsLarge_1__16,L2ResultsLarge_1__15,
                              L2ResultsLarge_1__14,L2ResultsLarge_1__13,
                              L2ResultsLarge_1__12,L2ResultsLarge_1__11,
                              L2ResultsLarge_1__10,L2ResultsLarge_1__9,
                              L2ResultsLarge_1__8,L2ResultsLarge_1__7,
                              L2ResultsLarge_1__6,L2ResultsLarge_1__5,
                              L2ResultsLarge_1__4,L2ResultsLarge_1__3,
                              L2ResultsLarge_1__2,L2ResultsLarge_1__1,
                              L2ResultsLarge_1__0}), .AdderBoothResult ({
                              \$dummy [508],
                              L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_15,
                              L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_14,
                              L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_13,
                              L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_12,
                              L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_11,
                              L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_10,
                              L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_9,
                              L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_8,
                              L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_7,
                              L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_6,
                              L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_5,
                              L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_4,
                              L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_3,
                              L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_2,
                              L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_1,
                              L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_0})) ;
    booth_unit_17 L1_2_L2_4_G2_MINI_ALU_BOOTH_UNIT (.CLK (CLK), .RST (RST), .Start (
                  Start), .Instr (Instr), .LoopingAndResultNotReady (nx3276), .Filter (
                  {FilterDin_2__4__7,FilterDin_2__4__6,FilterDin_2__4__5,
                  FilterDin_2__4__4,FilterDin_2__4__3,FilterDin_2__4__2,
                  FilterDin_2__4__1,FilterDin_2__4__0}), .Window ({
                  WindowDin_2__4__7,WindowDin_2__4__6,WindowDin_2__4__5,
                  WindowDin_2__4__4,WindowDin_2__4__3,WindowDin_2__4__2,
                  WindowDin_2__4__1,WindowDin_2__4__0}), .AdderBoothResult ({
                  L1FirstOperands_12__16,
                  L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_15,
                  L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_14,
                  L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_13,
                  L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_12,
                  L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_11,
                  L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_10,
                  L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_9,
                  L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_8,
                  L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_7,
                  L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_6,
                  L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_5,
                  L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_4,
                  L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_3,
                  L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_2,
                  L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_1,
                  L1_2_L2_4_G2_MINI_ALU_AdderBoothResult_0}), .BoothXORCheck (
                  L1_2_L2_4_G2_MINI_ALU_BoothXORCheck), .BoothResult ({
                  \$dummy [509],\$dummy [510],\$dummy [511],\$dummy [512],
                  \$dummy [513],\$dummy [514],\$dummy [515],\$dummy [516]}), .BoothAddingOperand (
                  {L1_2_L2_4_G2_MINI_ALU_BoothOperand_16,
                  L1_2_L2_4_G2_MINI_ALU_BoothOperand_15,
                  L1_2_L2_4_G2_MINI_ALU_BoothOperand_14,
                  L1_2_L2_4_G2_MINI_ALU_BoothOperand_13,
                  L1_2_L2_4_G2_MINI_ALU_BoothOperand_12,
                  L1_2_L2_4_G2_MINI_ALU_BoothOperand_11,
                  L1_2_L2_4_G2_MINI_ALU_BoothOperand_10,
                  L1_2_L2_4_G2_MINI_ALU_BoothOperand_9,\$dummy [517],
                  \$dummy [518],\$dummy [519],\$dummy [520],\$dummy [521],
                  \$dummy [522],\$dummy [523],\$dummy [524],\$dummy [525]}), .BoothP (
                  {L1_2_L2_4_G2_MINI_ALU_BoothP_16,
                  L1_2_L2_4_G2_MINI_ALU_BoothP_15,
                  L1_2_L2_4_G2_MINI_ALU_BoothP_14,
                  L1_2_L2_4_G2_MINI_ALU_BoothP_13,
                  L1_2_L2_4_G2_MINI_ALU_BoothP_12,
                  L1_2_L2_4_G2_MINI_ALU_BoothP_11,
                  L1_2_L2_4_G2_MINI_ALU_BoothP_10,L1_2_L2_4_G2_MINI_ALU_BoothP_9
                  ,L1_2_L2_4_G2_MINI_ALU_BoothP_8,L1_2_L2_4_G2_MINI_ALU_BoothP_7
                  ,L1_2_L2_4_G2_MINI_ALU_BoothP_6,L1_2_L2_4_G2_MINI_ALU_BoothP_5
                  ,L1_2_L2_4_G2_MINI_ALU_BoothP_4,L1_2_L2_4_G2_MINI_ALU_BoothP_3
                  ,L1_2_L2_4_G2_MINI_ALU_BoothP_2,L1_2_L2_4_G2_MINI_ALU_BoothP_1
                  ,L1_2_L2_4_G2_MINI_ALU_BoothP_0}), .LargeWindowShifted ({
                  \$dummy [526],\$dummy [527],\$dummy [528],\$dummy [529],
                  \$dummy [530],\$dummy [531],\$dummy [532],\$dummy [533],
                  \$dummy [534],\$dummy [535],\$dummy [536],\$dummy [537],
                  \$dummy [538],\$dummy [539],\$dummy [540],\$dummy [541],
                  \$dummy [542]})) ;
    booth_adder_17_unfolded16 L1_3_L2_0_G2_MINI_ALU_BOOTH_ADDER (.AdderFirstOperand (
                              {L1ResultsLarge_4__16,L1ResultsLarge_4__15,
                              L1ResultsLarge_4__14,L1ResultsLarge_4__13,
                              L1ResultsLarge_4__12,L1ResultsLarge_4__11,
                              L1ResultsLarge_4__10,L1ResultsLarge_4__9,
                              L1ResultsLarge_4__8,L1ResultsLarge_4__7,
                              L1ResultsLarge_4__6,L1ResultsLarge_4__5,
                              L1ResultsLarge_4__4,L1ResultsLarge_4__3,
                              L1ResultsLarge_4__2,L1ResultsLarge_4__1,
                              L1ResultsLarge_4__0}), .AdderSecondOperand ({
                              L1ResultsLarge_5__16,L1ResultsLarge_5__15,
                              L1ResultsLarge_5__14,L1ResultsLarge_5__13,
                              L1ResultsLarge_5__12,L1ResultsLarge_5__11,
                              L1ResultsLarge_5__10,L1ResultsLarge_5__9,
                              L1ResultsLarge_5__8,L1ResultsLarge_5__7,
                              L1ResultsLarge_5__6,L1ResultsLarge_5__5,
                              L1ResultsLarge_5__4,L1ResultsLarge_5__3,
                              L1ResultsLarge_5__2,L1ResultsLarge_5__1,
                              L1ResultsLarge_5__0}), .BoothOperand ({
                              L1_3_L2_0_G2_MINI_ALU_BoothOperand_16,
                              L1_3_L2_0_G2_MINI_ALU_BoothOperand_15,
                              L1_3_L2_0_G2_MINI_ALU_BoothOperand_14,
                              L1_3_L2_0_G2_MINI_ALU_BoothOperand_13,
                              L1_3_L2_0_G2_MINI_ALU_BoothOperand_12,
                              L1_3_L2_0_G2_MINI_ALU_BoothOperand_11,
                              L1_3_L2_0_G2_MINI_ALU_BoothOperand_10,
                              L1_3_L2_0_G2_MINI_ALU_BoothOperand_9,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16}), .BoothP ({
                              L1_3_L2_0_G2_MINI_ALU_BoothP_16,
                              L1_3_L2_0_G2_MINI_ALU_BoothP_15,
                              L1_3_L2_0_G2_MINI_ALU_BoothP_14,
                              L1_3_L2_0_G2_MINI_ALU_BoothP_13,
                              L1_3_L2_0_G2_MINI_ALU_BoothP_12,
                              L1_3_L2_0_G2_MINI_ALU_BoothP_11,
                              L1_3_L2_0_G2_MINI_ALU_BoothP_10,
                              L1_3_L2_0_G2_MINI_ALU_BoothP_9,
                              L1_3_L2_0_G2_MINI_ALU_BoothP_8,
                              L1_3_L2_0_G2_MINI_ALU_BoothP_7,
                              L1_3_L2_0_G2_MINI_ALU_BoothP_6,
                              L1_3_L2_0_G2_MINI_ALU_BoothP_5,
                              L1_3_L2_0_G2_MINI_ALU_BoothP_4,
                              L1_3_L2_0_G2_MINI_ALU_BoothP_3,
                              L1_3_L2_0_G2_MINI_ALU_BoothP_2,
                              L1_3_L2_0_G2_MINI_ALU_BoothP_1,
                              L1_3_L2_0_G2_MINI_ALU_BoothP_0}), .SelOperand (
                              nx3284), .Operation (
                              L1_3_L2_0_G2_MINI_ALU_BoothXORCheck), .AdderResult (
                              {L2ResultsLarge_2__16,L2ResultsLarge_2__15,
                              L2ResultsLarge_2__14,L2ResultsLarge_2__13,
                              L2ResultsLarge_2__12,L2ResultsLarge_2__11,
                              L2ResultsLarge_2__10,L2ResultsLarge_2__9,
                              L2ResultsLarge_2__8,L2ResultsLarge_2__7,
                              L2ResultsLarge_2__6,L2ResultsLarge_2__5,
                              L2ResultsLarge_2__4,L2ResultsLarge_2__3,
                              L2ResultsLarge_2__2,L2ResultsLarge_2__1,
                              L2ResultsLarge_2__0}), .AdderBoothResult ({
                              \$dummy [543],
                              L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_15,
                              L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_14,
                              L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_13,
                              L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_12,
                              L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_11,
                              L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_10,
                              L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_9,
                              L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_8,
                              L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_7,
                              L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_6,
                              L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_5,
                              L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_4,
                              L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_3,
                              L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_2,
                              L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_1,
                              L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_0})) ;
    booth_unit_17 L1_3_L2_0_G2_MINI_ALU_BOOTH_UNIT (.CLK (CLK), .RST (RST), .Start (
                  Start), .Instr (Instr), .LoopingAndResultNotReady (nx3276), .Filter (
                  {FilterDin_3__0__7,FilterDin_3__0__6,FilterDin_3__0__5,
                  FilterDin_3__0__4,FilterDin_3__0__3,FilterDin_3__0__2,
                  FilterDin_3__0__1,FilterDin_3__0__0}), .Window ({
                  WindowDin_3__0__7,WindowDin_3__0__6,WindowDin_3__0__5,
                  WindowDin_3__0__4,WindowDin_3__0__3,WindowDin_3__0__2,
                  WindowDin_3__0__1,WindowDin_3__0__0}), .AdderBoothResult ({
                  L1FirstOperands_12__16,
                  L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_15,
                  L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_14,
                  L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_13,
                  L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_12,
                  L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_11,
                  L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_10,
                  L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_9,
                  L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_8,
                  L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_7,
                  L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_6,
                  L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_5,
                  L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_4,
                  L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_3,
                  L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_2,
                  L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_1,
                  L1_3_L2_0_G2_MINI_ALU_AdderBoothResult_0}), .BoothXORCheck (
                  L1_3_L2_0_G2_MINI_ALU_BoothXORCheck), .BoothResult ({
                  \$dummy [544],\$dummy [545],\$dummy [546],\$dummy [547],
                  \$dummy [548],\$dummy [549],\$dummy [550],\$dummy [551]}), .BoothAddingOperand (
                  {L1_3_L2_0_G2_MINI_ALU_BoothOperand_16,
                  L1_3_L2_0_G2_MINI_ALU_BoothOperand_15,
                  L1_3_L2_0_G2_MINI_ALU_BoothOperand_14,
                  L1_3_L2_0_G2_MINI_ALU_BoothOperand_13,
                  L1_3_L2_0_G2_MINI_ALU_BoothOperand_12,
                  L1_3_L2_0_G2_MINI_ALU_BoothOperand_11,
                  L1_3_L2_0_G2_MINI_ALU_BoothOperand_10,
                  L1_3_L2_0_G2_MINI_ALU_BoothOperand_9,\$dummy [552],
                  \$dummy [553],\$dummy [554],\$dummy [555],\$dummy [556],
                  \$dummy [557],\$dummy [558],\$dummy [559],\$dummy [560]}), .BoothP (
                  {L1_3_L2_0_G2_MINI_ALU_BoothP_16,
                  L1_3_L2_0_G2_MINI_ALU_BoothP_15,
                  L1_3_L2_0_G2_MINI_ALU_BoothP_14,
                  L1_3_L2_0_G2_MINI_ALU_BoothP_13,
                  L1_3_L2_0_G2_MINI_ALU_BoothP_12,
                  L1_3_L2_0_G2_MINI_ALU_BoothP_11,
                  L1_3_L2_0_G2_MINI_ALU_BoothP_10,L1_3_L2_0_G2_MINI_ALU_BoothP_9
                  ,L1_3_L2_0_G2_MINI_ALU_BoothP_8,L1_3_L2_0_G2_MINI_ALU_BoothP_7
                  ,L1_3_L2_0_G2_MINI_ALU_BoothP_6,L1_3_L2_0_G2_MINI_ALU_BoothP_5
                  ,L1_3_L2_0_G2_MINI_ALU_BoothP_4,L1_3_L2_0_G2_MINI_ALU_BoothP_3
                  ,L1_3_L2_0_G2_MINI_ALU_BoothP_2,L1_3_L2_0_G2_MINI_ALU_BoothP_1
                  ,L1_3_L2_0_G2_MINI_ALU_BoothP_0}), .LargeWindowShifted ({
                  \$dummy [561],\$dummy [562],\$dummy [563],\$dummy [564],
                  \$dummy [565],\$dummy [566],\$dummy [567],\$dummy [568],
                  \$dummy [569],\$dummy [570],\$dummy [571],\$dummy [572],
                  \$dummy [573],\$dummy [574],\$dummy [575],\$dummy [576],
                  \$dummy [577]})) ;
    booth_adder_17_unfolded16 L1_3_L2_1_G2_MINI_ALU_BOOTH_ADDER (.AdderFirstOperand (
                              {L1ResultsLarge_6__16,L1ResultsLarge_6__15,
                              L1ResultsLarge_6__14,L1ResultsLarge_6__13,
                              L1ResultsLarge_6__12,L1ResultsLarge_6__11,
                              L1ResultsLarge_6__10,L1ResultsLarge_6__9,
                              L1ResultsLarge_6__8,L1ResultsLarge_6__7,
                              L1ResultsLarge_6__6,L1ResultsLarge_6__5,
                              L1ResultsLarge_6__4,L1ResultsLarge_6__3,
                              L1ResultsLarge_6__2,L1ResultsLarge_6__1,
                              L1ResultsLarge_6__0}), .AdderSecondOperand ({
                              L1ResultsLarge_7__16,L1ResultsLarge_7__15,
                              L1ResultsLarge_7__14,L1ResultsLarge_7__13,
                              L1ResultsLarge_7__12,L1ResultsLarge_7__11,
                              L1ResultsLarge_7__10,L1ResultsLarge_7__9,
                              L1ResultsLarge_7__8,L1ResultsLarge_7__7,
                              L1ResultsLarge_7__6,L1ResultsLarge_7__5,
                              L1ResultsLarge_7__4,L1ResultsLarge_7__3,
                              L1ResultsLarge_7__2,L1ResultsLarge_7__1,
                              L1ResultsLarge_7__0}), .BoothOperand ({
                              L1_3_L2_1_G2_MINI_ALU_BoothOperand_16,
                              L1_3_L2_1_G2_MINI_ALU_BoothOperand_15,
                              L1_3_L2_1_G2_MINI_ALU_BoothOperand_14,
                              L1_3_L2_1_G2_MINI_ALU_BoothOperand_13,
                              L1_3_L2_1_G2_MINI_ALU_BoothOperand_12,
                              L1_3_L2_1_G2_MINI_ALU_BoothOperand_11,
                              L1_3_L2_1_G2_MINI_ALU_BoothOperand_10,
                              L1_3_L2_1_G2_MINI_ALU_BoothOperand_9,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16}), .BoothP ({
                              L1_3_L2_1_G2_MINI_ALU_BoothP_16,
                              L1_3_L2_1_G2_MINI_ALU_BoothP_15,
                              L1_3_L2_1_G2_MINI_ALU_BoothP_14,
                              L1_3_L2_1_G2_MINI_ALU_BoothP_13,
                              L1_3_L2_1_G2_MINI_ALU_BoothP_12,
                              L1_3_L2_1_G2_MINI_ALU_BoothP_11,
                              L1_3_L2_1_G2_MINI_ALU_BoothP_10,
                              L1_3_L2_1_G2_MINI_ALU_BoothP_9,
                              L1_3_L2_1_G2_MINI_ALU_BoothP_8,
                              L1_3_L2_1_G2_MINI_ALU_BoothP_7,
                              L1_3_L2_1_G2_MINI_ALU_BoothP_6,
                              L1_3_L2_1_G2_MINI_ALU_BoothP_5,
                              L1_3_L2_1_G2_MINI_ALU_BoothP_4,
                              L1_3_L2_1_G2_MINI_ALU_BoothP_3,
                              L1_3_L2_1_G2_MINI_ALU_BoothP_2,
                              L1_3_L2_1_G2_MINI_ALU_BoothP_1,
                              L1_3_L2_1_G2_MINI_ALU_BoothP_0}), .SelOperand (
                              nx3282), .Operation (
                              L1_3_L2_1_G2_MINI_ALU_BoothXORCheck), .AdderResult (
                              {L2ResultsLarge_3__16,L2ResultsLarge_3__15,
                              L2ResultsLarge_3__14,L2ResultsLarge_3__13,
                              L2ResultsLarge_3__12,L2ResultsLarge_3__11,
                              L2ResultsLarge_3__10,L2ResultsLarge_3__9,
                              L2ResultsLarge_3__8,L2ResultsLarge_3__7,
                              L2ResultsLarge_3__6,L2ResultsLarge_3__5,
                              L2ResultsLarge_3__4,L2ResultsLarge_3__3,
                              L2ResultsLarge_3__2,L2ResultsLarge_3__1,
                              L2ResultsLarge_3__0}), .AdderBoothResult ({
                              \$dummy [578],
                              L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_15,
                              L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_14,
                              L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_13,
                              L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_12,
                              L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_11,
                              L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_10,
                              L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_9,
                              L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_8,
                              L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_7,
                              L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_6,
                              L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_5,
                              L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_4,
                              L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_3,
                              L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_2,
                              L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_1,
                              L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_0})) ;
    booth_unit_17 L1_3_L2_1_G2_MINI_ALU_BOOTH_UNIT (.CLK (CLK), .RST (RST), .Start (
                  Start), .Instr (Instr), .LoopingAndResultNotReady (nx3276), .Filter (
                  {FilterDin_3__1__7,FilterDin_3__1__6,FilterDin_3__1__5,
                  FilterDin_3__1__4,FilterDin_3__1__3,FilterDin_3__1__2,
                  FilterDin_3__1__1,FilterDin_3__1__0}), .Window ({
                  WindowDin_3__1__7,WindowDin_3__1__6,WindowDin_3__1__5,
                  WindowDin_3__1__4,WindowDin_3__1__3,WindowDin_3__1__2,
                  WindowDin_3__1__1,WindowDin_3__1__0}), .AdderBoothResult ({
                  L1FirstOperands_12__16,
                  L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_15,
                  L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_14,
                  L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_13,
                  L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_12,
                  L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_11,
                  L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_10,
                  L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_9,
                  L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_8,
                  L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_7,
                  L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_6,
                  L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_5,
                  L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_4,
                  L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_3,
                  L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_2,
                  L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_1,
                  L1_3_L2_1_G2_MINI_ALU_AdderBoothResult_0}), .BoothXORCheck (
                  L1_3_L2_1_G2_MINI_ALU_BoothXORCheck), .BoothResult ({
                  \$dummy [579],\$dummy [580],\$dummy [581],\$dummy [582],
                  \$dummy [583],\$dummy [584],\$dummy [585],\$dummy [586]}), .BoothAddingOperand (
                  {L1_3_L2_1_G2_MINI_ALU_BoothOperand_16,
                  L1_3_L2_1_G2_MINI_ALU_BoothOperand_15,
                  L1_3_L2_1_G2_MINI_ALU_BoothOperand_14,
                  L1_3_L2_1_G2_MINI_ALU_BoothOperand_13,
                  L1_3_L2_1_G2_MINI_ALU_BoothOperand_12,
                  L1_3_L2_1_G2_MINI_ALU_BoothOperand_11,
                  L1_3_L2_1_G2_MINI_ALU_BoothOperand_10,
                  L1_3_L2_1_G2_MINI_ALU_BoothOperand_9,\$dummy [587],
                  \$dummy [588],\$dummy [589],\$dummy [590],\$dummy [591],
                  \$dummy [592],\$dummy [593],\$dummy [594],\$dummy [595]}), .BoothP (
                  {L1_3_L2_1_G2_MINI_ALU_BoothP_16,
                  L1_3_L2_1_G2_MINI_ALU_BoothP_15,
                  L1_3_L2_1_G2_MINI_ALU_BoothP_14,
                  L1_3_L2_1_G2_MINI_ALU_BoothP_13,
                  L1_3_L2_1_G2_MINI_ALU_BoothP_12,
                  L1_3_L2_1_G2_MINI_ALU_BoothP_11,
                  L1_3_L2_1_G2_MINI_ALU_BoothP_10,L1_3_L2_1_G2_MINI_ALU_BoothP_9
                  ,L1_3_L2_1_G2_MINI_ALU_BoothP_8,L1_3_L2_1_G2_MINI_ALU_BoothP_7
                  ,L1_3_L2_1_G2_MINI_ALU_BoothP_6,L1_3_L2_1_G2_MINI_ALU_BoothP_5
                  ,L1_3_L2_1_G2_MINI_ALU_BoothP_4,L1_3_L2_1_G2_MINI_ALU_BoothP_3
                  ,L1_3_L2_1_G2_MINI_ALU_BoothP_2,L1_3_L2_1_G2_MINI_ALU_BoothP_1
                  ,L1_3_L2_1_G2_MINI_ALU_BoothP_0}), .LargeWindowShifted ({
                  \$dummy [596],\$dummy [597],\$dummy [598],\$dummy [599],
                  \$dummy [600],\$dummy [601],\$dummy [602],\$dummy [603],
                  \$dummy [604],\$dummy [605],\$dummy [606],\$dummy [607],
                  \$dummy [608],\$dummy [609],\$dummy [610],\$dummy [611],
                  \$dummy [612]})) ;
    booth_adder_17_unfolded16 L1_3_L2_2_G2_MINI_ALU_BOOTH_ADDER (.AdderFirstOperand (
                              {L1ResultsLarge_8__16,L1ResultsLarge_8__15,
                              L1ResultsLarge_8__14,L1ResultsLarge_8__13,
                              L1ResultsLarge_8__12,L1ResultsLarge_8__11,
                              L1ResultsLarge_8__10,L1ResultsLarge_8__9,
                              L1ResultsLarge_8__8,L1ResultsLarge_8__7,
                              L1ResultsLarge_8__6,L1ResultsLarge_8__5,
                              L1ResultsLarge_8__4,L1ResultsLarge_8__3,
                              L1ResultsLarge_8__2,L1ResultsLarge_8__1,
                              L1ResultsLarge_8__0}), .AdderSecondOperand ({
                              L1ResultsLarge_9__16,L1ResultsLarge_9__15,
                              L1ResultsLarge_9__14,L1ResultsLarge_9__13,
                              L1ResultsLarge_9__12,L1ResultsLarge_9__11,
                              L1ResultsLarge_9__10,L1ResultsLarge_9__9,
                              L1ResultsLarge_9__8,L1ResultsLarge_9__7,
                              L1ResultsLarge_9__6,L1ResultsLarge_9__5,
                              L1ResultsLarge_9__4,L1ResultsLarge_9__3,
                              L1ResultsLarge_9__2,L1ResultsLarge_9__1,
                              L1ResultsLarge_9__0}), .BoothOperand ({
                              L1_3_L2_2_G2_MINI_ALU_BoothOperand_16,
                              L1_3_L2_2_G2_MINI_ALU_BoothOperand_15,
                              L1_3_L2_2_G2_MINI_ALU_BoothOperand_14,
                              L1_3_L2_2_G2_MINI_ALU_BoothOperand_13,
                              L1_3_L2_2_G2_MINI_ALU_BoothOperand_12,
                              L1_3_L2_2_G2_MINI_ALU_BoothOperand_11,
                              L1_3_L2_2_G2_MINI_ALU_BoothOperand_10,
                              L1_3_L2_2_G2_MINI_ALU_BoothOperand_9,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16}), .BoothP ({
                              L1_3_L2_2_G2_MINI_ALU_BoothP_16,
                              L1_3_L2_2_G2_MINI_ALU_BoothP_15,
                              L1_3_L2_2_G2_MINI_ALU_BoothP_14,
                              L1_3_L2_2_G2_MINI_ALU_BoothP_13,
                              L1_3_L2_2_G2_MINI_ALU_BoothP_12,
                              L1_3_L2_2_G2_MINI_ALU_BoothP_11,
                              L1_3_L2_2_G2_MINI_ALU_BoothP_10,
                              L1_3_L2_2_G2_MINI_ALU_BoothP_9,
                              L1_3_L2_2_G2_MINI_ALU_BoothP_8,
                              L1_3_L2_2_G2_MINI_ALU_BoothP_7,
                              L1_3_L2_2_G2_MINI_ALU_BoothP_6,
                              L1_3_L2_2_G2_MINI_ALU_BoothP_5,
                              L1_3_L2_2_G2_MINI_ALU_BoothP_4,
                              L1_3_L2_2_G2_MINI_ALU_BoothP_3,
                              L1_3_L2_2_G2_MINI_ALU_BoothP_2,
                              L1_3_L2_2_G2_MINI_ALU_BoothP_1,
                              L1_3_L2_2_G2_MINI_ALU_BoothP_0}), .SelOperand (
                              nx3284), .Operation (
                              L1_3_L2_2_G2_MINI_ALU_BoothXORCheck), .AdderResult (
                              {L2ResultsLarge_4__16,L2ResultsLarge_4__15,
                              L2ResultsLarge_4__14,L2ResultsLarge_4__13,
                              L2ResultsLarge_4__12,L2ResultsLarge_4__11,
                              L2ResultsLarge_4__10,L2ResultsLarge_4__9,
                              L2ResultsLarge_4__8,L2ResultsLarge_4__7,
                              L2ResultsLarge_4__6,L2ResultsLarge_4__5,
                              L2ResultsLarge_4__4,L2ResultsLarge_4__3,
                              L2ResultsLarge_4__2,L2ResultsLarge_4__1,
                              L2ResultsLarge_4__0}), .AdderBoothResult ({
                              \$dummy [613],
                              L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_15,
                              L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_14,
                              L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_13,
                              L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_12,
                              L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_11,
                              L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_10,
                              L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_9,
                              L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_8,
                              L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_7,
                              L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_6,
                              L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_5,
                              L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_4,
                              L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_3,
                              L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_2,
                              L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_1,
                              L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_0})) ;
    booth_unit_17 L1_3_L2_2_G2_MINI_ALU_BOOTH_UNIT (.CLK (CLK), .RST (RST), .Start (
                  Start), .Instr (Instr), .LoopingAndResultNotReady (nx3276), .Filter (
                  {FilterDin_3__2__7,FilterDin_3__2__6,FilterDin_3__2__5,
                  FilterDin_3__2__4,FilterDin_3__2__3,FilterDin_3__2__2,
                  FilterDin_3__2__1,FilterDin_3__2__0}), .Window ({
                  WindowDin_3__2__7,WindowDin_3__2__6,WindowDin_3__2__5,
                  WindowDin_3__2__4,WindowDin_3__2__3,WindowDin_3__2__2,
                  WindowDin_3__2__1,WindowDin_3__2__0}), .AdderBoothResult ({
                  L1FirstOperands_12__16,
                  L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_15,
                  L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_14,
                  L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_13,
                  L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_12,
                  L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_11,
                  L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_10,
                  L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_9,
                  L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_8,
                  L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_7,
                  L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_6,
                  L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_5,
                  L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_4,
                  L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_3,
                  L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_2,
                  L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_1,
                  L1_3_L2_2_G2_MINI_ALU_AdderBoothResult_0}), .BoothXORCheck (
                  L1_3_L2_2_G2_MINI_ALU_BoothXORCheck), .BoothResult ({
                  \$dummy [614],\$dummy [615],\$dummy [616],\$dummy [617],
                  \$dummy [618],\$dummy [619],\$dummy [620],\$dummy [621]}), .BoothAddingOperand (
                  {L1_3_L2_2_G2_MINI_ALU_BoothOperand_16,
                  L1_3_L2_2_G2_MINI_ALU_BoothOperand_15,
                  L1_3_L2_2_G2_MINI_ALU_BoothOperand_14,
                  L1_3_L2_2_G2_MINI_ALU_BoothOperand_13,
                  L1_3_L2_2_G2_MINI_ALU_BoothOperand_12,
                  L1_3_L2_2_G2_MINI_ALU_BoothOperand_11,
                  L1_3_L2_2_G2_MINI_ALU_BoothOperand_10,
                  L1_3_L2_2_G2_MINI_ALU_BoothOperand_9,\$dummy [622],
                  \$dummy [623],\$dummy [624],\$dummy [625],\$dummy [626],
                  \$dummy [627],\$dummy [628],\$dummy [629],\$dummy [630]}), .BoothP (
                  {L1_3_L2_2_G2_MINI_ALU_BoothP_16,
                  L1_3_L2_2_G2_MINI_ALU_BoothP_15,
                  L1_3_L2_2_G2_MINI_ALU_BoothP_14,
                  L1_3_L2_2_G2_MINI_ALU_BoothP_13,
                  L1_3_L2_2_G2_MINI_ALU_BoothP_12,
                  L1_3_L2_2_G2_MINI_ALU_BoothP_11,
                  L1_3_L2_2_G2_MINI_ALU_BoothP_10,L1_3_L2_2_G2_MINI_ALU_BoothP_9
                  ,L1_3_L2_2_G2_MINI_ALU_BoothP_8,L1_3_L2_2_G2_MINI_ALU_BoothP_7
                  ,L1_3_L2_2_G2_MINI_ALU_BoothP_6,L1_3_L2_2_G2_MINI_ALU_BoothP_5
                  ,L1_3_L2_2_G2_MINI_ALU_BoothP_4,L1_3_L2_2_G2_MINI_ALU_BoothP_3
                  ,L1_3_L2_2_G2_MINI_ALU_BoothP_2,L1_3_L2_2_G2_MINI_ALU_BoothP_1
                  ,L1_3_L2_2_G2_MINI_ALU_BoothP_0}), .LargeWindowShifted ({
                  \$dummy [631],\$dummy [632],\$dummy [633],\$dummy [634],
                  \$dummy [635],\$dummy [636],\$dummy [637],\$dummy [638],
                  \$dummy [639],\$dummy [640],\$dummy [641],\$dummy [642],
                  \$dummy [643],\$dummy [644],\$dummy [645],\$dummy [646],
                  \$dummy [647]})) ;
    booth_adder_17_unfolded16 L1_3_L2_3_G2_MINI_ALU_BOOTH_ADDER (.AdderFirstOperand (
                              {L1ResultsLarge_10__16,L1ResultsLarge_10__15,
                              L1ResultsLarge_10__14,L1ResultsLarge_10__13,
                              L1ResultsLarge_10__12,L1ResultsLarge_10__11,
                              L1ResultsLarge_10__10,L1ResultsLarge_10__9,
                              L1ResultsLarge_10__8,L1ResultsLarge_10__7,
                              L1ResultsLarge_10__6,L1ResultsLarge_10__5,
                              L1ResultsLarge_10__4,L1ResultsLarge_10__3,
                              L1ResultsLarge_10__2,L1ResultsLarge_10__1,
                              L1ResultsLarge_10__0}), .AdderSecondOperand ({
                              L1ResultsLarge_11__16,L1ResultsLarge_11__15,
                              L1ResultsLarge_11__14,L1ResultsLarge_11__13,
                              L1ResultsLarge_11__12,L1ResultsLarge_11__11,
                              L1ResultsLarge_11__10,L1ResultsLarge_11__9,
                              L1ResultsLarge_11__8,L1ResultsLarge_11__7,
                              L1ResultsLarge_11__6,L1ResultsLarge_11__5,
                              L1ResultsLarge_11__4,L1ResultsLarge_11__3,
                              L1ResultsLarge_11__2,L1ResultsLarge_11__1,
                              L1ResultsLarge_11__0}), .BoothOperand ({
                              L1_3_L2_3_G2_MINI_ALU_BoothOperand_16,
                              L1_3_L2_3_G2_MINI_ALU_BoothOperand_15,
                              L1_3_L2_3_G2_MINI_ALU_BoothOperand_14,
                              L1_3_L2_3_G2_MINI_ALU_BoothOperand_13,
                              L1_3_L2_3_G2_MINI_ALU_BoothOperand_12,
                              L1_3_L2_3_G2_MINI_ALU_BoothOperand_11,
                              L1_3_L2_3_G2_MINI_ALU_BoothOperand_10,
                              L1_3_L2_3_G2_MINI_ALU_BoothOperand_9,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16}), .BoothP ({
                              L1_3_L2_3_G2_MINI_ALU_BoothP_16,
                              L1_3_L2_3_G2_MINI_ALU_BoothP_15,
                              L1_3_L2_3_G2_MINI_ALU_BoothP_14,
                              L1_3_L2_3_G2_MINI_ALU_BoothP_13,
                              L1_3_L2_3_G2_MINI_ALU_BoothP_12,
                              L1_3_L2_3_G2_MINI_ALU_BoothP_11,
                              L1_3_L2_3_G2_MINI_ALU_BoothP_10,
                              L1_3_L2_3_G2_MINI_ALU_BoothP_9,
                              L1_3_L2_3_G2_MINI_ALU_BoothP_8,
                              L1_3_L2_3_G2_MINI_ALU_BoothP_7,
                              L1_3_L2_3_G2_MINI_ALU_BoothP_6,
                              L1_3_L2_3_G2_MINI_ALU_BoothP_5,
                              L1_3_L2_3_G2_MINI_ALU_BoothP_4,
                              L1_3_L2_3_G2_MINI_ALU_BoothP_3,
                              L1_3_L2_3_G2_MINI_ALU_BoothP_2,
                              L1_3_L2_3_G2_MINI_ALU_BoothP_1,
                              L1_3_L2_3_G2_MINI_ALU_BoothP_0}), .SelOperand (
                              nx3284), .Operation (
                              L1_3_L2_3_G2_MINI_ALU_BoothXORCheck), .AdderResult (
                              {L2ResultsLarge_5__16,L2ResultsLarge_5__15,
                              L2ResultsLarge_5__14,L2ResultsLarge_5__13,
                              L2ResultsLarge_5__12,L2ResultsLarge_5__11,
                              L2ResultsLarge_5__10,L2ResultsLarge_5__9,
                              L2ResultsLarge_5__8,L2ResultsLarge_5__7,
                              L2ResultsLarge_5__6,L2ResultsLarge_5__5,
                              L2ResultsLarge_5__4,L2ResultsLarge_5__3,
                              L2ResultsLarge_5__2,L2ResultsLarge_5__1,
                              L2ResultsLarge_5__0}), .AdderBoothResult ({
                              \$dummy [648],
                              L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_15,
                              L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_14,
                              L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_13,
                              L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_12,
                              L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_11,
                              L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_10,
                              L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_9,
                              L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_8,
                              L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_7,
                              L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_6,
                              L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_5,
                              L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_4,
                              L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_3,
                              L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_2,
                              L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_1,
                              L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_0})) ;
    booth_unit_17 L1_3_L2_3_G2_MINI_ALU_BOOTH_UNIT (.CLK (CLK), .RST (RST), .Start (
                  Start), .Instr (Instr), .LoopingAndResultNotReady (nx3276), .Filter (
                  {FilterDin_3__3__7,FilterDin_3__3__6,FilterDin_3__3__5,
                  FilterDin_3__3__4,FilterDin_3__3__3,FilterDin_3__3__2,
                  FilterDin_3__3__1,FilterDin_3__3__0}), .Window ({
                  WindowDin_3__3__7,WindowDin_3__3__6,WindowDin_3__3__5,
                  WindowDin_3__3__4,WindowDin_3__3__3,WindowDin_3__3__2,
                  WindowDin_3__3__1,WindowDin_3__3__0}), .AdderBoothResult ({
                  L1FirstOperands_12__16,
                  L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_15,
                  L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_14,
                  L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_13,
                  L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_12,
                  L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_11,
                  L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_10,
                  L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_9,
                  L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_8,
                  L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_7,
                  L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_6,
                  L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_5,
                  L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_4,
                  L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_3,
                  L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_2,
                  L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_1,
                  L1_3_L2_3_G2_MINI_ALU_AdderBoothResult_0}), .BoothXORCheck (
                  L1_3_L2_3_G2_MINI_ALU_BoothXORCheck), .BoothResult ({
                  \$dummy [649],\$dummy [650],\$dummy [651],\$dummy [652],
                  \$dummy [653],\$dummy [654],\$dummy [655],\$dummy [656]}), .BoothAddingOperand (
                  {L1_3_L2_3_G2_MINI_ALU_BoothOperand_16,
                  L1_3_L2_3_G2_MINI_ALU_BoothOperand_15,
                  L1_3_L2_3_G2_MINI_ALU_BoothOperand_14,
                  L1_3_L2_3_G2_MINI_ALU_BoothOperand_13,
                  L1_3_L2_3_G2_MINI_ALU_BoothOperand_12,
                  L1_3_L2_3_G2_MINI_ALU_BoothOperand_11,
                  L1_3_L2_3_G2_MINI_ALU_BoothOperand_10,
                  L1_3_L2_3_G2_MINI_ALU_BoothOperand_9,\$dummy [657],
                  \$dummy [658],\$dummy [659],\$dummy [660],\$dummy [661],
                  \$dummy [662],\$dummy [663],\$dummy [664],\$dummy [665]}), .BoothP (
                  {L1_3_L2_3_G2_MINI_ALU_BoothP_16,
                  L1_3_L2_3_G2_MINI_ALU_BoothP_15,
                  L1_3_L2_3_G2_MINI_ALU_BoothP_14,
                  L1_3_L2_3_G2_MINI_ALU_BoothP_13,
                  L1_3_L2_3_G2_MINI_ALU_BoothP_12,
                  L1_3_L2_3_G2_MINI_ALU_BoothP_11,
                  L1_3_L2_3_G2_MINI_ALU_BoothP_10,L1_3_L2_3_G2_MINI_ALU_BoothP_9
                  ,L1_3_L2_3_G2_MINI_ALU_BoothP_8,L1_3_L2_3_G2_MINI_ALU_BoothP_7
                  ,L1_3_L2_3_G2_MINI_ALU_BoothP_6,L1_3_L2_3_G2_MINI_ALU_BoothP_5
                  ,L1_3_L2_3_G2_MINI_ALU_BoothP_4,L1_3_L2_3_G2_MINI_ALU_BoothP_3
                  ,L1_3_L2_3_G2_MINI_ALU_BoothP_2,L1_3_L2_3_G2_MINI_ALU_BoothP_1
                  ,L1_3_L2_3_G2_MINI_ALU_BoothP_0}), .LargeWindowShifted ({
                  \$dummy [666],\$dummy [667],\$dummy [668],\$dummy [669],
                  \$dummy [670],\$dummy [671],\$dummy [672],\$dummy [673],
                  \$dummy [674],\$dummy [675],\$dummy [676],\$dummy [677],
                  \$dummy [678],\$dummy [679],\$dummy [680],\$dummy [681],
                  \$dummy [682]})) ;
    booth_adder_17_unfolded16 L1_3_L2_4_G3_MINI_ALU_BOOTH_ADDER (.AdderFirstOperand (
                              {L2ResultsLarge_0__16,L2ResultsLarge_0__15,
                              L2ResultsLarge_0__14,L2ResultsLarge_0__13,
                              L2ResultsLarge_0__12,L2ResultsLarge_0__11,
                              L2ResultsLarge_0__10,L2ResultsLarge_0__9,
                              L2ResultsLarge_0__8,L2ResultsLarge_0__7,
                              L2ResultsLarge_0__6,L2ResultsLarge_0__5,
                              L2ResultsLarge_0__4,L2ResultsLarge_0__3,
                              L2ResultsLarge_0__2,L2ResultsLarge_0__1,
                              L2ResultsLarge_0__0}), .AdderSecondOperand ({
                              L2ResultsLarge_1__16,L2ResultsLarge_1__15,
                              L2ResultsLarge_1__14,L2ResultsLarge_1__13,
                              L2ResultsLarge_1__12,L2ResultsLarge_1__11,
                              L2ResultsLarge_1__10,L2ResultsLarge_1__9,
                              L2ResultsLarge_1__8,L2ResultsLarge_1__7,
                              L2ResultsLarge_1__6,L2ResultsLarge_1__5,
                              L2ResultsLarge_1__4,L2ResultsLarge_1__3,
                              L2ResultsLarge_1__2,L2ResultsLarge_1__1,
                              L2ResultsLarge_1__0}), .BoothOperand ({
                              L1_3_L2_4_G3_MINI_ALU_BoothOperand_16,
                              L1_3_L2_4_G3_MINI_ALU_BoothOperand_15,
                              L1_3_L2_4_G3_MINI_ALU_BoothOperand_14,
                              L1_3_L2_4_G3_MINI_ALU_BoothOperand_13,
                              L1_3_L2_4_G3_MINI_ALU_BoothOperand_12,
                              L1_3_L2_4_G3_MINI_ALU_BoothOperand_11,
                              L1_3_L2_4_G3_MINI_ALU_BoothOperand_10,
                              L1_3_L2_4_G3_MINI_ALU_BoothOperand_9,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16}), .BoothP ({
                              L1_3_L2_4_G3_MINI_ALU_BoothP_16,
                              L1_3_L2_4_G3_MINI_ALU_BoothP_15,
                              L1_3_L2_4_G3_MINI_ALU_BoothP_14,
                              L1_3_L2_4_G3_MINI_ALU_BoothP_13,
                              L1_3_L2_4_G3_MINI_ALU_BoothP_12,
                              L1_3_L2_4_G3_MINI_ALU_BoothP_11,
                              L1_3_L2_4_G3_MINI_ALU_BoothP_10,
                              L1_3_L2_4_G3_MINI_ALU_BoothP_9,
                              L1_3_L2_4_G3_MINI_ALU_BoothP_8,
                              L1_3_L2_4_G3_MINI_ALU_BoothP_7,
                              L1_3_L2_4_G3_MINI_ALU_BoothP_6,
                              L1_3_L2_4_G3_MINI_ALU_BoothP_5,
                              L1_3_L2_4_G3_MINI_ALU_BoothP_4,
                              L1_3_L2_4_G3_MINI_ALU_BoothP_3,
                              L1_3_L2_4_G3_MINI_ALU_BoothP_2,
                              L1_3_L2_4_G3_MINI_ALU_BoothP_1,
                              L1_3_L2_4_G3_MINI_ALU_BoothP_0}), .SelOperand (
                              nx3284), .Operation (
                              L1_3_L2_4_G3_MINI_ALU_BoothXORCheck), .AdderResult (
                              {L3ResultsLarge_0__16,L3ResultsLarge_0__15,
                              L3ResultsLarge_0__14,L3ResultsLarge_0__13,
                              L3ResultsLarge_0__12,L3ResultsLarge_0__11,
                              L3ResultsLarge_0__10,L3ResultsLarge_0__9,
                              L3ResultsLarge_0__8,L3ResultsLarge_0__7,
                              L3ResultsLarge_0__6,L3ResultsLarge_0__5,
                              L3ResultsLarge_0__4,L3ResultsLarge_0__3,
                              L3ResultsLarge_0__2,L3ResultsLarge_0__1,
                              L3ResultsLarge_0__0}), .AdderBoothResult ({
                              \$dummy [683],
                              L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_15,
                              L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_14,
                              L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_13,
                              L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_12,
                              L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_11,
                              L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_10,
                              L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_9,
                              L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_8,
                              L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_7,
                              L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_6,
                              L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_5,
                              L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_4,
                              L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_3,
                              L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_2,
                              L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_1,
                              L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_0})) ;
    booth_unit_17 L1_3_L2_4_G3_MINI_ALU_BOOTH_UNIT (.CLK (CLK), .RST (RST), .Start (
                  Start), .Instr (Instr), .LoopingAndResultNotReady (nx3276), .Filter (
                  {FilterDin_3__4__7,FilterDin_3__4__6,FilterDin_3__4__5,
                  FilterDin_3__4__4,FilterDin_3__4__3,FilterDin_3__4__2,
                  FilterDin_3__4__1,FilterDin_3__4__0}), .Window ({
                  WindowDin_3__4__7,WindowDin_3__4__6,WindowDin_3__4__5,
                  WindowDin_3__4__4,WindowDin_3__4__3,WindowDin_3__4__2,
                  WindowDin_3__4__1,WindowDin_3__4__0}), .AdderBoothResult ({
                  L1FirstOperands_12__16,
                  L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_15,
                  L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_14,
                  L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_13,
                  L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_12,
                  L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_11,
                  L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_10,
                  L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_9,
                  L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_8,
                  L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_7,
                  L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_6,
                  L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_5,
                  L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_4,
                  L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_3,
                  L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_2,
                  L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_1,
                  L1_3_L2_4_G3_MINI_ALU_AdderBoothResult_0}), .BoothXORCheck (
                  L1_3_L2_4_G3_MINI_ALU_BoothXORCheck), .BoothResult ({
                  \$dummy [684],\$dummy [685],\$dummy [686],\$dummy [687],
                  \$dummy [688],\$dummy [689],\$dummy [690],\$dummy [691]}), .BoothAddingOperand (
                  {L1_3_L2_4_G3_MINI_ALU_BoothOperand_16,
                  L1_3_L2_4_G3_MINI_ALU_BoothOperand_15,
                  L1_3_L2_4_G3_MINI_ALU_BoothOperand_14,
                  L1_3_L2_4_G3_MINI_ALU_BoothOperand_13,
                  L1_3_L2_4_G3_MINI_ALU_BoothOperand_12,
                  L1_3_L2_4_G3_MINI_ALU_BoothOperand_11,
                  L1_3_L2_4_G3_MINI_ALU_BoothOperand_10,
                  L1_3_L2_4_G3_MINI_ALU_BoothOperand_9,\$dummy [692],
                  \$dummy [693],\$dummy [694],\$dummy [695],\$dummy [696],
                  \$dummy [697],\$dummy [698],\$dummy [699],\$dummy [700]}), .BoothP (
                  {L1_3_L2_4_G3_MINI_ALU_BoothP_16,
                  L1_3_L2_4_G3_MINI_ALU_BoothP_15,
                  L1_3_L2_4_G3_MINI_ALU_BoothP_14,
                  L1_3_L2_4_G3_MINI_ALU_BoothP_13,
                  L1_3_L2_4_G3_MINI_ALU_BoothP_12,
                  L1_3_L2_4_G3_MINI_ALU_BoothP_11,
                  L1_3_L2_4_G3_MINI_ALU_BoothP_10,L1_3_L2_4_G3_MINI_ALU_BoothP_9
                  ,L1_3_L2_4_G3_MINI_ALU_BoothP_8,L1_3_L2_4_G3_MINI_ALU_BoothP_7
                  ,L1_3_L2_4_G3_MINI_ALU_BoothP_6,L1_3_L2_4_G3_MINI_ALU_BoothP_5
                  ,L1_3_L2_4_G3_MINI_ALU_BoothP_4,L1_3_L2_4_G3_MINI_ALU_BoothP_3
                  ,L1_3_L2_4_G3_MINI_ALU_BoothP_2,L1_3_L2_4_G3_MINI_ALU_BoothP_1
                  ,L1_3_L2_4_G3_MINI_ALU_BoothP_0}), .LargeWindowShifted ({
                  \$dummy [701],\$dummy [702],\$dummy [703],\$dummy [704],
                  \$dummy [705],\$dummy [706],\$dummy [707],\$dummy [708],
                  \$dummy [709],\$dummy [710],\$dummy [711],\$dummy [712],
                  \$dummy [713],\$dummy [714],\$dummy [715],\$dummy [716],
                  \$dummy [717]})) ;
    booth_adder_17_unfolded16 L1_4_L2_0_G3_MINI_ALU_BOOTH_ADDER (.AdderFirstOperand (
                              {L2ResultsLarge_2__16,L2ResultsLarge_2__15,
                              L2ResultsLarge_2__14,L2ResultsLarge_2__13,
                              L2ResultsLarge_2__12,L2ResultsLarge_2__11,
                              L2ResultsLarge_2__10,L2ResultsLarge_2__9,
                              L2ResultsLarge_2__8,L2ResultsLarge_2__7,
                              L2ResultsLarge_2__6,L2ResultsLarge_2__5,
                              L2ResultsLarge_2__4,L2ResultsLarge_2__3,
                              L2ResultsLarge_2__2,L2ResultsLarge_2__1,
                              L2ResultsLarge_2__0}), .AdderSecondOperand ({
                              L2ResultsLarge_3__16,L2ResultsLarge_3__15,
                              L2ResultsLarge_3__14,L2ResultsLarge_3__13,
                              L2ResultsLarge_3__12,L2ResultsLarge_3__11,
                              L2ResultsLarge_3__10,L2ResultsLarge_3__9,
                              L2ResultsLarge_3__8,L2ResultsLarge_3__7,
                              L2ResultsLarge_3__6,L2ResultsLarge_3__5,
                              L2ResultsLarge_3__4,L2ResultsLarge_3__3,
                              L2ResultsLarge_3__2,L2ResultsLarge_3__1,
                              L2ResultsLarge_3__0}), .BoothOperand ({
                              L1_4_L2_0_G3_MINI_ALU_BoothOperand_16,
                              L1_4_L2_0_G3_MINI_ALU_BoothOperand_15,
                              L1_4_L2_0_G3_MINI_ALU_BoothOperand_14,
                              L1_4_L2_0_G3_MINI_ALU_BoothOperand_13,
                              L1_4_L2_0_G3_MINI_ALU_BoothOperand_12,
                              L1_4_L2_0_G3_MINI_ALU_BoothOperand_11,
                              L1_4_L2_0_G3_MINI_ALU_BoothOperand_10,
                              L1_4_L2_0_G3_MINI_ALU_BoothOperand_9,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16}), .BoothP ({
                              L1_4_L2_0_G3_MINI_ALU_BoothP_16,
                              L1_4_L2_0_G3_MINI_ALU_BoothP_15,
                              L1_4_L2_0_G3_MINI_ALU_BoothP_14,
                              L1_4_L2_0_G3_MINI_ALU_BoothP_13,
                              L1_4_L2_0_G3_MINI_ALU_BoothP_12,
                              L1_4_L2_0_G3_MINI_ALU_BoothP_11,
                              L1_4_L2_0_G3_MINI_ALU_BoothP_10,
                              L1_4_L2_0_G3_MINI_ALU_BoothP_9,
                              L1_4_L2_0_G3_MINI_ALU_BoothP_8,
                              L1_4_L2_0_G3_MINI_ALU_BoothP_7,
                              L1_4_L2_0_G3_MINI_ALU_BoothP_6,
                              L1_4_L2_0_G3_MINI_ALU_BoothP_5,
                              L1_4_L2_0_G3_MINI_ALU_BoothP_4,
                              L1_4_L2_0_G3_MINI_ALU_BoothP_3,
                              L1_4_L2_0_G3_MINI_ALU_BoothP_2,
                              L1_4_L2_0_G3_MINI_ALU_BoothP_1,
                              L1_4_L2_0_G3_MINI_ALU_BoothP_0}), .SelOperand (
                              nx3284), .Operation (
                              L1_4_L2_0_G3_MINI_ALU_BoothXORCheck), .AdderResult (
                              {L3ResultsLarge_1__16,L3ResultsLarge_1__15,
                              L3ResultsLarge_1__14,L3ResultsLarge_1__13,
                              L3ResultsLarge_1__12,L3ResultsLarge_1__11,
                              L3ResultsLarge_1__10,L3ResultsLarge_1__9,
                              L3ResultsLarge_1__8,L3ResultsLarge_1__7,
                              L3ResultsLarge_1__6,L3ResultsLarge_1__5,
                              L3ResultsLarge_1__4,L3ResultsLarge_1__3,
                              L3ResultsLarge_1__2,L3ResultsLarge_1__1,
                              L3ResultsLarge_1__0}), .AdderBoothResult ({
                              \$dummy [718],
                              L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_15,
                              L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_14,
                              L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_13,
                              L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_12,
                              L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_11,
                              L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_10,
                              L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_9,
                              L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_8,
                              L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_7,
                              L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_6,
                              L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_5,
                              L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_4,
                              L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_3,
                              L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_2,
                              L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_1,
                              L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_0})) ;
    booth_unit_17 L1_4_L2_0_G3_MINI_ALU_BOOTH_UNIT (.CLK (CLK), .RST (RST), .Start (
                  Start), .Instr (Instr), .LoopingAndResultNotReady (nx3276), .Filter (
                  {FilterDin_4__0__7,FilterDin_4__0__6,FilterDin_4__0__5,
                  FilterDin_4__0__4,FilterDin_4__0__3,FilterDin_4__0__2,
                  FilterDin_4__0__1,FilterDin_4__0__0}), .Window ({
                  WindowDin_4__0__7,WindowDin_4__0__6,WindowDin_4__0__5,
                  WindowDin_4__0__4,WindowDin_4__0__3,WindowDin_4__0__2,
                  WindowDin_4__0__1,WindowDin_4__0__0}), .AdderBoothResult ({
                  L1FirstOperands_12__16,
                  L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_15,
                  L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_14,
                  L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_13,
                  L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_12,
                  L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_11,
                  L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_10,
                  L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_9,
                  L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_8,
                  L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_7,
                  L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_6,
                  L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_5,
                  L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_4,
                  L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_3,
                  L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_2,
                  L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_1,
                  L1_4_L2_0_G3_MINI_ALU_AdderBoothResult_0}), .BoothXORCheck (
                  L1_4_L2_0_G3_MINI_ALU_BoothXORCheck), .BoothResult ({
                  \$dummy [719],\$dummy [720],\$dummy [721],\$dummy [722],
                  \$dummy [723],\$dummy [724],\$dummy [725],\$dummy [726]}), .BoothAddingOperand (
                  {L1_4_L2_0_G3_MINI_ALU_BoothOperand_16,
                  L1_4_L2_0_G3_MINI_ALU_BoothOperand_15,
                  L1_4_L2_0_G3_MINI_ALU_BoothOperand_14,
                  L1_4_L2_0_G3_MINI_ALU_BoothOperand_13,
                  L1_4_L2_0_G3_MINI_ALU_BoothOperand_12,
                  L1_4_L2_0_G3_MINI_ALU_BoothOperand_11,
                  L1_4_L2_0_G3_MINI_ALU_BoothOperand_10,
                  L1_4_L2_0_G3_MINI_ALU_BoothOperand_9,\$dummy [727],
                  \$dummy [728],\$dummy [729],\$dummy [730],\$dummy [731],
                  \$dummy [732],\$dummy [733],\$dummy [734],\$dummy [735]}), .BoothP (
                  {L1_4_L2_0_G3_MINI_ALU_BoothP_16,
                  L1_4_L2_0_G3_MINI_ALU_BoothP_15,
                  L1_4_L2_0_G3_MINI_ALU_BoothP_14,
                  L1_4_L2_0_G3_MINI_ALU_BoothP_13,
                  L1_4_L2_0_G3_MINI_ALU_BoothP_12,
                  L1_4_L2_0_G3_MINI_ALU_BoothP_11,
                  L1_4_L2_0_G3_MINI_ALU_BoothP_10,L1_4_L2_0_G3_MINI_ALU_BoothP_9
                  ,L1_4_L2_0_G3_MINI_ALU_BoothP_8,L1_4_L2_0_G3_MINI_ALU_BoothP_7
                  ,L1_4_L2_0_G3_MINI_ALU_BoothP_6,L1_4_L2_0_G3_MINI_ALU_BoothP_5
                  ,L1_4_L2_0_G3_MINI_ALU_BoothP_4,L1_4_L2_0_G3_MINI_ALU_BoothP_3
                  ,L1_4_L2_0_G3_MINI_ALU_BoothP_2,L1_4_L2_0_G3_MINI_ALU_BoothP_1
                  ,L1_4_L2_0_G3_MINI_ALU_BoothP_0}), .LargeWindowShifted ({
                  \$dummy [736],\$dummy [737],\$dummy [738],\$dummy [739],
                  \$dummy [740],\$dummy [741],\$dummy [742],\$dummy [743],
                  \$dummy [744],\$dummy [745],\$dummy [746],\$dummy [747],
                  \$dummy [748],\$dummy [749],\$dummy [750],\$dummy [751],
                  \$dummy [752]})) ;
    booth_adder_17_unfolded16 L1_4_L2_1_G3_MINI_ALU_BOOTH_ADDER (.AdderFirstOperand (
                              {L2ResultsLarge_4__16,L2ResultsLarge_4__15,
                              L2ResultsLarge_4__14,L2ResultsLarge_4__13,
                              L2ResultsLarge_4__12,L2ResultsLarge_4__11,
                              L2ResultsLarge_4__10,L2ResultsLarge_4__9,
                              L2ResultsLarge_4__8,L2ResultsLarge_4__7,
                              L2ResultsLarge_4__6,L2ResultsLarge_4__5,
                              L2ResultsLarge_4__4,L2ResultsLarge_4__3,
                              L2ResultsLarge_4__2,L2ResultsLarge_4__1,
                              L2ResultsLarge_4__0}), .AdderSecondOperand ({
                              L2ResultsLarge_5__16,L2ResultsLarge_5__15,
                              L2ResultsLarge_5__14,L2ResultsLarge_5__13,
                              L2ResultsLarge_5__12,L2ResultsLarge_5__11,
                              L2ResultsLarge_5__10,L2ResultsLarge_5__9,
                              L2ResultsLarge_5__8,L2ResultsLarge_5__7,
                              L2ResultsLarge_5__6,L2ResultsLarge_5__5,
                              L2ResultsLarge_5__4,L2ResultsLarge_5__3,
                              L2ResultsLarge_5__2,L2ResultsLarge_5__1,
                              L2ResultsLarge_5__0}), .BoothOperand ({
                              L1_4_L2_1_G3_MINI_ALU_BoothOperand_16,
                              L1_4_L2_1_G3_MINI_ALU_BoothOperand_15,
                              L1_4_L2_1_G3_MINI_ALU_BoothOperand_14,
                              L1_4_L2_1_G3_MINI_ALU_BoothOperand_13,
                              L1_4_L2_1_G3_MINI_ALU_BoothOperand_12,
                              L1_4_L2_1_G3_MINI_ALU_BoothOperand_11,
                              L1_4_L2_1_G3_MINI_ALU_BoothOperand_10,
                              L1_4_L2_1_G3_MINI_ALU_BoothOperand_9,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16}), .BoothP ({
                              L1_4_L2_1_G3_MINI_ALU_BoothP_16,
                              L1_4_L2_1_G3_MINI_ALU_BoothP_15,
                              L1_4_L2_1_G3_MINI_ALU_BoothP_14,
                              L1_4_L2_1_G3_MINI_ALU_BoothP_13,
                              L1_4_L2_1_G3_MINI_ALU_BoothP_12,
                              L1_4_L2_1_G3_MINI_ALU_BoothP_11,
                              L1_4_L2_1_G3_MINI_ALU_BoothP_10,
                              L1_4_L2_1_G3_MINI_ALU_BoothP_9,
                              L1_4_L2_1_G3_MINI_ALU_BoothP_8,
                              L1_4_L2_1_G3_MINI_ALU_BoothP_7,
                              L1_4_L2_1_G3_MINI_ALU_BoothP_6,
                              L1_4_L2_1_G3_MINI_ALU_BoothP_5,
                              L1_4_L2_1_G3_MINI_ALU_BoothP_4,
                              L1_4_L2_1_G3_MINI_ALU_BoothP_3,
                              L1_4_L2_1_G3_MINI_ALU_BoothP_2,
                              L1_4_L2_1_G3_MINI_ALU_BoothP_1,
                              L1_4_L2_1_G3_MINI_ALU_BoothP_0}), .SelOperand (
                              nx3286), .Operation (
                              L1_4_L2_1_G3_MINI_ALU_BoothXORCheck), .AdderResult (
                              {L3ResultsLarge_2__16,L3ResultsLarge_2__15,
                              L3ResultsLarge_2__14,L3ResultsLarge_2__13,
                              L3ResultsLarge_2__12,L3ResultsLarge_2__11,
                              L3ResultsLarge_2__10,L3ResultsLarge_2__9,
                              L3ResultsLarge_2__8,L3ResultsLarge_2__7,
                              L3ResultsLarge_2__6,L3ResultsLarge_2__5,
                              L3ResultsLarge_2__4,L3ResultsLarge_2__3,
                              L3ResultsLarge_2__2,L3ResultsLarge_2__1,
                              L3ResultsLarge_2__0}), .AdderBoothResult ({
                              \$dummy [753],
                              L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_15,
                              L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_14,
                              L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_13,
                              L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_12,
                              L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_11,
                              L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_10,
                              L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_9,
                              L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_8,
                              L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_7,
                              L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_6,
                              L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_5,
                              L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_4,
                              L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_3,
                              L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_2,
                              L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_1,
                              L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_0})) ;
    booth_unit_17 L1_4_L2_1_G3_MINI_ALU_BOOTH_UNIT (.CLK (CLK), .RST (RST), .Start (
                  Start), .Instr (Instr), .LoopingAndResultNotReady (nx3278), .Filter (
                  {FilterDin_4__1__7,FilterDin_4__1__6,FilterDin_4__1__5,
                  FilterDin_4__1__4,FilterDin_4__1__3,FilterDin_4__1__2,
                  FilterDin_4__1__1,FilterDin_4__1__0}), .Window ({
                  WindowDin_4__1__7,WindowDin_4__1__6,WindowDin_4__1__5,
                  WindowDin_4__1__4,WindowDin_4__1__3,WindowDin_4__1__2,
                  WindowDin_4__1__1,WindowDin_4__1__0}), .AdderBoothResult ({
                  L1FirstOperands_12__16,
                  L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_15,
                  L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_14,
                  L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_13,
                  L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_12,
                  L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_11,
                  L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_10,
                  L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_9,
                  L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_8,
                  L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_7,
                  L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_6,
                  L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_5,
                  L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_4,
                  L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_3,
                  L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_2,
                  L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_1,
                  L1_4_L2_1_G3_MINI_ALU_AdderBoothResult_0}), .BoothXORCheck (
                  L1_4_L2_1_G3_MINI_ALU_BoothXORCheck), .BoothResult ({
                  \$dummy [754],\$dummy [755],\$dummy [756],\$dummy [757],
                  \$dummy [758],\$dummy [759],\$dummy [760],\$dummy [761]}), .BoothAddingOperand (
                  {L1_4_L2_1_G3_MINI_ALU_BoothOperand_16,
                  L1_4_L2_1_G3_MINI_ALU_BoothOperand_15,
                  L1_4_L2_1_G3_MINI_ALU_BoothOperand_14,
                  L1_4_L2_1_G3_MINI_ALU_BoothOperand_13,
                  L1_4_L2_1_G3_MINI_ALU_BoothOperand_12,
                  L1_4_L2_1_G3_MINI_ALU_BoothOperand_11,
                  L1_4_L2_1_G3_MINI_ALU_BoothOperand_10,
                  L1_4_L2_1_G3_MINI_ALU_BoothOperand_9,\$dummy [762],
                  \$dummy [763],\$dummy [764],\$dummy [765],\$dummy [766],
                  \$dummy [767],\$dummy [768],\$dummy [769],\$dummy [770]}), .BoothP (
                  {L1_4_L2_1_G3_MINI_ALU_BoothP_16,
                  L1_4_L2_1_G3_MINI_ALU_BoothP_15,
                  L1_4_L2_1_G3_MINI_ALU_BoothP_14,
                  L1_4_L2_1_G3_MINI_ALU_BoothP_13,
                  L1_4_L2_1_G3_MINI_ALU_BoothP_12,
                  L1_4_L2_1_G3_MINI_ALU_BoothP_11,
                  L1_4_L2_1_G3_MINI_ALU_BoothP_10,L1_4_L2_1_G3_MINI_ALU_BoothP_9
                  ,L1_4_L2_1_G3_MINI_ALU_BoothP_8,L1_4_L2_1_G3_MINI_ALU_BoothP_7
                  ,L1_4_L2_1_G3_MINI_ALU_BoothP_6,L1_4_L2_1_G3_MINI_ALU_BoothP_5
                  ,L1_4_L2_1_G3_MINI_ALU_BoothP_4,L1_4_L2_1_G3_MINI_ALU_BoothP_3
                  ,L1_4_L2_1_G3_MINI_ALU_BoothP_2,L1_4_L2_1_G3_MINI_ALU_BoothP_1
                  ,L1_4_L2_1_G3_MINI_ALU_BoothP_0}), .LargeWindowShifted ({
                  \$dummy [771],\$dummy [772],\$dummy [773],\$dummy [774],
                  \$dummy [775],\$dummy [776],\$dummy [777],\$dummy [778],
                  \$dummy [779],\$dummy [780],\$dummy [781],\$dummy [782],
                  \$dummy [783],\$dummy [784],\$dummy [785],\$dummy [786],
                  \$dummy [787]})) ;
    booth_adder_17_unfolded16 L1_4_L2_2_G4_MINI_ALU_BOOTH_ADDER (.AdderFirstOperand (
                              {L3ResultsLarge_0__16,L3ResultsLarge_0__15,
                              L3ResultsLarge_0__14,L3ResultsLarge_0__13,
                              L3ResultsLarge_0__12,L3ResultsLarge_0__11,
                              L3ResultsLarge_0__10,L3ResultsLarge_0__9,
                              L3ResultsLarge_0__8,L3ResultsLarge_0__7,
                              L3ResultsLarge_0__6,L3ResultsLarge_0__5,
                              L3ResultsLarge_0__4,L3ResultsLarge_0__3,
                              L3ResultsLarge_0__2,L3ResultsLarge_0__1,
                              L3ResultsLarge_0__0}), .AdderSecondOperand ({
                              L3ResultsLarge_1__16,L3ResultsLarge_1__15,
                              L3ResultsLarge_1__14,L3ResultsLarge_1__13,
                              L3ResultsLarge_1__12,L3ResultsLarge_1__11,
                              L3ResultsLarge_1__10,L3ResultsLarge_1__9,
                              L3ResultsLarge_1__8,L3ResultsLarge_1__7,
                              L3ResultsLarge_1__6,L3ResultsLarge_1__5,
                              L3ResultsLarge_1__4,L3ResultsLarge_1__3,
                              L3ResultsLarge_1__2,L3ResultsLarge_1__1,
                              L3ResultsLarge_1__0}), .BoothOperand ({
                              L1_4_L2_2_G4_MINI_ALU_BoothOperand_16,
                              L1_4_L2_2_G4_MINI_ALU_BoothOperand_15,
                              L1_4_L2_2_G4_MINI_ALU_BoothOperand_14,
                              L1_4_L2_2_G4_MINI_ALU_BoothOperand_13,
                              L1_4_L2_2_G4_MINI_ALU_BoothOperand_12,
                              L1_4_L2_2_G4_MINI_ALU_BoothOperand_11,
                              L1_4_L2_2_G4_MINI_ALU_BoothOperand_10,
                              L1_4_L2_2_G4_MINI_ALU_BoothOperand_9,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16}), .BoothP ({
                              L1_4_L2_2_G4_MINI_ALU_BoothP_16,
                              L1_4_L2_2_G4_MINI_ALU_BoothP_15,
                              L1_4_L2_2_G4_MINI_ALU_BoothP_14,
                              L1_4_L2_2_G4_MINI_ALU_BoothP_13,
                              L1_4_L2_2_G4_MINI_ALU_BoothP_12,
                              L1_4_L2_2_G4_MINI_ALU_BoothP_11,
                              L1_4_L2_2_G4_MINI_ALU_BoothP_10,
                              L1_4_L2_2_G4_MINI_ALU_BoothP_9,
                              L1_4_L2_2_G4_MINI_ALU_BoothP_8,
                              L1_4_L2_2_G4_MINI_ALU_BoothP_7,
                              L1_4_L2_2_G4_MINI_ALU_BoothP_6,
                              L1_4_L2_2_G4_MINI_ALU_BoothP_5,
                              L1_4_L2_2_G4_MINI_ALU_BoothP_4,
                              L1_4_L2_2_G4_MINI_ALU_BoothP_3,
                              L1_4_L2_2_G4_MINI_ALU_BoothP_2,
                              L1_4_L2_2_G4_MINI_ALU_BoothP_1,
                              L1_4_L2_2_G4_MINI_ALU_BoothP_0}), .SelOperand (
                              nx3286), .Operation (
                              L1_4_L2_2_G4_MINI_ALU_BoothXORCheck), .AdderResult (
                              {L4ResultsLarge_0__16,L4ResultsLarge_0__15,
                              L4ResultsLarge_0__14,L4ResultsLarge_0__13,
                              L4ResultsLarge_0__12,L4ResultsLarge_0__11,
                              L4ResultsLarge_0__10,L4ResultsLarge_0__9,
                              L4ResultsLarge_0__8,L4ResultsLarge_0__7,
                              L4ResultsLarge_0__6,L4ResultsLarge_0__5,
                              L4ResultsLarge_0__4,L4ResultsLarge_0__3,
                              L4ResultsLarge_0__2,L4ResultsLarge_0__1,
                              L4ResultsLarge_0__0}), .AdderBoothResult ({
                              \$dummy [788],
                              L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_15,
                              L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_14,
                              L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_13,
                              L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_12,
                              L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_11,
                              L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_10,
                              L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_9,
                              L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_8,
                              L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_7,
                              L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_6,
                              L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_5,
                              L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_4,
                              L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_3,
                              L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_2,
                              L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_1,
                              L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_0})) ;
    booth_unit_17 L1_4_L2_2_G4_MINI_ALU_BOOTH_UNIT (.CLK (CLK), .RST (RST), .Start (
                  Start), .Instr (Instr), .LoopingAndResultNotReady (nx3278), .Filter (
                  {FilterDin_4__2__7,FilterDin_4__2__6,FilterDin_4__2__5,
                  FilterDin_4__2__4,FilterDin_4__2__3,FilterDin_4__2__2,
                  FilterDin_4__2__1,FilterDin_4__2__0}), .Window ({
                  WindowDin_4__2__7,WindowDin_4__2__6,WindowDin_4__2__5,
                  WindowDin_4__2__4,WindowDin_4__2__3,WindowDin_4__2__2,
                  WindowDin_4__2__1,WindowDin_4__2__0}), .AdderBoothResult ({
                  L1FirstOperands_12__16,
                  L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_15,
                  L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_14,
                  L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_13,
                  L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_12,
                  L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_11,
                  L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_10,
                  L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_9,
                  L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_8,
                  L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_7,
                  L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_6,
                  L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_5,
                  L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_4,
                  L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_3,
                  L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_2,
                  L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_1,
                  L1_4_L2_2_G4_MINI_ALU_AdderBoothResult_0}), .BoothXORCheck (
                  L1_4_L2_2_G4_MINI_ALU_BoothXORCheck), .BoothResult ({
                  \$dummy [789],\$dummy [790],\$dummy [791],\$dummy [792],
                  \$dummy [793],\$dummy [794],\$dummy [795],\$dummy [796]}), .BoothAddingOperand (
                  {L1_4_L2_2_G4_MINI_ALU_BoothOperand_16,
                  L1_4_L2_2_G4_MINI_ALU_BoothOperand_15,
                  L1_4_L2_2_G4_MINI_ALU_BoothOperand_14,
                  L1_4_L2_2_G4_MINI_ALU_BoothOperand_13,
                  L1_4_L2_2_G4_MINI_ALU_BoothOperand_12,
                  L1_4_L2_2_G4_MINI_ALU_BoothOperand_11,
                  L1_4_L2_2_G4_MINI_ALU_BoothOperand_10,
                  L1_4_L2_2_G4_MINI_ALU_BoothOperand_9,\$dummy [797],
                  \$dummy [798],\$dummy [799],\$dummy [800],\$dummy [801],
                  \$dummy [802],\$dummy [803],\$dummy [804],\$dummy [805]}), .BoothP (
                  {L1_4_L2_2_G4_MINI_ALU_BoothP_16,
                  L1_4_L2_2_G4_MINI_ALU_BoothP_15,
                  L1_4_L2_2_G4_MINI_ALU_BoothP_14,
                  L1_4_L2_2_G4_MINI_ALU_BoothP_13,
                  L1_4_L2_2_G4_MINI_ALU_BoothP_12,
                  L1_4_L2_2_G4_MINI_ALU_BoothP_11,
                  L1_4_L2_2_G4_MINI_ALU_BoothP_10,L1_4_L2_2_G4_MINI_ALU_BoothP_9
                  ,L1_4_L2_2_G4_MINI_ALU_BoothP_8,L1_4_L2_2_G4_MINI_ALU_BoothP_7
                  ,L1_4_L2_2_G4_MINI_ALU_BoothP_6,L1_4_L2_2_G4_MINI_ALU_BoothP_5
                  ,L1_4_L2_2_G4_MINI_ALU_BoothP_4,L1_4_L2_2_G4_MINI_ALU_BoothP_3
                  ,L1_4_L2_2_G4_MINI_ALU_BoothP_2,L1_4_L2_2_G4_MINI_ALU_BoothP_1
                  ,L1_4_L2_2_G4_MINI_ALU_BoothP_0}), .LargeWindowShifted ({
                  \$dummy [806],\$dummy [807],\$dummy [808],\$dummy [809],
                  \$dummy [810],\$dummy [811],\$dummy [812],\$dummy [813],
                  \$dummy [814],\$dummy [815],\$dummy [816],\$dummy [817],
                  \$dummy [818],\$dummy [819],\$dummy [820],\$dummy [821],
                  \$dummy [822]})) ;
    booth_adder_17_unfolded16 L1_4_L2_3_G5_MINI_ALU_BOOTH_ADDER (.AdderFirstOperand (
                              {L4ResultsLarge_0__16,L4ResultsLarge_0__15,
                              L4ResultsLarge_0__14,L4ResultsLarge_0__13,
                              L4ResultsLarge_0__12,L4ResultsLarge_0__11,
                              L4ResultsLarge_0__10,L4ResultsLarge_0__9,
                              L4ResultsLarge_0__8,L4ResultsLarge_0__7,
                              L4ResultsLarge_0__6,L4ResultsLarge_0__5,
                              L4ResultsLarge_0__4,L4ResultsLarge_0__3,
                              L4ResultsLarge_0__2,L4ResultsLarge_0__1,
                              L4ResultsLarge_0__0}), .AdderSecondOperand ({
                              L3ResultsLarge_2__16,L3ResultsLarge_2__15,
                              L3ResultsLarge_2__14,L3ResultsLarge_2__13,
                              L3ResultsLarge_2__12,L3ResultsLarge_2__11,
                              L3ResultsLarge_2__10,L3ResultsLarge_2__9,
                              L3ResultsLarge_2__8,L3ResultsLarge_2__7,
                              L3ResultsLarge_2__6,L3ResultsLarge_2__5,
                              L3ResultsLarge_2__4,L3ResultsLarge_2__3,
                              L3ResultsLarge_2__2,L3ResultsLarge_2__1,
                              L3ResultsLarge_2__0}), .BoothOperand ({
                              L1_4_L2_3_G5_MINI_ALU_BoothOperand_16,
                              L1_4_L2_3_G5_MINI_ALU_BoothOperand_15,
                              L1_4_L2_3_G5_MINI_ALU_BoothOperand_14,
                              L1_4_L2_3_G5_MINI_ALU_BoothOperand_13,
                              L1_4_L2_3_G5_MINI_ALU_BoothOperand_12,
                              L1_4_L2_3_G5_MINI_ALU_BoothOperand_11,
                              L1_4_L2_3_G5_MINI_ALU_BoothOperand_10,
                              L1_4_L2_3_G5_MINI_ALU_BoothOperand_9,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16}), .BoothP ({
                              L1_4_L2_3_G5_MINI_ALU_BoothP_16,
                              L1_4_L2_3_G5_MINI_ALU_BoothP_15,
                              L1_4_L2_3_G5_MINI_ALU_BoothP_14,
                              L1_4_L2_3_G5_MINI_ALU_BoothP_13,
                              L1_4_L2_3_G5_MINI_ALU_BoothP_12,
                              L1_4_L2_3_G5_MINI_ALU_BoothP_11,
                              L1_4_L2_3_G5_MINI_ALU_BoothP_10,
                              L1_4_L2_3_G5_MINI_ALU_BoothP_9,
                              L1_4_L2_3_G5_MINI_ALU_BoothP_8,
                              L1_4_L2_3_G5_MINI_ALU_BoothP_7,
                              L1_4_L2_3_G5_MINI_ALU_BoothP_6,
                              L1_4_L2_3_G5_MINI_ALU_BoothP_5,
                              L1_4_L2_3_G5_MINI_ALU_BoothP_4,
                              L1_4_L2_3_G5_MINI_ALU_BoothP_3,
                              L1_4_L2_3_G5_MINI_ALU_BoothP_2,
                              L1_4_L2_3_G5_MINI_ALU_BoothP_1,
                              L1_4_L2_3_G5_MINI_ALU_BoothP_0}), .SelOperand (
                              nx3286), .Operation (
                              L1_4_L2_3_G5_MINI_ALU_BoothXORCheck), .AdderResult (
                              {L5FirstOperands_1__16,L5FirstOperands_1__15,
                              L5FirstOperands_1__14,L5FirstOperands_1__13,
                              L5FirstOperands_1__12,L5FirstOperands_1__11,
                              L5FirstOperands_1__10,L5FirstOperands_1__9,
                              L5FirstOperands_1__8,L5FirstOperands_1__7,
                              L5FirstOperands_1__6,L5FirstOperands_1__5,
                              L5FirstOperands_1__4,L5FirstOperands_1__3,
                              L5FirstOperands_1__2,L5FirstOperands_1__1,
                              L5FirstOperands_1__0}), .AdderBoothResult ({
                              \$dummy [823],
                              L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_15,
                              L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_14,
                              L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_13,
                              L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_12,
                              L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_11,
                              L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_10,
                              L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_9,
                              L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_8,
                              L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_7,
                              L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_6,
                              L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_5,
                              L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_4,
                              L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_3,
                              L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_2,
                              L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_1,
                              L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_0})) ;
    booth_unit_17 L1_4_L2_3_G5_MINI_ALU_BOOTH_UNIT (.CLK (CLK), .RST (RST), .Start (
                  Start), .Instr (Instr), .LoopingAndResultNotReady (nx3278), .Filter (
                  {FilterDin_4__3__7,FilterDin_4__3__6,FilterDin_4__3__5,
                  FilterDin_4__3__4,FilterDin_4__3__3,FilterDin_4__3__2,
                  FilterDin_4__3__1,FilterDin_4__3__0}), .Window ({
                  WindowDin_4__3__7,WindowDin_4__3__6,WindowDin_4__3__5,
                  WindowDin_4__3__4,WindowDin_4__3__3,WindowDin_4__3__2,
                  WindowDin_4__3__1,WindowDin_4__3__0}), .AdderBoothResult ({
                  L1FirstOperands_12__16,
                  L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_15,
                  L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_14,
                  L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_13,
                  L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_12,
                  L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_11,
                  L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_10,
                  L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_9,
                  L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_8,
                  L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_7,
                  L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_6,
                  L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_5,
                  L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_4,
                  L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_3,
                  L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_2,
                  L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_1,
                  L1_4_L2_3_G5_MINI_ALU_AdderBoothResult_0}), .BoothXORCheck (
                  L1_4_L2_3_G5_MINI_ALU_BoothXORCheck), .BoothResult ({
                  \$dummy [824],\$dummy [825],\$dummy [826],\$dummy [827],
                  \$dummy [828],\$dummy [829],\$dummy [830],\$dummy [831]}), .BoothAddingOperand (
                  {L1_4_L2_3_G5_MINI_ALU_BoothOperand_16,
                  L1_4_L2_3_G5_MINI_ALU_BoothOperand_15,
                  L1_4_L2_3_G5_MINI_ALU_BoothOperand_14,
                  L1_4_L2_3_G5_MINI_ALU_BoothOperand_13,
                  L1_4_L2_3_G5_MINI_ALU_BoothOperand_12,
                  L1_4_L2_3_G5_MINI_ALU_BoothOperand_11,
                  L1_4_L2_3_G5_MINI_ALU_BoothOperand_10,
                  L1_4_L2_3_G5_MINI_ALU_BoothOperand_9,\$dummy [832],
                  \$dummy [833],\$dummy [834],\$dummy [835],\$dummy [836],
                  \$dummy [837],\$dummy [838],\$dummy [839],\$dummy [840]}), .BoothP (
                  {L1_4_L2_3_G5_MINI_ALU_BoothP_16,
                  L1_4_L2_3_G5_MINI_ALU_BoothP_15,
                  L1_4_L2_3_G5_MINI_ALU_BoothP_14,
                  L1_4_L2_3_G5_MINI_ALU_BoothP_13,
                  L1_4_L2_3_G5_MINI_ALU_BoothP_12,
                  L1_4_L2_3_G5_MINI_ALU_BoothP_11,
                  L1_4_L2_3_G5_MINI_ALU_BoothP_10,L1_4_L2_3_G5_MINI_ALU_BoothP_9
                  ,L1_4_L2_3_G5_MINI_ALU_BoothP_8,L1_4_L2_3_G5_MINI_ALU_BoothP_7
                  ,L1_4_L2_3_G5_MINI_ALU_BoothP_6,L1_4_L2_3_G5_MINI_ALU_BoothP_5
                  ,L1_4_L2_3_G5_MINI_ALU_BoothP_4,L1_4_L2_3_G5_MINI_ALU_BoothP_3
                  ,L1_4_L2_3_G5_MINI_ALU_BoothP_2,L1_4_L2_3_G5_MINI_ALU_BoothP_1
                  ,L1_4_L2_3_G5_MINI_ALU_BoothP_0}), .LargeWindowShifted ({
                  \$dummy [841],\$dummy [842],\$dummy [843],\$dummy [844],
                  \$dummy [845],\$dummy [846],\$dummy [847],\$dummy [848],
                  \$dummy [849],\$dummy [850],\$dummy [851],\$dummy [852],
                  \$dummy [853],\$dummy [854],\$dummy [855],\$dummy [856],
                  \$dummy [857]})) ;
    booth_adder_17_unfolded17 L1_4_L2_4_G5_MINI_ALU_BOOTH_ADDER (.AdderFirstOperand (
                              {L5FirstOperands_1__16,L5FirstOperands_1__15,
                              L5FirstOperands_1__14,L5FirstOperands_1__13,
                              L5FirstOperands_1__12,L5FirstOperands_1__11,
                              L5FirstOperands_1__10,L5FirstOperands_1__9,
                              L5FirstOperands_1__8,L5FirstOperands_1__7,
                              L5FirstOperands_1__6,L5FirstOperands_1__5,
                              L5FirstOperands_1__4,L5FirstOperands_1__3,
                              L5FirstOperands_1__2,L5FirstOperands_1__1,
                              L5FirstOperands_1__0}), .AdderSecondOperand ({
                              L1FirstOperands_12__16,
                              L1_4_L2_4_G5_MINI_ALU_OperationResult_15,
                              L1_4_L2_4_G5_MINI_ALU_OperationResult_14,
                              L1_4_L2_4_G5_MINI_ALU_OperationResult_13,
                              L1_4_L2_4_G5_MINI_ALU_OperationResult_12,
                              L1_4_L2_4_G5_MINI_ALU_OperationResult_11,
                              L1_4_L2_4_G5_MINI_ALU_OperationResult_10,
                              L1_4_L2_4_G5_MINI_ALU_OperationResult_9,
                              L1_4_L2_4_G5_MINI_ALU_OperationResult_8,
                              L1_4_L2_4_G5_MINI_ALU_OperationResult_7,
                              L1_4_L2_4_G5_MINI_ALU_OperationResult_6,
                              L1_4_L2_4_G5_MINI_ALU_OperationResult_5,
                              L1_4_L2_4_G5_MINI_ALU_OperationResult_4,
                              L1_4_L2_4_G5_MINI_ALU_OperationResult_3,
                              L1_4_L2_4_G5_MINI_ALU_OperationResult_2,
                              L1_4_L2_4_G5_MINI_ALU_OperationResult_1,
                              L1_4_L2_4_G5_MINI_ALU_OperationResult_0}), .BoothOperand (
                              {L1_4_L2_4_G5_MINI_ALU_BoothOperand_16,
                              L1_4_L2_4_G5_MINI_ALU_BoothOperand_15,
                              L1_4_L2_4_G5_MINI_ALU_BoothOperand_14,
                              L1_4_L2_4_G5_MINI_ALU_BoothOperand_13,
                              L1_4_L2_4_G5_MINI_ALU_BoothOperand_12,
                              L1_4_L2_4_G5_MINI_ALU_BoothOperand_11,
                              L1_4_L2_4_G5_MINI_ALU_BoothOperand_10,
                              L1_4_L2_4_G5_MINI_ALU_BoothOperand_9,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16,L1FirstOperands_12__16,
                              L1FirstOperands_12__16}), .BoothP ({
                              L1_4_L2_4_G5_MINI_ALU_BoothP_16,
                              L1_4_L2_4_G5_MINI_ALU_BoothP_15,
                              L1_4_L2_4_G5_MINI_ALU_BoothP_14,
                              L1_4_L2_4_G5_MINI_ALU_BoothP_13,
                              L1_4_L2_4_G5_MINI_ALU_BoothP_12,
                              L1_4_L2_4_G5_MINI_ALU_BoothP_11,
                              L1_4_L2_4_G5_MINI_ALU_BoothP_10,
                              L1_4_L2_4_G5_MINI_ALU_BoothP_9,
                              L1_4_L2_4_G5_MINI_ALU_BoothP_8,
                              L1_4_L2_4_G5_MINI_ALU_BoothP_7,
                              L1_4_L2_4_G5_MINI_ALU_BoothP_6,
                              L1_4_L2_4_G5_MINI_ALU_BoothP_5,
                              L1_4_L2_4_G5_MINI_ALU_BoothP_4,
                              L1_4_L2_4_G5_MINI_ALU_BoothP_3,
                              L1_4_L2_4_G5_MINI_ALU_BoothP_2,
                              L1_4_L2_4_G5_MINI_ALU_BoothP_1,
                              L1_4_L2_4_G5_MINI_ALU_BoothP_0}), .SelOperand (
                              nx3286), .Operation (
                              L1_4_L2_4_G5_MINI_ALU_BoothXORCheck), .AdderResult (
                              {\$dummy [858],\$dummy [859],\$dummy [860],
                              \$dummy [861],\$dummy [862],\$dummy [863],
                              \$dummy [864],\$dummy [865],\$dummy [866],
                              L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_7,
                              L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_6,
                              L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_5,
                              L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_4,
                              L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_3,
                              L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_2,
                              L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_1,
                              L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_0}), .AdderBoothResult (
                              {\$dummy [867],
                              L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_15,
                              L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_14,
                              L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_13,
                              L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_12,
                              L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_11,
                              L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_10,
                              L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_9,
                              L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_8,
                              L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_7,
                              L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_6,
                              L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_5,
                              L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_4,
                              L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_3,
                              L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_2,
                              L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_1,
                              L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_0})) ;
    booth_unit_17 L1_4_L2_4_G5_MINI_ALU_BOOTH_UNIT (.CLK (CLK), .RST (RST), .Start (
                  Start), .Instr (Instr), .LoopingAndResultNotReady (nx3278), .Filter (
                  {FilterDin_4__4__7,FilterDin_4__4__6,FilterDin_4__4__5,
                  FilterDin_4__4__4,FilterDin_4__4__3,FilterDin_4__4__2,
                  FilterDin_4__4__1,FilterDin_4__4__0}), .Window ({
                  WindowDin_4__4__7,WindowDin_4__4__6,WindowDin_4__4__5,
                  WindowDin_4__4__4,WindowDin_4__4__3,WindowDin_4__4__2,
                  WindowDin_4__4__1,WindowDin_4__4__0}), .AdderBoothResult ({
                  L1FirstOperands_12__16,
                  L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_15,
                  L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_14,
                  L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_13,
                  L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_12,
                  L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_11,
                  L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_10,
                  L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_9,
                  L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_8,
                  L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_7,
                  L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_6,
                  L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_5,
                  L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_4,
                  L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_3,
                  L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_2,
                  L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_1,
                  L1_4_L2_4_G5_MINI_ALU_AdderBoothResult_0}), .BoothXORCheck (
                  L1_4_L2_4_G5_MINI_ALU_BoothXORCheck), .BoothResult ({
                  \$dummy [868],\$dummy [869],\$dummy [870],\$dummy [871],
                  \$dummy [872],\$dummy [873],\$dummy [874],\$dummy [875]}), .BoothAddingOperand (
                  {L1_4_L2_4_G5_MINI_ALU_BoothOperand_16,
                  L1_4_L2_4_G5_MINI_ALU_BoothOperand_15,
                  L1_4_L2_4_G5_MINI_ALU_BoothOperand_14,
                  L1_4_L2_4_G5_MINI_ALU_BoothOperand_13,
                  L1_4_L2_4_G5_MINI_ALU_BoothOperand_12,
                  L1_4_L2_4_G5_MINI_ALU_BoothOperand_11,
                  L1_4_L2_4_G5_MINI_ALU_BoothOperand_10,
                  L1_4_L2_4_G5_MINI_ALU_BoothOperand_9,\$dummy [876],
                  \$dummy [877],\$dummy [878],\$dummy [879],\$dummy [880],
                  \$dummy [881],\$dummy [882],\$dummy [883],\$dummy [884]}), .BoothP (
                  {L1_4_L2_4_G5_MINI_ALU_BoothP_16,
                  L1_4_L2_4_G5_MINI_ALU_BoothP_15,
                  L1_4_L2_4_G5_MINI_ALU_BoothP_14,
                  L1_4_L2_4_G5_MINI_ALU_BoothP_13,
                  L1_4_L2_4_G5_MINI_ALU_BoothP_12,
                  L1_4_L2_4_G5_MINI_ALU_BoothP_11,
                  L1_4_L2_4_G5_MINI_ALU_BoothP_10,L1_4_L2_4_G5_MINI_ALU_BoothP_9
                  ,L1_4_L2_4_G5_MINI_ALU_BoothP_8,L1_4_L2_4_G5_MINI_ALU_BoothP_7
                  ,L1_4_L2_4_G5_MINI_ALU_BoothP_6,L1_4_L2_4_G5_MINI_ALU_BoothP_5
                  ,L1_4_L2_4_G5_MINI_ALU_BoothP_4,L1_4_L2_4_G5_MINI_ALU_BoothP_3
                  ,L1_4_L2_4_G5_MINI_ALU_BoothP_2,L1_4_L2_4_G5_MINI_ALU_BoothP_1
                  ,L1_4_L2_4_G5_MINI_ALU_BoothP_0}), .LargeWindowShifted ({
                  \$dummy [885],\$dummy [886],\$dummy [887],\$dummy [888],
                  \$dummy [889],\$dummy [890],\$dummy [891],\$dummy [892],
                  \$dummy [893],\$dummy [894],\$dummy [895],\$dummy [896],
                  \$dummy [897],\$dummy [898],\$dummy [899],\$dummy [900],
                  \$dummy [901]})) ;
    nor02ii ix2852 (.Y (NOT__145383), .A0 (Instr), .A1 (nx2853)) ;
    nand03 ix2854 (.Y (nx2853), .A0 (CounterOut_0), .A1 (CounterOut_3), .A2 (
           nx2873)) ;
    dffr reg_CounterOut_0 (.Q (CounterOut_0), .QB (NOT_CounterOut_0), .D (
         NOT_CounterOut_0), .CLK (nx1032), .R (nx1036)) ;
    or02 ix1037 (.Y (nx1036), .A0 (Start), .A1 (RST)) ;
    dffr reg_CounterOut_3 (.Q (CounterOut_3), .QB (\$dummy [902]), .D (nx1066), 
         .CLK (nx1032), .R (nx1036)) ;
    xnor2 ix1067 (.Y (nx1066), .A0 (CounterOut_3), .A1 (nx2865)) ;
    nand03 ix2866 (.Y (nx2865), .A0 (CounterOut_2), .A1 (CounterOut_1), .A2 (
           CounterOut_0)) ;
    dffr reg_CounterOut_2 (.Q (CounterOut_2), .QB (\$dummy [903]), .D (nx1058), 
         .CLK (nx1032), .R (nx1036)) ;
    xnor2 ix1059 (.Y (nx1058), .A0 (CounterOut_2), .A1 (nx2869)) ;
    dffr reg_CounterOut_1 (.Q (CounterOut_1), .QB (nx2873), .D (nx1046), .CLK (
         nx1032), .R (nx1036)) ;
    fake_gnd ix2302 (.Y (L1FirstOperands_12__16)) ;
    mux21_ni ix109 (.Y (L1_4_L2_4_G5_MINI_ALU_OperationResult_0), .A0 (
             L1_4_L2_4_G5_MINI_ALU_BoothP_1), .A1 (WindowDin_4__4__0), .S0 (
             Instr)) ;
    mux21_ni ix117 (.Y (L1_4_L2_4_G5_MINI_ALU_OperationResult_1), .A0 (
             L1_4_L2_4_G5_MINI_ALU_BoothP_2), .A1 (WindowDin_4__4__1), .S0 (
             Instr)) ;
    mux21_ni ix125 (.Y (L1_4_L2_4_G5_MINI_ALU_OperationResult_2), .A0 (
             L1_4_L2_4_G5_MINI_ALU_BoothP_3), .A1 (WindowDin_4__4__2), .S0 (
             Instr)) ;
    mux21_ni ix133 (.Y (L1_4_L2_4_G5_MINI_ALU_OperationResult_3), .A0 (
             L1_4_L2_4_G5_MINI_ALU_BoothP_4), .A1 (WindowDin_4__4__3), .S0 (
             Instr)) ;
    mux21_ni ix141 (.Y (L1_4_L2_4_G5_MINI_ALU_OperationResult_4), .A0 (
             L1_4_L2_4_G5_MINI_ALU_BoothP_5), .A1 (WindowDin_4__4__4), .S0 (
             Instr)) ;
    mux21_ni ix149 (.Y (L1_4_L2_4_G5_MINI_ALU_OperationResult_5), .A0 (
             L1_4_L2_4_G5_MINI_ALU_BoothP_6), .A1 (WindowDin_4__4__5), .S0 (
             Instr)) ;
    mux21_ni ix157 (.Y (L1_4_L2_4_G5_MINI_ALU_OperationResult_6), .A0 (
             L1_4_L2_4_G5_MINI_ALU_BoothP_7), .A1 (WindowDin_4__4__6), .S0 (
             Instr)) ;
    mux21_ni ix165 (.Y (L1_4_L2_4_G5_MINI_ALU_OperationResult_7), .A0 (
             L1_4_L2_4_G5_MINI_ALU_BoothP_8), .A1 (WindowDin_4__4__7), .S0 (
             Instr)) ;
    nor02ii ix73 (.Y (L1_4_L2_4_G5_MINI_ALU_OperationResult_8), .A0 (Instr), .A1 (
            L1_4_L2_4_G5_MINI_ALU_BoothP_9)) ;
    nor02ii ix77 (.Y (L1_4_L2_4_G5_MINI_ALU_OperationResult_9), .A0 (Instr), .A1 (
            L1_4_L2_4_G5_MINI_ALU_BoothP_10)) ;
    nor02ii ix81 (.Y (L1_4_L2_4_G5_MINI_ALU_OperationResult_10), .A0 (Instr), .A1 (
            L1_4_L2_4_G5_MINI_ALU_BoothP_11)) ;
    nor02ii ix85 (.Y (L1_4_L2_4_G5_MINI_ALU_OperationResult_11), .A0 (Instr), .A1 (
            L1_4_L2_4_G5_MINI_ALU_BoothP_12)) ;
    nor02ii ix89 (.Y (L1_4_L2_4_G5_MINI_ALU_OperationResult_12), .A0 (Instr), .A1 (
            L1_4_L2_4_G5_MINI_ALU_BoothP_13)) ;
    nor02ii ix93 (.Y (L1_4_L2_4_G5_MINI_ALU_OperationResult_13), .A0 (Instr), .A1 (
            L1_4_L2_4_G5_MINI_ALU_BoothP_14)) ;
    nor02ii ix97 (.Y (L1_4_L2_4_G5_MINI_ALU_OperationResult_14), .A0 (Instr), .A1 (
            L1_4_L2_4_G5_MINI_ALU_BoothP_15)) ;
    nor02ii ix101 (.Y (L1_4_L2_4_G5_MINI_ALU_OperationResult_15), .A0 (Instr), .A1 (
            L1_4_L2_4_G5_MINI_ALU_BoothP_16)) ;
    mux21_ni ix1121 (.Y (L1_2_L2_1_G1_MINI_ALU_OperationResult_0), .A0 (
             L1_2_L2_1_G1_MINI_ALU_BoothP_1), .A1 (WindowDin_2__1__0), .S0 (
             Instr)) ;
    mux21_ni ix1129 (.Y (L1_2_L2_1_G1_MINI_ALU_OperationResult_1), .A0 (
             L1_2_L2_1_G1_MINI_ALU_BoothP_2), .A1 (WindowDin_2__1__1), .S0 (
             Instr)) ;
    mux21_ni ix1137 (.Y (L1_2_L2_1_G1_MINI_ALU_OperationResult_2), .A0 (
             L1_2_L2_1_G1_MINI_ALU_BoothP_3), .A1 (WindowDin_2__1__2), .S0 (
             Instr)) ;
    mux21_ni ix1145 (.Y (L1_2_L2_1_G1_MINI_ALU_OperationResult_3), .A0 (
             L1_2_L2_1_G1_MINI_ALU_BoothP_4), .A1 (WindowDin_2__1__3), .S0 (
             Instr)) ;
    mux21_ni ix1153 (.Y (L1_2_L2_1_G1_MINI_ALU_OperationResult_4), .A0 (
             L1_2_L2_1_G1_MINI_ALU_BoothP_5), .A1 (WindowDin_2__1__4), .S0 (
             Instr)) ;
    mux21_ni ix1161 (.Y (L1_2_L2_1_G1_MINI_ALU_OperationResult_5), .A0 (
             L1_2_L2_1_G1_MINI_ALU_BoothP_6), .A1 (WindowDin_2__1__5), .S0 (
             Instr)) ;
    mux21_ni ix1169 (.Y (L1_2_L2_1_G1_MINI_ALU_OperationResult_6), .A0 (
             L1_2_L2_1_G1_MINI_ALU_BoothP_7), .A1 (WindowDin_2__1__6), .S0 (
             Instr)) ;
    mux21_ni ix1177 (.Y (L1_2_L2_1_G1_MINI_ALU_OperationResult_7), .A0 (
             L1_2_L2_1_G1_MINI_ALU_BoothP_8), .A1 (WindowDin_2__1__7), .S0 (
             Instr)) ;
    nor02ii ix1085 (.Y (L1_2_L2_1_G1_MINI_ALU_OperationResult_8), .A0 (Instr), .A1 (
            L1_2_L2_1_G1_MINI_ALU_BoothP_9)) ;
    nor02ii ix1089 (.Y (L1_2_L2_1_G1_MINI_ALU_OperationResult_9), .A0 (Instr), .A1 (
            L1_2_L2_1_G1_MINI_ALU_BoothP_10)) ;
    nor02ii ix1093 (.Y (L1_2_L2_1_G1_MINI_ALU_OperationResult_10), .A0 (Instr), 
            .A1 (L1_2_L2_1_G1_MINI_ALU_BoothP_11)) ;
    nor02ii ix1097 (.Y (L1_2_L2_1_G1_MINI_ALU_OperationResult_11), .A0 (Instr), 
            .A1 (L1_2_L2_1_G1_MINI_ALU_BoothP_12)) ;
    nor02ii ix1101 (.Y (L1_2_L2_1_G1_MINI_ALU_OperationResult_12), .A0 (Instr), 
            .A1 (L1_2_L2_1_G1_MINI_ALU_BoothP_13)) ;
    nor02ii ix1105 (.Y (L1_2_L2_1_G1_MINI_ALU_OperationResult_13), .A0 (Instr), 
            .A1 (L1_2_L2_1_G1_MINI_ALU_BoothP_14)) ;
    nor02ii ix1109 (.Y (L1_2_L2_1_G1_MINI_ALU_OperationResult_14), .A0 (Instr), 
            .A1 (L1_2_L2_1_G1_MINI_ALU_BoothP_15)) ;
    nor02ii ix1113 (.Y (L1_2_L2_1_G1_MINI_ALU_OperationResult_15), .A0 (Instr), 
            .A1 (L1_2_L2_1_G1_MINI_ALU_BoothP_16)) ;
    mux21_ni ix1217 (.Y (L1_2_L2_0_G1_MINI_ALU_OperationResult_0), .A0 (
             L1_2_L2_0_G1_MINI_ALU_BoothP_1), .A1 (WindowDin_2__0__0), .S0 (
             Instr)) ;
    mux21_ni ix1225 (.Y (L1_2_L2_0_G1_MINI_ALU_OperationResult_1), .A0 (
             L1_2_L2_0_G1_MINI_ALU_BoothP_2), .A1 (WindowDin_2__0__1), .S0 (
             Instr)) ;
    mux21_ni ix1233 (.Y (L1_2_L2_0_G1_MINI_ALU_OperationResult_2), .A0 (
             L1_2_L2_0_G1_MINI_ALU_BoothP_3), .A1 (WindowDin_2__0__2), .S0 (
             Instr)) ;
    mux21_ni ix1241 (.Y (L1_2_L2_0_G1_MINI_ALU_OperationResult_3), .A0 (
             L1_2_L2_0_G1_MINI_ALU_BoothP_4), .A1 (WindowDin_2__0__3), .S0 (
             Instr)) ;
    mux21_ni ix1249 (.Y (L1_2_L2_0_G1_MINI_ALU_OperationResult_4), .A0 (
             L1_2_L2_0_G1_MINI_ALU_BoothP_5), .A1 (WindowDin_2__0__4), .S0 (
             Instr)) ;
    mux21_ni ix1257 (.Y (L1_2_L2_0_G1_MINI_ALU_OperationResult_5), .A0 (
             L1_2_L2_0_G1_MINI_ALU_BoothP_6), .A1 (WindowDin_2__0__5), .S0 (
             Instr)) ;
    mux21_ni ix1265 (.Y (L1_2_L2_0_G1_MINI_ALU_OperationResult_6), .A0 (
             L1_2_L2_0_G1_MINI_ALU_BoothP_7), .A1 (WindowDin_2__0__6), .S0 (
             Instr)) ;
    mux21_ni ix1273 (.Y (L1_2_L2_0_G1_MINI_ALU_OperationResult_7), .A0 (
             L1_2_L2_0_G1_MINI_ALU_BoothP_8), .A1 (WindowDin_2__0__7), .S0 (
             Instr)) ;
    nor02ii ix1181 (.Y (L1_2_L2_0_G1_MINI_ALU_OperationResult_8), .A0 (Instr), .A1 (
            L1_2_L2_0_G1_MINI_ALU_BoothP_9)) ;
    nor02ii ix1185 (.Y (L1_2_L2_0_G1_MINI_ALU_OperationResult_9), .A0 (Instr), .A1 (
            L1_2_L2_0_G1_MINI_ALU_BoothP_10)) ;
    nor02ii ix1189 (.Y (L1_2_L2_0_G1_MINI_ALU_OperationResult_10), .A0 (Instr), 
            .A1 (L1_2_L2_0_G1_MINI_ALU_BoothP_11)) ;
    nor02ii ix1193 (.Y (L1_2_L2_0_G1_MINI_ALU_OperationResult_11), .A0 (Instr), 
            .A1 (L1_2_L2_0_G1_MINI_ALU_BoothP_12)) ;
    nor02ii ix1197 (.Y (L1_2_L2_0_G1_MINI_ALU_OperationResult_12), .A0 (Instr), 
            .A1 (L1_2_L2_0_G1_MINI_ALU_BoothP_13)) ;
    nor02ii ix1201 (.Y (L1_2_L2_0_G1_MINI_ALU_OperationResult_13), .A0 (Instr), 
            .A1 (L1_2_L2_0_G1_MINI_ALU_BoothP_14)) ;
    nor02ii ix1205 (.Y (L1_2_L2_0_G1_MINI_ALU_OperationResult_14), .A0 (Instr), 
            .A1 (L1_2_L2_0_G1_MINI_ALU_BoothP_15)) ;
    nor02ii ix1209 (.Y (L1_2_L2_0_G1_MINI_ALU_OperationResult_15), .A0 (Instr), 
            .A1 (L1_2_L2_0_G1_MINI_ALU_BoothP_16)) ;
    mux21_ni ix1313 (.Y (L1_1_L2_4_G1_MINI_ALU_OperationResult_0), .A0 (
             L1_1_L2_4_G1_MINI_ALU_BoothP_1), .A1 (WindowDin_1__4__0), .S0 (
             Instr)) ;
    mux21_ni ix1321 (.Y (L1_1_L2_4_G1_MINI_ALU_OperationResult_1), .A0 (
             L1_1_L2_4_G1_MINI_ALU_BoothP_2), .A1 (WindowDin_1__4__1), .S0 (
             Instr)) ;
    mux21_ni ix1329 (.Y (L1_1_L2_4_G1_MINI_ALU_OperationResult_2), .A0 (
             L1_1_L2_4_G1_MINI_ALU_BoothP_3), .A1 (WindowDin_1__4__2), .S0 (
             Instr)) ;
    mux21_ni ix1337 (.Y (L1_1_L2_4_G1_MINI_ALU_OperationResult_3), .A0 (
             L1_1_L2_4_G1_MINI_ALU_BoothP_4), .A1 (WindowDin_1__4__3), .S0 (
             Instr)) ;
    mux21_ni ix1345 (.Y (L1_1_L2_4_G1_MINI_ALU_OperationResult_4), .A0 (
             L1_1_L2_4_G1_MINI_ALU_BoothP_5), .A1 (WindowDin_1__4__4), .S0 (
             Instr)) ;
    mux21_ni ix1353 (.Y (L1_1_L2_4_G1_MINI_ALU_OperationResult_5), .A0 (
             L1_1_L2_4_G1_MINI_ALU_BoothP_6), .A1 (WindowDin_1__4__5), .S0 (
             Instr)) ;
    mux21_ni ix1361 (.Y (L1_1_L2_4_G1_MINI_ALU_OperationResult_6), .A0 (
             L1_1_L2_4_G1_MINI_ALU_BoothP_7), .A1 (WindowDin_1__4__6), .S0 (
             Instr)) ;
    mux21_ni ix1369 (.Y (L1_1_L2_4_G1_MINI_ALU_OperationResult_7), .A0 (
             L1_1_L2_4_G1_MINI_ALU_BoothP_8), .A1 (WindowDin_1__4__7), .S0 (
             Instr)) ;
    nor02ii ix1277 (.Y (L1_1_L2_4_G1_MINI_ALU_OperationResult_8), .A0 (Instr), .A1 (
            L1_1_L2_4_G1_MINI_ALU_BoothP_9)) ;
    nor02ii ix1281 (.Y (L1_1_L2_4_G1_MINI_ALU_OperationResult_9), .A0 (Instr), .A1 (
            L1_1_L2_4_G1_MINI_ALU_BoothP_10)) ;
    nor02ii ix1285 (.Y (L1_1_L2_4_G1_MINI_ALU_OperationResult_10), .A0 (Instr), 
            .A1 (L1_1_L2_4_G1_MINI_ALU_BoothP_11)) ;
    nor02ii ix1289 (.Y (L1_1_L2_4_G1_MINI_ALU_OperationResult_11), .A0 (Instr), 
            .A1 (L1_1_L2_4_G1_MINI_ALU_BoothP_12)) ;
    nor02ii ix1293 (.Y (L1_1_L2_4_G1_MINI_ALU_OperationResult_12), .A0 (Instr), 
            .A1 (L1_1_L2_4_G1_MINI_ALU_BoothP_13)) ;
    nor02ii ix1297 (.Y (L1_1_L2_4_G1_MINI_ALU_OperationResult_13), .A0 (Instr), 
            .A1 (L1_1_L2_4_G1_MINI_ALU_BoothP_14)) ;
    nor02ii ix1301 (.Y (L1_1_L2_4_G1_MINI_ALU_OperationResult_14), .A0 (Instr), 
            .A1 (L1_1_L2_4_G1_MINI_ALU_BoothP_15)) ;
    nor02ii ix1305 (.Y (L1_1_L2_4_G1_MINI_ALU_OperationResult_15), .A0 (Instr), 
            .A1 (L1_1_L2_4_G1_MINI_ALU_BoothP_16)) ;
    mux21_ni ix1409 (.Y (L1_1_L2_3_G1_MINI_ALU_OperationResult_0), .A0 (
             L1_1_L2_3_G1_MINI_ALU_BoothP_1), .A1 (WindowDin_1__3__0), .S0 (
             Instr)) ;
    mux21_ni ix1417 (.Y (L1_1_L2_3_G1_MINI_ALU_OperationResult_1), .A0 (
             L1_1_L2_3_G1_MINI_ALU_BoothP_2), .A1 (WindowDin_1__3__1), .S0 (
             Instr)) ;
    mux21_ni ix1425 (.Y (L1_1_L2_3_G1_MINI_ALU_OperationResult_2), .A0 (
             L1_1_L2_3_G1_MINI_ALU_BoothP_3), .A1 (WindowDin_1__3__2), .S0 (
             Instr)) ;
    mux21_ni ix1433 (.Y (L1_1_L2_3_G1_MINI_ALU_OperationResult_3), .A0 (
             L1_1_L2_3_G1_MINI_ALU_BoothP_4), .A1 (WindowDin_1__3__3), .S0 (
             Instr)) ;
    mux21_ni ix1441 (.Y (L1_1_L2_3_G1_MINI_ALU_OperationResult_4), .A0 (
             L1_1_L2_3_G1_MINI_ALU_BoothP_5), .A1 (WindowDin_1__3__4), .S0 (
             Instr)) ;
    mux21_ni ix1449 (.Y (L1_1_L2_3_G1_MINI_ALU_OperationResult_5), .A0 (
             L1_1_L2_3_G1_MINI_ALU_BoothP_6), .A1 (WindowDin_1__3__5), .S0 (
             Instr)) ;
    mux21_ni ix1457 (.Y (L1_1_L2_3_G1_MINI_ALU_OperationResult_6), .A0 (
             L1_1_L2_3_G1_MINI_ALU_BoothP_7), .A1 (WindowDin_1__3__6), .S0 (
             Instr)) ;
    mux21_ni ix1465 (.Y (L1_1_L2_3_G1_MINI_ALU_OperationResult_7), .A0 (
             L1_1_L2_3_G1_MINI_ALU_BoothP_8), .A1 (WindowDin_1__3__7), .S0 (
             Instr)) ;
    nor02ii ix1373 (.Y (L1_1_L2_3_G1_MINI_ALU_OperationResult_8), .A0 (Instr), .A1 (
            L1_1_L2_3_G1_MINI_ALU_BoothP_9)) ;
    nor02ii ix1377 (.Y (L1_1_L2_3_G1_MINI_ALU_OperationResult_9), .A0 (Instr), .A1 (
            L1_1_L2_3_G1_MINI_ALU_BoothP_10)) ;
    nor02ii ix1381 (.Y (L1_1_L2_3_G1_MINI_ALU_OperationResult_10), .A0 (Instr), 
            .A1 (L1_1_L2_3_G1_MINI_ALU_BoothP_11)) ;
    nor02ii ix1385 (.Y (L1_1_L2_3_G1_MINI_ALU_OperationResult_11), .A0 (Instr), 
            .A1 (L1_1_L2_3_G1_MINI_ALU_BoothP_12)) ;
    nor02ii ix1389 (.Y (L1_1_L2_3_G1_MINI_ALU_OperationResult_12), .A0 (Instr), 
            .A1 (L1_1_L2_3_G1_MINI_ALU_BoothP_13)) ;
    nor02ii ix1393 (.Y (L1_1_L2_3_G1_MINI_ALU_OperationResult_13), .A0 (Instr), 
            .A1 (L1_1_L2_3_G1_MINI_ALU_BoothP_14)) ;
    nor02ii ix1397 (.Y (L1_1_L2_3_G1_MINI_ALU_OperationResult_14), .A0 (Instr), 
            .A1 (L1_1_L2_3_G1_MINI_ALU_BoothP_15)) ;
    nor02ii ix1401 (.Y (L1_1_L2_3_G1_MINI_ALU_OperationResult_15), .A0 (Instr), 
            .A1 (L1_1_L2_3_G1_MINI_ALU_BoothP_16)) ;
    mux21_ni ix1505 (.Y (L1_1_L2_2_G1_MINI_ALU_OperationResult_0), .A0 (
             L1_1_L2_2_G1_MINI_ALU_BoothP_1), .A1 (WindowDin_1__2__0), .S0 (
             Instr)) ;
    mux21_ni ix1513 (.Y (L1_1_L2_2_G1_MINI_ALU_OperationResult_1), .A0 (
             L1_1_L2_2_G1_MINI_ALU_BoothP_2), .A1 (WindowDin_1__2__1), .S0 (
             Instr)) ;
    mux21_ni ix1521 (.Y (L1_1_L2_2_G1_MINI_ALU_OperationResult_2), .A0 (
             L1_1_L2_2_G1_MINI_ALU_BoothP_3), .A1 (WindowDin_1__2__2), .S0 (
             Instr)) ;
    mux21_ni ix1529 (.Y (L1_1_L2_2_G1_MINI_ALU_OperationResult_3), .A0 (
             L1_1_L2_2_G1_MINI_ALU_BoothP_4), .A1 (WindowDin_1__2__3), .S0 (
             Instr)) ;
    mux21_ni ix1537 (.Y (L1_1_L2_2_G1_MINI_ALU_OperationResult_4), .A0 (
             L1_1_L2_2_G1_MINI_ALU_BoothP_5), .A1 (WindowDin_1__2__4), .S0 (
             Instr)) ;
    mux21_ni ix1545 (.Y (L1_1_L2_2_G1_MINI_ALU_OperationResult_5), .A0 (
             L1_1_L2_2_G1_MINI_ALU_BoothP_6), .A1 (WindowDin_1__2__5), .S0 (
             Instr)) ;
    mux21_ni ix1553 (.Y (L1_1_L2_2_G1_MINI_ALU_OperationResult_6), .A0 (
             L1_1_L2_2_G1_MINI_ALU_BoothP_7), .A1 (WindowDin_1__2__6), .S0 (
             Instr)) ;
    mux21_ni ix1561 (.Y (L1_1_L2_2_G1_MINI_ALU_OperationResult_7), .A0 (
             L1_1_L2_2_G1_MINI_ALU_BoothP_8), .A1 (WindowDin_1__2__7), .S0 (
             Instr)) ;
    nor02ii ix1469 (.Y (L1_1_L2_2_G1_MINI_ALU_OperationResult_8), .A0 (Instr), .A1 (
            L1_1_L2_2_G1_MINI_ALU_BoothP_9)) ;
    nor02ii ix1473 (.Y (L1_1_L2_2_G1_MINI_ALU_OperationResult_9), .A0 (Instr), .A1 (
            L1_1_L2_2_G1_MINI_ALU_BoothP_10)) ;
    nor02ii ix1477 (.Y (L1_1_L2_2_G1_MINI_ALU_OperationResult_10), .A0 (Instr), 
            .A1 (L1_1_L2_2_G1_MINI_ALU_BoothP_11)) ;
    nor02ii ix1481 (.Y (L1_1_L2_2_G1_MINI_ALU_OperationResult_11), .A0 (Instr), 
            .A1 (L1_1_L2_2_G1_MINI_ALU_BoothP_12)) ;
    nor02ii ix1485 (.Y (L1_1_L2_2_G1_MINI_ALU_OperationResult_12), .A0 (Instr), 
            .A1 (L1_1_L2_2_G1_MINI_ALU_BoothP_13)) ;
    nor02ii ix1489 (.Y (L1_1_L2_2_G1_MINI_ALU_OperationResult_13), .A0 (Instr), 
            .A1 (L1_1_L2_2_G1_MINI_ALU_BoothP_14)) ;
    nor02ii ix1493 (.Y (L1_1_L2_2_G1_MINI_ALU_OperationResult_14), .A0 (Instr), 
            .A1 (L1_1_L2_2_G1_MINI_ALU_BoothP_15)) ;
    nor02ii ix1497 (.Y (L1_1_L2_2_G1_MINI_ALU_OperationResult_15), .A0 (Instr), 
            .A1 (L1_1_L2_2_G1_MINI_ALU_BoothP_16)) ;
    mux21_ni ix1601 (.Y (L1_1_L2_1_G1_MINI_ALU_OperationResult_0), .A0 (
             L1_1_L2_1_G1_MINI_ALU_BoothP_1), .A1 (WindowDin_1__1__0), .S0 (
             Instr)) ;
    mux21_ni ix1609 (.Y (L1_1_L2_1_G1_MINI_ALU_OperationResult_1), .A0 (
             L1_1_L2_1_G1_MINI_ALU_BoothP_2), .A1 (WindowDin_1__1__1), .S0 (
             Instr)) ;
    mux21_ni ix1617 (.Y (L1_1_L2_1_G1_MINI_ALU_OperationResult_2), .A0 (
             L1_1_L2_1_G1_MINI_ALU_BoothP_3), .A1 (WindowDin_1__1__2), .S0 (
             Instr)) ;
    mux21_ni ix1625 (.Y (L1_1_L2_1_G1_MINI_ALU_OperationResult_3), .A0 (
             L1_1_L2_1_G1_MINI_ALU_BoothP_4), .A1 (WindowDin_1__1__3), .S0 (
             Instr)) ;
    mux21_ni ix1633 (.Y (L1_1_L2_1_G1_MINI_ALU_OperationResult_4), .A0 (
             L1_1_L2_1_G1_MINI_ALU_BoothP_5), .A1 (WindowDin_1__1__4), .S0 (
             Instr)) ;
    mux21_ni ix1641 (.Y (L1_1_L2_1_G1_MINI_ALU_OperationResult_5), .A0 (
             L1_1_L2_1_G1_MINI_ALU_BoothP_6), .A1 (WindowDin_1__1__5), .S0 (
             Instr)) ;
    mux21_ni ix1649 (.Y (L1_1_L2_1_G1_MINI_ALU_OperationResult_6), .A0 (
             L1_1_L2_1_G1_MINI_ALU_BoothP_7), .A1 (WindowDin_1__1__6), .S0 (
             Instr)) ;
    mux21_ni ix1657 (.Y (L1_1_L2_1_G1_MINI_ALU_OperationResult_7), .A0 (
             L1_1_L2_1_G1_MINI_ALU_BoothP_8), .A1 (WindowDin_1__1__7), .S0 (
             Instr)) ;
    nor02ii ix1565 (.Y (L1_1_L2_1_G1_MINI_ALU_OperationResult_8), .A0 (Instr), .A1 (
            L1_1_L2_1_G1_MINI_ALU_BoothP_9)) ;
    nor02ii ix1569 (.Y (L1_1_L2_1_G1_MINI_ALU_OperationResult_9), .A0 (Instr), .A1 (
            L1_1_L2_1_G1_MINI_ALU_BoothP_10)) ;
    nor02ii ix1573 (.Y (L1_1_L2_1_G1_MINI_ALU_OperationResult_10), .A0 (Instr), 
            .A1 (L1_1_L2_1_G1_MINI_ALU_BoothP_11)) ;
    nor02ii ix1577 (.Y (L1_1_L2_1_G1_MINI_ALU_OperationResult_11), .A0 (Instr), 
            .A1 (L1_1_L2_1_G1_MINI_ALU_BoothP_12)) ;
    nor02ii ix1581 (.Y (L1_1_L2_1_G1_MINI_ALU_OperationResult_12), .A0 (Instr), 
            .A1 (L1_1_L2_1_G1_MINI_ALU_BoothP_13)) ;
    nor02ii ix1585 (.Y (L1_1_L2_1_G1_MINI_ALU_OperationResult_13), .A0 (Instr), 
            .A1 (L1_1_L2_1_G1_MINI_ALU_BoothP_14)) ;
    nor02ii ix1589 (.Y (L1_1_L2_1_G1_MINI_ALU_OperationResult_14), .A0 (Instr), 
            .A1 (L1_1_L2_1_G1_MINI_ALU_BoothP_15)) ;
    nor02ii ix1593 (.Y (L1_1_L2_1_G1_MINI_ALU_OperationResult_15), .A0 (Instr), 
            .A1 (L1_1_L2_1_G1_MINI_ALU_BoothP_16)) ;
    mux21_ni ix1697 (.Y (L1_1_L2_0_G1_MINI_ALU_OperationResult_0), .A0 (
             L1_1_L2_0_G1_MINI_ALU_BoothP_1), .A1 (WindowDin_1__0__0), .S0 (
             Instr)) ;
    mux21_ni ix1705 (.Y (L1_1_L2_0_G1_MINI_ALU_OperationResult_1), .A0 (
             L1_1_L2_0_G1_MINI_ALU_BoothP_2), .A1 (WindowDin_1__0__1), .S0 (
             Instr)) ;
    mux21_ni ix1713 (.Y (L1_1_L2_0_G1_MINI_ALU_OperationResult_2), .A0 (
             L1_1_L2_0_G1_MINI_ALU_BoothP_3), .A1 (WindowDin_1__0__2), .S0 (
             Instr)) ;
    mux21_ni ix1721 (.Y (L1_1_L2_0_G1_MINI_ALU_OperationResult_3), .A0 (
             L1_1_L2_0_G1_MINI_ALU_BoothP_4), .A1 (WindowDin_1__0__3), .S0 (
             Instr)) ;
    mux21_ni ix1729 (.Y (L1_1_L2_0_G1_MINI_ALU_OperationResult_4), .A0 (
             L1_1_L2_0_G1_MINI_ALU_BoothP_5), .A1 (WindowDin_1__0__4), .S0 (
             Instr)) ;
    mux21_ni ix1737 (.Y (L1_1_L2_0_G1_MINI_ALU_OperationResult_5), .A0 (
             L1_1_L2_0_G1_MINI_ALU_BoothP_6), .A1 (WindowDin_1__0__5), .S0 (
             Instr)) ;
    mux21_ni ix1745 (.Y (L1_1_L2_0_G1_MINI_ALU_OperationResult_6), .A0 (
             L1_1_L2_0_G1_MINI_ALU_BoothP_7), .A1 (WindowDin_1__0__6), .S0 (
             Instr)) ;
    mux21_ni ix1753 (.Y (L1_1_L2_0_G1_MINI_ALU_OperationResult_7), .A0 (
             L1_1_L2_0_G1_MINI_ALU_BoothP_8), .A1 (WindowDin_1__0__7), .S0 (
             Instr)) ;
    nor02ii ix1661 (.Y (L1_1_L2_0_G1_MINI_ALU_OperationResult_8), .A0 (Instr), .A1 (
            L1_1_L2_0_G1_MINI_ALU_BoothP_9)) ;
    nor02ii ix1665 (.Y (L1_1_L2_0_G1_MINI_ALU_OperationResult_9), .A0 (Instr), .A1 (
            L1_1_L2_0_G1_MINI_ALU_BoothP_10)) ;
    nor02ii ix1669 (.Y (L1_1_L2_0_G1_MINI_ALU_OperationResult_10), .A0 (Instr), 
            .A1 (L1_1_L2_0_G1_MINI_ALU_BoothP_11)) ;
    nor02ii ix1673 (.Y (L1_1_L2_0_G1_MINI_ALU_OperationResult_11), .A0 (Instr), 
            .A1 (L1_1_L2_0_G1_MINI_ALU_BoothP_12)) ;
    nor02ii ix1677 (.Y (L1_1_L2_0_G1_MINI_ALU_OperationResult_12), .A0 (Instr), 
            .A1 (L1_1_L2_0_G1_MINI_ALU_BoothP_13)) ;
    nor02ii ix1681 (.Y (L1_1_L2_0_G1_MINI_ALU_OperationResult_13), .A0 (Instr), 
            .A1 (L1_1_L2_0_G1_MINI_ALU_BoothP_14)) ;
    nor02ii ix1685 (.Y (L1_1_L2_0_G1_MINI_ALU_OperationResult_14), .A0 (Instr), 
            .A1 (L1_1_L2_0_G1_MINI_ALU_BoothP_15)) ;
    nor02ii ix1689 (.Y (L1_1_L2_0_G1_MINI_ALU_OperationResult_15), .A0 (Instr), 
            .A1 (L1_1_L2_0_G1_MINI_ALU_BoothP_16)) ;
    mux21_ni ix1793 (.Y (L1_0_L2_4_G1_MINI_ALU_OperationResult_0), .A0 (
             L1_0_L2_4_G1_MINI_ALU_BoothP_1), .A1 (WindowDin_0__4__0), .S0 (
             Instr)) ;
    mux21_ni ix1801 (.Y (L1_0_L2_4_G1_MINI_ALU_OperationResult_1), .A0 (
             L1_0_L2_4_G1_MINI_ALU_BoothP_2), .A1 (WindowDin_0__4__1), .S0 (
             Instr)) ;
    mux21_ni ix1809 (.Y (L1_0_L2_4_G1_MINI_ALU_OperationResult_2), .A0 (
             L1_0_L2_4_G1_MINI_ALU_BoothP_3), .A1 (WindowDin_0__4__2), .S0 (
             Instr)) ;
    mux21_ni ix1817 (.Y (L1_0_L2_4_G1_MINI_ALU_OperationResult_3), .A0 (
             L1_0_L2_4_G1_MINI_ALU_BoothP_4), .A1 (WindowDin_0__4__3), .S0 (
             Instr)) ;
    mux21_ni ix1825 (.Y (L1_0_L2_4_G1_MINI_ALU_OperationResult_4), .A0 (
             L1_0_L2_4_G1_MINI_ALU_BoothP_5), .A1 (WindowDin_0__4__4), .S0 (
             Instr)) ;
    mux21_ni ix1833 (.Y (L1_0_L2_4_G1_MINI_ALU_OperationResult_5), .A0 (
             L1_0_L2_4_G1_MINI_ALU_BoothP_6), .A1 (WindowDin_0__4__5), .S0 (
             Instr)) ;
    mux21_ni ix1841 (.Y (L1_0_L2_4_G1_MINI_ALU_OperationResult_6), .A0 (
             L1_0_L2_4_G1_MINI_ALU_BoothP_7), .A1 (WindowDin_0__4__6), .S0 (
             Instr)) ;
    mux21_ni ix1849 (.Y (L1_0_L2_4_G1_MINI_ALU_OperationResult_7), .A0 (
             L1_0_L2_4_G1_MINI_ALU_BoothP_8), .A1 (WindowDin_0__4__7), .S0 (
             Instr)) ;
    nor02ii ix1757 (.Y (L1_0_L2_4_G1_MINI_ALU_OperationResult_8), .A0 (Instr), .A1 (
            L1_0_L2_4_G1_MINI_ALU_BoothP_9)) ;
    nor02ii ix1761 (.Y (L1_0_L2_4_G1_MINI_ALU_OperationResult_9), .A0 (Instr), .A1 (
            L1_0_L2_4_G1_MINI_ALU_BoothP_10)) ;
    nor02ii ix1765 (.Y (L1_0_L2_4_G1_MINI_ALU_OperationResult_10), .A0 (Instr), 
            .A1 (L1_0_L2_4_G1_MINI_ALU_BoothP_11)) ;
    nor02ii ix1769 (.Y (L1_0_L2_4_G1_MINI_ALU_OperationResult_11), .A0 (Instr), 
            .A1 (L1_0_L2_4_G1_MINI_ALU_BoothP_12)) ;
    nor02ii ix1773 (.Y (L1_0_L2_4_G1_MINI_ALU_OperationResult_12), .A0 (Instr), 
            .A1 (L1_0_L2_4_G1_MINI_ALU_BoothP_13)) ;
    nor02ii ix1777 (.Y (L1_0_L2_4_G1_MINI_ALU_OperationResult_13), .A0 (Instr), 
            .A1 (L1_0_L2_4_G1_MINI_ALU_BoothP_14)) ;
    nor02ii ix1781 (.Y (L1_0_L2_4_G1_MINI_ALU_OperationResult_14), .A0 (Instr), 
            .A1 (L1_0_L2_4_G1_MINI_ALU_BoothP_15)) ;
    nor02ii ix1785 (.Y (L1_0_L2_4_G1_MINI_ALU_OperationResult_15), .A0 (Instr), 
            .A1 (L1_0_L2_4_G1_MINI_ALU_BoothP_16)) ;
    mux21_ni ix1889 (.Y (L1_0_L2_3_G1_MINI_ALU_OperationResult_0), .A0 (
             L1_0_L2_3_G1_MINI_ALU_BoothP_1), .A1 (WindowDin_0__3__0), .S0 (
             Instr)) ;
    mux21_ni ix1897 (.Y (L1_0_L2_3_G1_MINI_ALU_OperationResult_1), .A0 (
             L1_0_L2_3_G1_MINI_ALU_BoothP_2), .A1 (WindowDin_0__3__1), .S0 (
             Instr)) ;
    mux21_ni ix1905 (.Y (L1_0_L2_3_G1_MINI_ALU_OperationResult_2), .A0 (
             L1_0_L2_3_G1_MINI_ALU_BoothP_3), .A1 (WindowDin_0__3__2), .S0 (
             Instr)) ;
    mux21_ni ix1913 (.Y (L1_0_L2_3_G1_MINI_ALU_OperationResult_3), .A0 (
             L1_0_L2_3_G1_MINI_ALU_BoothP_4), .A1 (WindowDin_0__3__3), .S0 (
             Instr)) ;
    mux21_ni ix1921 (.Y (L1_0_L2_3_G1_MINI_ALU_OperationResult_4), .A0 (
             L1_0_L2_3_G1_MINI_ALU_BoothP_5), .A1 (WindowDin_0__3__4), .S0 (
             Instr)) ;
    mux21_ni ix1929 (.Y (L1_0_L2_3_G1_MINI_ALU_OperationResult_5), .A0 (
             L1_0_L2_3_G1_MINI_ALU_BoothP_6), .A1 (WindowDin_0__3__5), .S0 (
             Instr)) ;
    mux21_ni ix1937 (.Y (L1_0_L2_3_G1_MINI_ALU_OperationResult_6), .A0 (
             L1_0_L2_3_G1_MINI_ALU_BoothP_7), .A1 (WindowDin_0__3__6), .S0 (
             Instr)) ;
    mux21_ni ix1945 (.Y (L1_0_L2_3_G1_MINI_ALU_OperationResult_7), .A0 (
             L1_0_L2_3_G1_MINI_ALU_BoothP_8), .A1 (WindowDin_0__3__7), .S0 (
             Instr)) ;
    nor02ii ix1853 (.Y (L1_0_L2_3_G1_MINI_ALU_OperationResult_8), .A0 (Instr), .A1 (
            L1_0_L2_3_G1_MINI_ALU_BoothP_9)) ;
    nor02ii ix1857 (.Y (L1_0_L2_3_G1_MINI_ALU_OperationResult_9), .A0 (Instr), .A1 (
            L1_0_L2_3_G1_MINI_ALU_BoothP_10)) ;
    nor02ii ix1861 (.Y (L1_0_L2_3_G1_MINI_ALU_OperationResult_10), .A0 (Instr), 
            .A1 (L1_0_L2_3_G1_MINI_ALU_BoothP_11)) ;
    nor02ii ix1865 (.Y (L1_0_L2_3_G1_MINI_ALU_OperationResult_11), .A0 (Instr), 
            .A1 (L1_0_L2_3_G1_MINI_ALU_BoothP_12)) ;
    nor02ii ix1869 (.Y (L1_0_L2_3_G1_MINI_ALU_OperationResult_12), .A0 (Instr), 
            .A1 (L1_0_L2_3_G1_MINI_ALU_BoothP_13)) ;
    nor02ii ix1873 (.Y (L1_0_L2_3_G1_MINI_ALU_OperationResult_13), .A0 (Instr), 
            .A1 (L1_0_L2_3_G1_MINI_ALU_BoothP_14)) ;
    nor02ii ix1877 (.Y (L1_0_L2_3_G1_MINI_ALU_OperationResult_14), .A0 (Instr), 
            .A1 (L1_0_L2_3_G1_MINI_ALU_BoothP_15)) ;
    nor02ii ix1881 (.Y (L1_0_L2_3_G1_MINI_ALU_OperationResult_15), .A0 (Instr), 
            .A1 (L1_0_L2_3_G1_MINI_ALU_BoothP_16)) ;
    mux21_ni ix1985 (.Y (L1_0_L2_2_G1_MINI_ALU_OperationResult_0), .A0 (
             L1_0_L2_2_G1_MINI_ALU_BoothP_1), .A1 (WindowDin_0__2__0), .S0 (
             Instr)) ;
    mux21_ni ix1993 (.Y (L1_0_L2_2_G1_MINI_ALU_OperationResult_1), .A0 (
             L1_0_L2_2_G1_MINI_ALU_BoothP_2), .A1 (WindowDin_0__2__1), .S0 (
             Instr)) ;
    mux21_ni ix2001 (.Y (L1_0_L2_2_G1_MINI_ALU_OperationResult_2), .A0 (
             L1_0_L2_2_G1_MINI_ALU_BoothP_3), .A1 (WindowDin_0__2__2), .S0 (
             Instr)) ;
    mux21_ni ix2009 (.Y (L1_0_L2_2_G1_MINI_ALU_OperationResult_3), .A0 (
             L1_0_L2_2_G1_MINI_ALU_BoothP_4), .A1 (WindowDin_0__2__3), .S0 (
             Instr)) ;
    mux21_ni ix2017 (.Y (L1_0_L2_2_G1_MINI_ALU_OperationResult_4), .A0 (
             L1_0_L2_2_G1_MINI_ALU_BoothP_5), .A1 (WindowDin_0__2__4), .S0 (
             Instr)) ;
    mux21_ni ix2025 (.Y (L1_0_L2_2_G1_MINI_ALU_OperationResult_5), .A0 (
             L1_0_L2_2_G1_MINI_ALU_BoothP_6), .A1 (WindowDin_0__2__5), .S0 (
             Instr)) ;
    mux21_ni ix2033 (.Y (L1_0_L2_2_G1_MINI_ALU_OperationResult_6), .A0 (
             L1_0_L2_2_G1_MINI_ALU_BoothP_7), .A1 (WindowDin_0__2__6), .S0 (
             Instr)) ;
    mux21_ni ix2041 (.Y (L1_0_L2_2_G1_MINI_ALU_OperationResult_7), .A0 (
             L1_0_L2_2_G1_MINI_ALU_BoothP_8), .A1 (WindowDin_0__2__7), .S0 (
             Instr)) ;
    nor02ii ix1949 (.Y (L1_0_L2_2_G1_MINI_ALU_OperationResult_8), .A0 (Instr), .A1 (
            L1_0_L2_2_G1_MINI_ALU_BoothP_9)) ;
    nor02ii ix1953 (.Y (L1_0_L2_2_G1_MINI_ALU_OperationResult_9), .A0 (Instr), .A1 (
            L1_0_L2_2_G1_MINI_ALU_BoothP_10)) ;
    nor02ii ix1957 (.Y (L1_0_L2_2_G1_MINI_ALU_OperationResult_10), .A0 (Instr), 
            .A1 (L1_0_L2_2_G1_MINI_ALU_BoothP_11)) ;
    nor02ii ix1961 (.Y (L1_0_L2_2_G1_MINI_ALU_OperationResult_11), .A0 (Instr), 
            .A1 (L1_0_L2_2_G1_MINI_ALU_BoothP_12)) ;
    nor02ii ix1965 (.Y (L1_0_L2_2_G1_MINI_ALU_OperationResult_12), .A0 (Instr), 
            .A1 (L1_0_L2_2_G1_MINI_ALU_BoothP_13)) ;
    nor02ii ix1969 (.Y (L1_0_L2_2_G1_MINI_ALU_OperationResult_13), .A0 (Instr), 
            .A1 (L1_0_L2_2_G1_MINI_ALU_BoothP_14)) ;
    nor02ii ix1973 (.Y (L1_0_L2_2_G1_MINI_ALU_OperationResult_14), .A0 (Instr), 
            .A1 (L1_0_L2_2_G1_MINI_ALU_BoothP_15)) ;
    nor02ii ix1977 (.Y (L1_0_L2_2_G1_MINI_ALU_OperationResult_15), .A0 (Instr), 
            .A1 (L1_0_L2_2_G1_MINI_ALU_BoothP_16)) ;
    mux21_ni ix2081 (.Y (L1_0_L2_1_G1_MINI_ALU_OperationResult_0), .A0 (
             L1_0_L2_1_G1_MINI_ALU_BoothP_1), .A1 (WindowDin_0__1__0), .S0 (
             Instr)) ;
    mux21_ni ix2089 (.Y (L1_0_L2_1_G1_MINI_ALU_OperationResult_1), .A0 (
             L1_0_L2_1_G1_MINI_ALU_BoothP_2), .A1 (WindowDin_0__1__1), .S0 (
             Instr)) ;
    mux21_ni ix2097 (.Y (L1_0_L2_1_G1_MINI_ALU_OperationResult_2), .A0 (
             L1_0_L2_1_G1_MINI_ALU_BoothP_3), .A1 (WindowDin_0__1__2), .S0 (
             Instr)) ;
    mux21_ni ix2105 (.Y (L1_0_L2_1_G1_MINI_ALU_OperationResult_3), .A0 (
             L1_0_L2_1_G1_MINI_ALU_BoothP_4), .A1 (WindowDin_0__1__3), .S0 (
             Instr)) ;
    mux21_ni ix2113 (.Y (L1_0_L2_1_G1_MINI_ALU_OperationResult_4), .A0 (
             L1_0_L2_1_G1_MINI_ALU_BoothP_5), .A1 (WindowDin_0__1__4), .S0 (
             Instr)) ;
    mux21_ni ix2121 (.Y (L1_0_L2_1_G1_MINI_ALU_OperationResult_5), .A0 (
             L1_0_L2_1_G1_MINI_ALU_BoothP_6), .A1 (WindowDin_0__1__5), .S0 (
             Instr)) ;
    mux21_ni ix2129 (.Y (L1_0_L2_1_G1_MINI_ALU_OperationResult_6), .A0 (
             L1_0_L2_1_G1_MINI_ALU_BoothP_7), .A1 (WindowDin_0__1__6), .S0 (
             Instr)) ;
    mux21_ni ix2137 (.Y (L1_0_L2_1_G1_MINI_ALU_OperationResult_7), .A0 (
             L1_0_L2_1_G1_MINI_ALU_BoothP_8), .A1 (WindowDin_0__1__7), .S0 (
             Instr)) ;
    nor02ii ix2045 (.Y (L1_0_L2_1_G1_MINI_ALU_OperationResult_8), .A0 (Instr), .A1 (
            L1_0_L2_1_G1_MINI_ALU_BoothP_9)) ;
    nor02ii ix2049 (.Y (L1_0_L2_1_G1_MINI_ALU_OperationResult_9), .A0 (Instr), .A1 (
            L1_0_L2_1_G1_MINI_ALU_BoothP_10)) ;
    nor02ii ix2053 (.Y (L1_0_L2_1_G1_MINI_ALU_OperationResult_10), .A0 (Instr), 
            .A1 (L1_0_L2_1_G1_MINI_ALU_BoothP_11)) ;
    nor02ii ix2057 (.Y (L1_0_L2_1_G1_MINI_ALU_OperationResult_11), .A0 (Instr), 
            .A1 (L1_0_L2_1_G1_MINI_ALU_BoothP_12)) ;
    nor02ii ix2061 (.Y (L1_0_L2_1_G1_MINI_ALU_OperationResult_12), .A0 (Instr), 
            .A1 (L1_0_L2_1_G1_MINI_ALU_BoothP_13)) ;
    nor02ii ix2065 (.Y (L1_0_L2_1_G1_MINI_ALU_OperationResult_13), .A0 (Instr), 
            .A1 (L1_0_L2_1_G1_MINI_ALU_BoothP_14)) ;
    nor02ii ix2069 (.Y (L1_0_L2_1_G1_MINI_ALU_OperationResult_14), .A0 (Instr), 
            .A1 (L1_0_L2_1_G1_MINI_ALU_BoothP_15)) ;
    nor02ii ix2073 (.Y (L1_0_L2_1_G1_MINI_ALU_OperationResult_15), .A0 (Instr), 
            .A1 (L1_0_L2_1_G1_MINI_ALU_BoothP_16)) ;
    mux21_ni ix2177 (.Y (L1_0_L2_0_G1_MINI_ALU_OperationResult_0), .A0 (
             L1_0_L2_0_G1_MINI_ALU_BoothP_1), .A1 (WindowDin_0__0__0), .S0 (
             Instr)) ;
    mux21_ni ix2185 (.Y (L1_0_L2_0_G1_MINI_ALU_OperationResult_1), .A0 (
             L1_0_L2_0_G1_MINI_ALU_BoothP_2), .A1 (WindowDin_0__0__1), .S0 (
             Instr)) ;
    mux21_ni ix2193 (.Y (L1_0_L2_0_G1_MINI_ALU_OperationResult_2), .A0 (
             L1_0_L2_0_G1_MINI_ALU_BoothP_3), .A1 (WindowDin_0__0__2), .S0 (
             Instr)) ;
    mux21_ni ix2201 (.Y (L1_0_L2_0_G1_MINI_ALU_OperationResult_3), .A0 (
             L1_0_L2_0_G1_MINI_ALU_BoothP_4), .A1 (WindowDin_0__0__3), .S0 (
             Instr)) ;
    mux21_ni ix2209 (.Y (L1_0_L2_0_G1_MINI_ALU_OperationResult_4), .A0 (
             L1_0_L2_0_G1_MINI_ALU_BoothP_5), .A1 (WindowDin_0__0__4), .S0 (
             Instr)) ;
    mux21_ni ix2217 (.Y (L1_0_L2_0_G1_MINI_ALU_OperationResult_5), .A0 (
             L1_0_L2_0_G1_MINI_ALU_BoothP_6), .A1 (WindowDin_0__0__5), .S0 (
             Instr)) ;
    mux21_ni ix2225 (.Y (L1_0_L2_0_G1_MINI_ALU_OperationResult_6), .A0 (
             L1_0_L2_0_G1_MINI_ALU_BoothP_7), .A1 (WindowDin_0__0__6), .S0 (
             Instr)) ;
    mux21_ni ix2233 (.Y (L1_0_L2_0_G1_MINI_ALU_OperationResult_7), .A0 (
             L1_0_L2_0_G1_MINI_ALU_BoothP_8), .A1 (WindowDin_0__0__7), .S0 (
             Instr)) ;
    nor02ii ix2141 (.Y (L1_0_L2_0_G1_MINI_ALU_OperationResult_8), .A0 (Instr), .A1 (
            L1_0_L2_0_G1_MINI_ALU_BoothP_9)) ;
    nor02ii ix2145 (.Y (L1_0_L2_0_G1_MINI_ALU_OperationResult_9), .A0 (Instr), .A1 (
            L1_0_L2_0_G1_MINI_ALU_BoothP_10)) ;
    nor02ii ix2149 (.Y (L1_0_L2_0_G1_MINI_ALU_OperationResult_10), .A0 (Instr), 
            .A1 (L1_0_L2_0_G1_MINI_ALU_BoothP_11)) ;
    nor02ii ix2153 (.Y (L1_0_L2_0_G1_MINI_ALU_OperationResult_11), .A0 (Instr), 
            .A1 (L1_0_L2_0_G1_MINI_ALU_BoothP_12)) ;
    nor02ii ix2157 (.Y (L1_0_L2_0_G1_MINI_ALU_OperationResult_12), .A0 (Instr), 
            .A1 (L1_0_L2_0_G1_MINI_ALU_BoothP_13)) ;
    nor02ii ix2161 (.Y (L1_0_L2_0_G1_MINI_ALU_OperationResult_13), .A0 (Instr), 
            .A1 (L1_0_L2_0_G1_MINI_ALU_BoothP_14)) ;
    nor02ii ix2165 (.Y (L1_0_L2_0_G1_MINI_ALU_OperationResult_14), .A0 (Instr), 
            .A1 (L1_0_L2_0_G1_MINI_ALU_BoothP_15)) ;
    nor02ii ix2169 (.Y (L1_0_L2_0_G1_MINI_ALU_OperationResult_15), .A0 (Instr), 
            .A1 (L1_0_L2_0_G1_MINI_ALU_BoothP_16)) ;
    mux21_ni ix973 (.Y (L1FirstOperands_11__0), .A0 (
             L1_2_L2_2_G1_MINI_ALU_BoothP_1), .A1 (WindowDin_2__2__0), .S0 (
             Instr)) ;
    mux21_ni ix981 (.Y (L1FirstOperands_11__1), .A0 (
             L1_2_L2_2_G1_MINI_ALU_BoothP_2), .A1 (WindowDin_2__2__1), .S0 (
             Instr)) ;
    mux21_ni ix989 (.Y (L1FirstOperands_11__2), .A0 (
             L1_2_L2_2_G1_MINI_ALU_BoothP_3), .A1 (WindowDin_2__2__2), .S0 (
             Instr)) ;
    mux21_ni ix997 (.Y (L1FirstOperands_11__3), .A0 (
             L1_2_L2_2_G1_MINI_ALU_BoothP_4), .A1 (WindowDin_2__2__3), .S0 (
             Instr)) ;
    mux21_ni ix1005 (.Y (L1FirstOperands_11__4), .A0 (
             L1_2_L2_2_G1_MINI_ALU_BoothP_5), .A1 (WindowDin_2__2__4), .S0 (
             Instr)) ;
    mux21_ni ix1013 (.Y (L1FirstOperands_11__5), .A0 (
             L1_2_L2_2_G1_MINI_ALU_BoothP_6), .A1 (WindowDin_2__2__5), .S0 (
             Instr)) ;
    mux21_ni ix1021 (.Y (L1FirstOperands_11__6), .A0 (
             L1_2_L2_2_G1_MINI_ALU_BoothP_7), .A1 (WindowDin_2__2__6), .S0 (
             Instr)) ;
    mux21_ni ix1029 (.Y (L1FirstOperands_11__7), .A0 (
             L1_2_L2_2_G1_MINI_ALU_BoothP_8), .A1 (WindowDin_2__2__7), .S0 (
             Instr)) ;
    nor02ii ix937 (.Y (L1FirstOperands_11__8), .A0 (Instr), .A1 (
            L1_2_L2_2_G1_MINI_ALU_BoothP_9)) ;
    nor02ii ix941 (.Y (L1FirstOperands_11__9), .A0 (Instr), .A1 (
            L1_2_L2_2_G1_MINI_ALU_BoothP_10)) ;
    nor02ii ix945 (.Y (L1FirstOperands_11__10), .A0 (Instr), .A1 (
            L1_2_L2_2_G1_MINI_ALU_BoothP_11)) ;
    nor02ii ix949 (.Y (L1FirstOperands_11__11), .A0 (Instr), .A1 (
            L1_2_L2_2_G1_MINI_ALU_BoothP_12)) ;
    nor02ii ix953 (.Y (L1FirstOperands_11__12), .A0 (Instr), .A1 (
            L1_2_L2_2_G1_MINI_ALU_BoothP_13)) ;
    nor02ii ix957 (.Y (L1FirstOperands_11__13), .A0 (Instr), .A1 (
            L1_2_L2_2_G1_MINI_ALU_BoothP_14)) ;
    nor02ii ix961 (.Y (L1FirstOperands_11__14), .A0 (Instr), .A1 (
            L1_2_L2_2_G1_MINI_ALU_BoothP_15)) ;
    nor02ii ix965 (.Y (L1FirstOperands_11__15), .A0 (Instr), .A1 (
            L1_2_L2_2_G1_MINI_ALU_BoothP_16)) ;
    mux21_ni ix397 (.Y (L1FirstOperands_10__0), .A0 (
             L1_3_L2_3_G2_MINI_ALU_BoothP_1), .A1 (WindowDin_3__3__0), .S0 (
             Instr)) ;
    mux21_ni ix405 (.Y (L1FirstOperands_10__1), .A0 (
             L1_3_L2_3_G2_MINI_ALU_BoothP_2), .A1 (WindowDin_3__3__1), .S0 (
             Instr)) ;
    mux21_ni ix413 (.Y (L1FirstOperands_10__2), .A0 (
             L1_3_L2_3_G2_MINI_ALU_BoothP_3), .A1 (WindowDin_3__3__2), .S0 (
             Instr)) ;
    mux21_ni ix421 (.Y (L1FirstOperands_10__3), .A0 (
             L1_3_L2_3_G2_MINI_ALU_BoothP_4), .A1 (WindowDin_3__3__3), .S0 (
             Instr)) ;
    mux21_ni ix429 (.Y (L1FirstOperands_10__4), .A0 (
             L1_3_L2_3_G2_MINI_ALU_BoothP_5), .A1 (WindowDin_3__3__4), .S0 (
             Instr)) ;
    mux21_ni ix437 (.Y (L1FirstOperands_10__5), .A0 (
             L1_3_L2_3_G2_MINI_ALU_BoothP_6), .A1 (WindowDin_3__3__5), .S0 (
             Instr)) ;
    mux21_ni ix445 (.Y (L1FirstOperands_10__6), .A0 (
             L1_3_L2_3_G2_MINI_ALU_BoothP_7), .A1 (WindowDin_3__3__6), .S0 (
             Instr)) ;
    mux21_ni ix453 (.Y (L1FirstOperands_10__7), .A0 (
             L1_3_L2_3_G2_MINI_ALU_BoothP_8), .A1 (WindowDin_3__3__7), .S0 (
             Instr)) ;
    nor02ii ix361 (.Y (L1FirstOperands_10__8), .A0 (Instr), .A1 (
            L1_3_L2_3_G2_MINI_ALU_BoothP_9)) ;
    nor02ii ix365 (.Y (L1FirstOperands_10__9), .A0 (Instr), .A1 (
            L1_3_L2_3_G2_MINI_ALU_BoothP_10)) ;
    nor02ii ix369 (.Y (L1FirstOperands_10__10), .A0 (Instr), .A1 (
            L1_3_L2_3_G2_MINI_ALU_BoothP_11)) ;
    nor02ii ix373 (.Y (L1FirstOperands_10__11), .A0 (Instr), .A1 (
            L1_3_L2_3_G2_MINI_ALU_BoothP_12)) ;
    nor02ii ix377 (.Y (L1FirstOperands_10__12), .A0 (Instr), .A1 (
            L1_3_L2_3_G2_MINI_ALU_BoothP_13)) ;
    nor02ii ix381 (.Y (L1FirstOperands_10__13), .A0 (Instr), .A1 (
            L1_3_L2_3_G2_MINI_ALU_BoothP_14)) ;
    nor02ii ix385 (.Y (L1FirstOperands_10__14), .A0 (Instr), .A1 (
            L1_3_L2_3_G2_MINI_ALU_BoothP_15)) ;
    nor02ii ix389 (.Y (L1FirstOperands_10__15), .A0 (Instr), .A1 (
            L1_3_L2_3_G2_MINI_ALU_BoothP_16)) ;
    mux21_ni ix493 (.Y (L1FirstOperands_8__0), .A0 (
             L1_3_L2_2_G2_MINI_ALU_BoothP_1), .A1 (WindowDin_3__2__0), .S0 (
             Instr)) ;
    mux21_ni ix501 (.Y (L1FirstOperands_8__1), .A0 (
             L1_3_L2_2_G2_MINI_ALU_BoothP_2), .A1 (WindowDin_3__2__1), .S0 (
             Instr)) ;
    mux21_ni ix509 (.Y (L1FirstOperands_8__2), .A0 (
             L1_3_L2_2_G2_MINI_ALU_BoothP_3), .A1 (WindowDin_3__2__2), .S0 (
             Instr)) ;
    mux21_ni ix517 (.Y (L1FirstOperands_8__3), .A0 (
             L1_3_L2_2_G2_MINI_ALU_BoothP_4), .A1 (WindowDin_3__2__3), .S0 (
             Instr)) ;
    mux21_ni ix525 (.Y (L1FirstOperands_8__4), .A0 (
             L1_3_L2_2_G2_MINI_ALU_BoothP_5), .A1 (WindowDin_3__2__4), .S0 (
             Instr)) ;
    mux21_ni ix533 (.Y (L1FirstOperands_8__5), .A0 (
             L1_3_L2_2_G2_MINI_ALU_BoothP_6), .A1 (WindowDin_3__2__5), .S0 (
             Instr)) ;
    mux21_ni ix541 (.Y (L1FirstOperands_8__6), .A0 (
             L1_3_L2_2_G2_MINI_ALU_BoothP_7), .A1 (WindowDin_3__2__6), .S0 (
             Instr)) ;
    mux21_ni ix549 (.Y (L1FirstOperands_8__7), .A0 (
             L1_3_L2_2_G2_MINI_ALU_BoothP_8), .A1 (WindowDin_3__2__7), .S0 (
             Instr)) ;
    nor02ii ix457 (.Y (L1FirstOperands_8__8), .A0 (Instr), .A1 (
            L1_3_L2_2_G2_MINI_ALU_BoothP_9)) ;
    nor02ii ix461 (.Y (L1FirstOperands_8__9), .A0 (Instr), .A1 (
            L1_3_L2_2_G2_MINI_ALU_BoothP_10)) ;
    nor02ii ix465 (.Y (L1FirstOperands_8__10), .A0 (Instr), .A1 (
            L1_3_L2_2_G2_MINI_ALU_BoothP_11)) ;
    nor02ii ix469 (.Y (L1FirstOperands_8__11), .A0 (Instr), .A1 (
            L1_3_L2_2_G2_MINI_ALU_BoothP_12)) ;
    nor02ii ix473 (.Y (L1FirstOperands_8__12), .A0 (Instr), .A1 (
            L1_3_L2_2_G2_MINI_ALU_BoothP_13)) ;
    nor02ii ix477 (.Y (L1FirstOperands_8__13), .A0 (Instr), .A1 (
            L1_3_L2_2_G2_MINI_ALU_BoothP_14)) ;
    nor02ii ix481 (.Y (L1FirstOperands_8__14), .A0 (Instr), .A1 (
            L1_3_L2_2_G2_MINI_ALU_BoothP_15)) ;
    nor02ii ix485 (.Y (L1FirstOperands_8__15), .A0 (Instr), .A1 (
            L1_3_L2_2_G2_MINI_ALU_BoothP_16)) ;
    mux21_ni ix205 (.Y (L1FirstOperands_7__0), .A0 (
             L1_4_L2_3_G5_MINI_ALU_BoothP_1), .A1 (WindowDin_4__3__0), .S0 (
             Instr)) ;
    mux21_ni ix213 (.Y (L1FirstOperands_7__1), .A0 (
             L1_4_L2_3_G5_MINI_ALU_BoothP_2), .A1 (WindowDin_4__3__1), .S0 (
             Instr)) ;
    mux21_ni ix221 (.Y (L1FirstOperands_7__2), .A0 (
             L1_4_L2_3_G5_MINI_ALU_BoothP_3), .A1 (WindowDin_4__3__2), .S0 (
             Instr)) ;
    mux21_ni ix229 (.Y (L1FirstOperands_7__3), .A0 (
             L1_4_L2_3_G5_MINI_ALU_BoothP_4), .A1 (WindowDin_4__3__3), .S0 (
             Instr)) ;
    mux21_ni ix237 (.Y (L1FirstOperands_7__4), .A0 (
             L1_4_L2_3_G5_MINI_ALU_BoothP_5), .A1 (WindowDin_4__3__4), .S0 (
             Instr)) ;
    mux21_ni ix245 (.Y (L1FirstOperands_7__5), .A0 (
             L1_4_L2_3_G5_MINI_ALU_BoothP_6), .A1 (WindowDin_4__3__5), .S0 (
             Instr)) ;
    mux21_ni ix253 (.Y (L1FirstOperands_7__6), .A0 (
             L1_4_L2_3_G5_MINI_ALU_BoothP_7), .A1 (WindowDin_4__3__6), .S0 (
             Instr)) ;
    mux21_ni ix261 (.Y (L1FirstOperands_7__7), .A0 (
             L1_4_L2_3_G5_MINI_ALU_BoothP_8), .A1 (WindowDin_4__3__7), .S0 (
             Instr)) ;
    nor02ii ix169 (.Y (L1FirstOperands_7__8), .A0 (Instr), .A1 (
            L1_4_L2_3_G5_MINI_ALU_BoothP_9)) ;
    nor02ii ix173 (.Y (L1FirstOperands_7__9), .A0 (Instr), .A1 (
            L1_4_L2_3_G5_MINI_ALU_BoothP_10)) ;
    nor02ii ix177 (.Y (L1FirstOperands_7__10), .A0 (Instr), .A1 (
            L1_4_L2_3_G5_MINI_ALU_BoothP_11)) ;
    nor02ii ix181 (.Y (L1FirstOperands_7__11), .A0 (Instr), .A1 (
            L1_4_L2_3_G5_MINI_ALU_BoothP_12)) ;
    nor02ii ix185 (.Y (L1FirstOperands_7__12), .A0 (Instr), .A1 (
            L1_4_L2_3_G5_MINI_ALU_BoothP_13)) ;
    nor02ii ix189 (.Y (L1FirstOperands_7__13), .A0 (Instr), .A1 (
            L1_4_L2_3_G5_MINI_ALU_BoothP_14)) ;
    nor02ii ix193 (.Y (L1FirstOperands_7__14), .A0 (Instr), .A1 (
            L1_4_L2_3_G5_MINI_ALU_BoothP_15)) ;
    nor02ii ix197 (.Y (L1FirstOperands_7__15), .A0 (Instr), .A1 (
            L1_4_L2_3_G5_MINI_ALU_BoothP_16)) ;
    mux21_ni ix589 (.Y (L1FirstOperands_6__0), .A0 (
             L1_3_L2_1_G2_MINI_ALU_BoothP_1), .A1 (WindowDin_3__1__0), .S0 (
             Instr)) ;
    mux21_ni ix597 (.Y (L1FirstOperands_6__1), .A0 (
             L1_3_L2_1_G2_MINI_ALU_BoothP_2), .A1 (WindowDin_3__1__1), .S0 (
             Instr)) ;
    mux21_ni ix605 (.Y (L1FirstOperands_6__2), .A0 (
             L1_3_L2_1_G2_MINI_ALU_BoothP_3), .A1 (WindowDin_3__1__2), .S0 (
             Instr)) ;
    mux21_ni ix613 (.Y (L1FirstOperands_6__3), .A0 (
             L1_3_L2_1_G2_MINI_ALU_BoothP_4), .A1 (WindowDin_3__1__3), .S0 (
             Instr)) ;
    mux21_ni ix621 (.Y (L1FirstOperands_6__4), .A0 (
             L1_3_L2_1_G2_MINI_ALU_BoothP_5), .A1 (WindowDin_3__1__4), .S0 (
             Instr)) ;
    mux21_ni ix629 (.Y (L1FirstOperands_6__5), .A0 (
             L1_3_L2_1_G2_MINI_ALU_BoothP_6), .A1 (WindowDin_3__1__5), .S0 (
             Instr)) ;
    mux21_ni ix637 (.Y (L1FirstOperands_6__6), .A0 (
             L1_3_L2_1_G2_MINI_ALU_BoothP_7), .A1 (WindowDin_3__1__6), .S0 (
             Instr)) ;
    mux21_ni ix645 (.Y (L1FirstOperands_6__7), .A0 (
             L1_3_L2_1_G2_MINI_ALU_BoothP_8), .A1 (WindowDin_3__1__7), .S0 (
             Instr)) ;
    nor02ii ix553 (.Y (L1FirstOperands_6__8), .A0 (Instr), .A1 (
            L1_3_L2_1_G2_MINI_ALU_BoothP_9)) ;
    nor02ii ix557 (.Y (L1FirstOperands_6__9), .A0 (Instr), .A1 (
            L1_3_L2_1_G2_MINI_ALU_BoothP_10)) ;
    nor02ii ix561 (.Y (L1FirstOperands_6__10), .A0 (Instr), .A1 (
            L1_3_L2_1_G2_MINI_ALU_BoothP_11)) ;
    nor02ii ix565 (.Y (L1FirstOperands_6__11), .A0 (Instr), .A1 (
            L1_3_L2_1_G2_MINI_ALU_BoothP_12)) ;
    nor02ii ix569 (.Y (L1FirstOperands_6__12), .A0 (Instr), .A1 (
            L1_3_L2_1_G2_MINI_ALU_BoothP_13)) ;
    nor02ii ix573 (.Y (L1FirstOperands_6__13), .A0 (Instr), .A1 (
            L1_3_L2_1_G2_MINI_ALU_BoothP_14)) ;
    nor02ii ix577 (.Y (L1FirstOperands_6__14), .A0 (Instr), .A1 (
            L1_3_L2_1_G2_MINI_ALU_BoothP_15)) ;
    nor02ii ix581 (.Y (L1FirstOperands_6__15), .A0 (Instr), .A1 (
            L1_3_L2_1_G2_MINI_ALU_BoothP_16)) ;
    mux21_ni ix685 (.Y (L1FirstOperands_4__0), .A0 (
             L1_3_L2_0_G2_MINI_ALU_BoothP_1), .A1 (WindowDin_3__0__0), .S0 (
             Instr)) ;
    mux21_ni ix693 (.Y (L1FirstOperands_4__1), .A0 (
             L1_3_L2_0_G2_MINI_ALU_BoothP_2), .A1 (WindowDin_3__0__1), .S0 (
             Instr)) ;
    mux21_ni ix701 (.Y (L1FirstOperands_4__2), .A0 (
             L1_3_L2_0_G2_MINI_ALU_BoothP_3), .A1 (WindowDin_3__0__2), .S0 (
             Instr)) ;
    mux21_ni ix709 (.Y (L1FirstOperands_4__3), .A0 (
             L1_3_L2_0_G2_MINI_ALU_BoothP_4), .A1 (WindowDin_3__0__3), .S0 (
             Instr)) ;
    mux21_ni ix717 (.Y (L1FirstOperands_4__4), .A0 (
             L1_3_L2_0_G2_MINI_ALU_BoothP_5), .A1 (WindowDin_3__0__4), .S0 (
             Instr)) ;
    mux21_ni ix725 (.Y (L1FirstOperands_4__5), .A0 (
             L1_3_L2_0_G2_MINI_ALU_BoothP_6), .A1 (WindowDin_3__0__5), .S0 (
             Instr)) ;
    mux21_ni ix733 (.Y (L1FirstOperands_4__6), .A0 (
             L1_3_L2_0_G2_MINI_ALU_BoothP_7), .A1 (WindowDin_3__0__6), .S0 (
             Instr)) ;
    mux21_ni ix741 (.Y (L1FirstOperands_4__7), .A0 (
             L1_3_L2_0_G2_MINI_ALU_BoothP_8), .A1 (WindowDin_3__0__7), .S0 (
             Instr)) ;
    nor02ii ix649 (.Y (L1FirstOperands_4__8), .A0 (Instr), .A1 (
            L1_3_L2_0_G2_MINI_ALU_BoothP_9)) ;
    nor02ii ix653 (.Y (L1FirstOperands_4__9), .A0 (Instr), .A1 (
            L1_3_L2_0_G2_MINI_ALU_BoothP_10)) ;
    nor02ii ix657 (.Y (L1FirstOperands_4__10), .A0 (Instr), .A1 (
            L1_3_L2_0_G2_MINI_ALU_BoothP_11)) ;
    nor02ii ix661 (.Y (L1FirstOperands_4__11), .A0 (Instr), .A1 (
            L1_3_L2_0_G2_MINI_ALU_BoothP_12)) ;
    nor02ii ix665 (.Y (L1FirstOperands_4__12), .A0 (Instr), .A1 (
            L1_3_L2_0_G2_MINI_ALU_BoothP_13)) ;
    nor02ii ix669 (.Y (L1FirstOperands_4__13), .A0 (Instr), .A1 (
            L1_3_L2_0_G2_MINI_ALU_BoothP_14)) ;
    nor02ii ix673 (.Y (L1FirstOperands_4__14), .A0 (Instr), .A1 (
            L1_3_L2_0_G2_MINI_ALU_BoothP_15)) ;
    nor02ii ix677 (.Y (L1FirstOperands_4__15), .A0 (Instr), .A1 (
            L1_3_L2_0_G2_MINI_ALU_BoothP_16)) ;
    mux21_ni ix301 (.Y (L1FirstOperands_3__0), .A0 (
             L1_4_L2_2_G4_MINI_ALU_BoothP_1), .A1 (WindowDin_4__2__0), .S0 (
             Instr)) ;
    mux21_ni ix309 (.Y (L1FirstOperands_3__1), .A0 (
             L1_4_L2_2_G4_MINI_ALU_BoothP_2), .A1 (WindowDin_4__2__1), .S0 (
             Instr)) ;
    mux21_ni ix317 (.Y (L1FirstOperands_3__2), .A0 (
             L1_4_L2_2_G4_MINI_ALU_BoothP_3), .A1 (WindowDin_4__2__2), .S0 (
             Instr)) ;
    mux21_ni ix325 (.Y (L1FirstOperands_3__3), .A0 (
             L1_4_L2_2_G4_MINI_ALU_BoothP_4), .A1 (WindowDin_4__2__3), .S0 (
             Instr)) ;
    mux21_ni ix333 (.Y (L1FirstOperands_3__4), .A0 (
             L1_4_L2_2_G4_MINI_ALU_BoothP_5), .A1 (WindowDin_4__2__4), .S0 (
             Instr)) ;
    mux21_ni ix341 (.Y (L1FirstOperands_3__5), .A0 (
             L1_4_L2_2_G4_MINI_ALU_BoothP_6), .A1 (WindowDin_4__2__5), .S0 (
             Instr)) ;
    mux21_ni ix349 (.Y (L1FirstOperands_3__6), .A0 (
             L1_4_L2_2_G4_MINI_ALU_BoothP_7), .A1 (WindowDin_4__2__6), .S0 (
             Instr)) ;
    mux21_ni ix357 (.Y (L1FirstOperands_3__7), .A0 (
             L1_4_L2_2_G4_MINI_ALU_BoothP_8), .A1 (WindowDin_4__2__7), .S0 (
             Instr)) ;
    nor02ii ix265 (.Y (L1FirstOperands_3__8), .A0 (Instr), .A1 (
            L1_4_L2_2_G4_MINI_ALU_BoothP_9)) ;
    nor02ii ix269 (.Y (L1FirstOperands_3__9), .A0 (Instr), .A1 (
            L1_4_L2_2_G4_MINI_ALU_BoothP_10)) ;
    nor02ii ix273 (.Y (L1FirstOperands_3__10), .A0 (Instr), .A1 (
            L1_4_L2_2_G4_MINI_ALU_BoothP_11)) ;
    nor02ii ix277 (.Y (L1FirstOperands_3__11), .A0 (Instr), .A1 (
            L1_4_L2_2_G4_MINI_ALU_BoothP_12)) ;
    nor02ii ix281 (.Y (L1FirstOperands_3__12), .A0 (Instr), .A1 (
            L1_4_L2_2_G4_MINI_ALU_BoothP_13)) ;
    nor02ii ix285 (.Y (L1FirstOperands_3__13), .A0 (Instr), .A1 (
            L1_4_L2_2_G4_MINI_ALU_BoothP_14)) ;
    nor02ii ix289 (.Y (L1FirstOperands_3__14), .A0 (Instr), .A1 (
            L1_4_L2_2_G4_MINI_ALU_BoothP_15)) ;
    nor02ii ix293 (.Y (L1FirstOperands_3__15), .A0 (Instr), .A1 (
            L1_4_L2_2_G4_MINI_ALU_BoothP_16)) ;
    mux21_ni ix781 (.Y (L1FirstOperands_2__0), .A0 (
             L1_2_L2_4_G2_MINI_ALU_BoothP_1), .A1 (WindowDin_2__4__0), .S0 (
             Instr)) ;
    mux21_ni ix789 (.Y (L1FirstOperands_2__1), .A0 (
             L1_2_L2_4_G2_MINI_ALU_BoothP_2), .A1 (WindowDin_2__4__1), .S0 (
             Instr)) ;
    mux21_ni ix797 (.Y (L1FirstOperands_2__2), .A0 (
             L1_2_L2_4_G2_MINI_ALU_BoothP_3), .A1 (WindowDin_2__4__2), .S0 (
             Instr)) ;
    mux21_ni ix805 (.Y (L1FirstOperands_2__3), .A0 (
             L1_2_L2_4_G2_MINI_ALU_BoothP_4), .A1 (WindowDin_2__4__3), .S0 (
             Instr)) ;
    mux21_ni ix813 (.Y (L1FirstOperands_2__4), .A0 (
             L1_2_L2_4_G2_MINI_ALU_BoothP_5), .A1 (WindowDin_2__4__4), .S0 (
             Instr)) ;
    mux21_ni ix821 (.Y (L1FirstOperands_2__5), .A0 (
             L1_2_L2_4_G2_MINI_ALU_BoothP_6), .A1 (WindowDin_2__4__5), .S0 (
             Instr)) ;
    mux21_ni ix829 (.Y (L1FirstOperands_2__6), .A0 (
             L1_2_L2_4_G2_MINI_ALU_BoothP_7), .A1 (WindowDin_2__4__6), .S0 (
             Instr)) ;
    mux21_ni ix837 (.Y (L1FirstOperands_2__7), .A0 (
             L1_2_L2_4_G2_MINI_ALU_BoothP_8), .A1 (WindowDin_2__4__7), .S0 (
             Instr)) ;
    nor02ii ix745 (.Y (L1FirstOperands_2__8), .A0 (Instr), .A1 (
            L1_2_L2_4_G2_MINI_ALU_BoothP_9)) ;
    nor02ii ix749 (.Y (L1FirstOperands_2__9), .A0 (Instr), .A1 (
            L1_2_L2_4_G2_MINI_ALU_BoothP_10)) ;
    nor02ii ix753 (.Y (L1FirstOperands_2__10), .A0 (Instr), .A1 (
            L1_2_L2_4_G2_MINI_ALU_BoothP_11)) ;
    nor02ii ix757 (.Y (L1FirstOperands_2__11), .A0 (Instr), .A1 (
            L1_2_L2_4_G2_MINI_ALU_BoothP_12)) ;
    nor02ii ix761 (.Y (L1FirstOperands_2__12), .A0 (Instr), .A1 (
            L1_2_L2_4_G2_MINI_ALU_BoothP_13)) ;
    nor02ii ix765 (.Y (L1FirstOperands_2__13), .A0 (Instr), .A1 (
            L1_2_L2_4_G2_MINI_ALU_BoothP_14)) ;
    nor02ii ix769 (.Y (L1FirstOperands_2__14), .A0 (Instr), .A1 (
            L1_2_L2_4_G2_MINI_ALU_BoothP_15)) ;
    nor02ii ix773 (.Y (L1FirstOperands_2__15), .A0 (Instr), .A1 (
            L1_2_L2_4_G2_MINI_ALU_BoothP_16)) ;
    mux21_ni ix877 (.Y (L1FirstOperands_0__0), .A0 (
             L1_2_L2_3_G2_MINI_ALU_BoothP_1), .A1 (WindowDin_2__3__0), .S0 (
             Instr)) ;
    mux21_ni ix885 (.Y (L1FirstOperands_0__1), .A0 (
             L1_2_L2_3_G2_MINI_ALU_BoothP_2), .A1 (WindowDin_2__3__1), .S0 (
             Instr)) ;
    mux21_ni ix893 (.Y (L1FirstOperands_0__2), .A0 (
             L1_2_L2_3_G2_MINI_ALU_BoothP_3), .A1 (WindowDin_2__3__2), .S0 (
             Instr)) ;
    mux21_ni ix901 (.Y (L1FirstOperands_0__3), .A0 (
             L1_2_L2_3_G2_MINI_ALU_BoothP_4), .A1 (WindowDin_2__3__3), .S0 (
             Instr)) ;
    mux21_ni ix909 (.Y (L1FirstOperands_0__4), .A0 (
             L1_2_L2_3_G2_MINI_ALU_BoothP_5), .A1 (WindowDin_2__3__4), .S0 (
             Instr)) ;
    mux21_ni ix917 (.Y (L1FirstOperands_0__5), .A0 (
             L1_2_L2_3_G2_MINI_ALU_BoothP_6), .A1 (WindowDin_2__3__5), .S0 (
             Instr)) ;
    mux21_ni ix925 (.Y (L1FirstOperands_0__6), .A0 (
             L1_2_L2_3_G2_MINI_ALU_BoothP_7), .A1 (WindowDin_2__3__6), .S0 (
             Instr)) ;
    mux21_ni ix933 (.Y (L1FirstOperands_0__7), .A0 (
             L1_2_L2_3_G2_MINI_ALU_BoothP_8), .A1 (WindowDin_2__3__7), .S0 (
             Instr)) ;
    nor02ii ix841 (.Y (L1FirstOperands_0__8), .A0 (Instr), .A1 (
            L1_2_L2_3_G2_MINI_ALU_BoothP_9)) ;
    nor02ii ix845 (.Y (L1FirstOperands_0__9), .A0 (Instr), .A1 (
            L1_2_L2_3_G2_MINI_ALU_BoothP_10)) ;
    nor02ii ix849 (.Y (L1FirstOperands_0__10), .A0 (Instr), .A1 (
            L1_2_L2_3_G2_MINI_ALU_BoothP_11)) ;
    nor02ii ix853 (.Y (L1FirstOperands_0__11), .A0 (Instr), .A1 (
            L1_2_L2_3_G2_MINI_ALU_BoothP_12)) ;
    nor02ii ix857 (.Y (L1FirstOperands_0__12), .A0 (Instr), .A1 (
            L1_2_L2_3_G2_MINI_ALU_BoothP_13)) ;
    nor02ii ix861 (.Y (L1FirstOperands_0__13), .A0 (Instr), .A1 (
            L1_2_L2_3_G2_MINI_ALU_BoothP_14)) ;
    nor02ii ix865 (.Y (L1FirstOperands_0__14), .A0 (Instr), .A1 (
            L1_2_L2_3_G2_MINI_ALU_BoothP_15)) ;
    nor02ii ix869 (.Y (L1FirstOperands_0__15), .A0 (Instr), .A1 (
            L1_2_L2_3_G2_MINI_ALU_BoothP_16)) ;
    nor02ii ix2243 (.Y (LoopingAndResultNotReady), .A0 (nx3230), .A1 (nx2853)) ;
    nor04 ix3231 (.Y (nx3230), .A0 (CounterOut_0), .A1 (CounterOut_1), .A2 (
          CounterOut_2), .A3 (CounterOut_3)) ;
    oai21 ix29 (.Y (Result[0]), .A0 (nx3233), .A1 (Instr), .B0 (nx3235)) ;
    inv01 ix3234 (.Y (nx3233), .A (L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_0)) ;
    aoi32 ix3236 (.Y (nx3235), .A0 (L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_5), .A1 (
          FilterSize), .A2 (Instr), .B0 (
          L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_3), .B1 (nx22)) ;
    nor02ii ix23 (.Y (nx22), .A0 (FilterSize), .A1 (Instr)) ;
    oai21 ix41 (.Y (Result[1]), .A0 (nx3239), .A1 (Instr), .B0 (nx3241)) ;
    inv01 ix3240 (.Y (nx3239), .A (L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_1)) ;
    aoi32 ix3242 (.Y (nx3241), .A0 (L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_6), .A1 (
          FilterSize), .A2 (Instr), .B0 (
          L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_4), .B1 (nx22)) ;
    oai21 ix53 (.Y (Result[2]), .A0 (nx3244), .A1 (Instr), .B0 (nx3246)) ;
    inv01 ix3245 (.Y (nx3244), .A (L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_2)) ;
    aoi32 ix3247 (.Y (nx3246), .A0 (L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_7), .A1 (
          FilterSize), .A2 (Instr), .B0 (
          L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_5), .B1 (nx22)) ;
    nor02ii ix3 (.Y (Result[5]), .A0 (Instr), .A1 (
            L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_5)) ;
    nor02ii ix7 (.Y (Result[6]), .A0 (Instr), .A1 (
            L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_6)) ;
    nor02ii ix11 (.Y (Result[7]), .A0 (Instr), .A1 (
            L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_7)) ;
    inv01 ix1079 (.Y (Done), .A (NOT__145383)) ;
    inv01 ix3269 (.Y (nx3270), .A (LoopingAndResultNotReady)) ;
    inv01 ix3271 (.Y (nx3272), .A (nx3270)) ;
    inv01 ix3273 (.Y (nx3274), .A (nx3270)) ;
    inv01 ix3275 (.Y (nx3276), .A (nx3270)) ;
    inv01 ix3277 (.Y (nx3278), .A (nx3270)) ;
    inv01 ix3279 (.Y (nx3280), .A (Done)) ;
    inv01 ix3281 (.Y (nx3282), .A (Done)) ;
    inv01 ix3283 (.Y (nx3284), .A (Done)) ;
    inv01 ix3285 (.Y (nx3286), .A (Done)) ;
    and02 ix1033 (.Y (nx1032), .A0 (NOT__145383), .A1 (CLK)) ;
    or02 ix2870 (.Y (nx2869), .A0 (nx2873), .A1 (NOT_CounterOut_0)) ;
    xnor2 ix1047 (.Y (nx1046), .A0 (nx2873), .A1 (CounterOut_0)) ;
    ao22 ix61 (.Y (Result[3]), .A0 (L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_6), .A1 (
         nx22), .B0 (L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_3), .B1 (nx3292)) ;
    inv01 ix3291 (.Y (nx3292), .A (Instr)) ;
    ao22 ix69 (.Y (Result[4]), .A0 (L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_7), .A1 (
         nx22), .B0 (L1_4_L2_4_G5_MINI_ALU_AdderResultLarge_4), .B1 (nx3292)) ;
endmodule


module booth_adder_17_unfolded17 ( AdderFirstOperand, AdderSecondOperand, 
                                   BoothOperand, BoothP, SelOperand, Operation, 
                                   AdderResult, AdderBoothResult ) ;

    input [16:0]AdderFirstOperand ;
    input [16:0]AdderSecondOperand ;
    input [16:0]BoothOperand ;
    input [16:0]BoothP ;
    input SelOperand ;
    input Operation ;
    output [16:0]AdderResult ;
    output [16:0]AdderBoothResult ;

    wire AdderResult_16_rename, AdderResult_15_rename, AdderResult_14_rename, 
         AdderResult_13_rename, AdderResult_12_rename, AdderResult_11_rename, 
         AdderResult_10_rename, AdderResult_9_rename, AdderResult_8_rename, 
         FirstOperand_16, FirstOperand_15, FirstOperand_14, FirstOperand_13, 
         FirstOperand_12, FirstOperand_11, FirstOperand_10, FirstOperand_9, 
         FirstOperand_8, FirstOperand_7, FirstOperand_6, FirstOperand_5, 
         FirstOperand_4, FirstOperand_3, FirstOperand_2, FirstOperand_1, 
         FirstOperand_0, SecondOperand_16, SecondOperand_15, SecondOperand_14, 
         SecondOperand_13, SecondOperand_12, SecondOperand_11, SecondOperand_10, 
         SecondOperand_9, SecondOperand_8, SecondOperand_7, SecondOperand_6, 
         SecondOperand_5, SecondOperand_4, SecondOperand_3, SecondOperand_2, 
         SecondOperand_1, SecondOperand_0, nx224, nx227, nx229, nx231, nx233, 
         nx235, nx237, nx239, nx241, nx243;
    wire [0:0] \$dummy ;




    assign AdderResult[16] = AdderBoothResult[16] ;
    assign AdderResult[15] = AdderBoothResult[16] ;
    assign AdderResult[14] = AdderBoothResult[16] ;
    assign AdderResult[13] = AdderBoothResult[16] ;
    assign AdderResult[12] = AdderBoothResult[16] ;
    assign AdderResult[11] = AdderBoothResult[16] ;
    assign AdderResult[10] = AdderBoothResult[16] ;
    assign AdderResult[9] = AdderBoothResult[16] ;
    assign AdderResult[8] = AdderBoothResult[16] ;
    adder_17 ADDER (.A ({FirstOperand_16,FirstOperand_15,FirstOperand_14,
             FirstOperand_13,FirstOperand_12,FirstOperand_11,FirstOperand_10,
             FirstOperand_9,FirstOperand_8,FirstOperand_7,FirstOperand_6,
             FirstOperand_5,FirstOperand_4,FirstOperand_3,FirstOperand_2,
             FirstOperand_1,FirstOperand_0}), .B ({SecondOperand_16,
             SecondOperand_15,SecondOperand_14,SecondOperand_13,SecondOperand_12
             ,SecondOperand_11,SecondOperand_10,SecondOperand_9,SecondOperand_8,
             SecondOperand_7,SecondOperand_6,SecondOperand_5,SecondOperand_4,
             SecondOperand_3,SecondOperand_2,SecondOperand_1,SecondOperand_0}), 
             .Cin (AdderBoothResult[16]), .Sum ({AdderResult_16_rename,
             AdderResult_15_rename,AdderResult_14_rename,AdderResult_13_rename,
             AdderResult_12_rename,AdderResult_11_rename,AdderResult_10_rename,
             AdderResult_9_rename,AdderResult_8_rename,AdderResult[7],
             AdderResult[6],AdderResult[5],AdderResult[4],AdderResult[3],
             AdderResult[2],AdderResult[1],AdderResult[0]}), .Cout (\$dummy [0])
             ) ;
    fake_gnd ix47 (.Y (AdderBoothResult[16])) ;
    mux21_ni ix137 (.Y (SecondOperand_0), .A0 (AdderSecondOperand[0]), .A1 (
             BoothP[0]), .S0 (nx235)) ;
    mux21_ni ix145 (.Y (SecondOperand_1), .A0 (AdderSecondOperand[1]), .A1 (
             BoothP[1]), .S0 (nx235)) ;
    mux21_ni ix153 (.Y (SecondOperand_2), .A0 (AdderSecondOperand[2]), .A1 (
             BoothP[2]), .S0 (nx235)) ;
    mux21_ni ix161 (.Y (SecondOperand_3), .A0 (AdderSecondOperand[3]), .A1 (
             BoothP[3]), .S0 (nx235)) ;
    mux21_ni ix169 (.Y (SecondOperand_4), .A0 (AdderSecondOperand[4]), .A1 (
             BoothP[4]), .S0 (nx235)) ;
    mux21_ni ix177 (.Y (SecondOperand_5), .A0 (AdderSecondOperand[5]), .A1 (
             BoothP[5]), .S0 (nx235)) ;
    mux21_ni ix185 (.Y (SecondOperand_6), .A0 (AdderSecondOperand[6]), .A1 (
             BoothP[6]), .S0 (nx235)) ;
    mux21_ni ix193 (.Y (SecondOperand_7), .A0 (AdderSecondOperand[7]), .A1 (
             BoothP[7]), .S0 (nx237)) ;
    mux21_ni ix201 (.Y (SecondOperand_8), .A0 (AdderSecondOperand[8]), .A1 (
             BoothP[8]), .S0 (nx237)) ;
    mux21_ni ix209 (.Y (SecondOperand_9), .A0 (AdderSecondOperand[9]), .A1 (
             BoothP[9]), .S0 (nx237)) ;
    mux21_ni ix217 (.Y (SecondOperand_10), .A0 (AdderSecondOperand[10]), .A1 (
             BoothP[10]), .S0 (nx237)) ;
    mux21_ni ix225 (.Y (SecondOperand_11), .A0 (AdderSecondOperand[11]), .A1 (
             BoothP[11]), .S0 (nx237)) ;
    mux21_ni ix233 (.Y (SecondOperand_12), .A0 (AdderSecondOperand[12]), .A1 (
             BoothP[12]), .S0 (nx237)) ;
    mux21_ni ix241 (.Y (SecondOperand_13), .A0 (AdderSecondOperand[13]), .A1 (
             BoothP[13]), .S0 (nx237)) ;
    mux21_ni ix249 (.Y (SecondOperand_14), .A0 (AdderSecondOperand[14]), .A1 (
             BoothP[14]), .S0 (nx239)) ;
    mux21_ni ix257 (.Y (SecondOperand_15), .A0 (AdderSecondOperand[15]), .A1 (
             BoothP[15]), .S0 (nx239)) ;
    nor02ii ix261 (.Y (FirstOperand_0), .A0 (nx239), .A1 (AdderFirstOperand[0])
            ) ;
    nor02ii ix265 (.Y (FirstOperand_1), .A0 (nx239), .A1 (AdderFirstOperand[1])
            ) ;
    nor02ii ix269 (.Y (FirstOperand_2), .A0 (nx239), .A1 (AdderFirstOperand[2])
            ) ;
    nor02ii ix273 (.Y (FirstOperand_3), .A0 (nx239), .A1 (AdderFirstOperand[3])
            ) ;
    nor02ii ix277 (.Y (FirstOperand_4), .A0 (nx239), .A1 (AdderFirstOperand[4])
            ) ;
    nor02ii ix281 (.Y (FirstOperand_5), .A0 (nx241), .A1 (AdderFirstOperand[5])
            ) ;
    nor02ii ix285 (.Y (FirstOperand_6), .A0 (nx241), .A1 (AdderFirstOperand[6])
            ) ;
    nor02ii ix289 (.Y (FirstOperand_7), .A0 (nx241), .A1 (AdderFirstOperand[7])
            ) ;
    nor02ii ix293 (.Y (FirstOperand_8), .A0 (nx241), .A1 (AdderFirstOperand[8])
            ) ;
    mux21_ni ix301 (.Y (FirstOperand_9), .A0 (AdderFirstOperand[9]), .A1 (
             BoothOperand[9]), .S0 (nx241)) ;
    mux21_ni ix309 (.Y (FirstOperand_10), .A0 (AdderFirstOperand[10]), .A1 (
             BoothOperand[10]), .S0 (nx241)) ;
    mux21_ni ix317 (.Y (FirstOperand_11), .A0 (AdderFirstOperand[11]), .A1 (
             BoothOperand[11]), .S0 (nx241)) ;
    mux21_ni ix325 (.Y (FirstOperand_12), .A0 (AdderFirstOperand[12]), .A1 (
             BoothOperand[12]), .S0 (nx243)) ;
    mux21_ni ix333 (.Y (FirstOperand_13), .A0 (AdderFirstOperand[13]), .A1 (
             BoothOperand[13]), .S0 (nx243)) ;
    mux21_ni ix341 (.Y (FirstOperand_14), .A0 (AdderFirstOperand[14]), .A1 (
             BoothOperand[14]), .S0 (nx243)) ;
    mux21_ni ix349 (.Y (FirstOperand_15), .A0 (AdderFirstOperand[15]), .A1 (
             BoothOperand[15]), .S0 (nx243)) ;
    mux21_ni ix357 (.Y (FirstOperand_16), .A0 (AdderFirstOperand[16]), .A1 (
             BoothOperand[16]), .S0 (nx243)) ;
    mux21_ni ix7 (.Y (AdderBoothResult[0]), .A0 (BoothP[1]), .A1 (AdderResult[1]
             ), .S0 (nx227)) ;
    mux21_ni ix15 (.Y (AdderBoothResult[1]), .A0 (BoothP[2]), .A1 (
             AdderResult[2]), .S0 (nx227)) ;
    mux21_ni ix23 (.Y (AdderBoothResult[2]), .A0 (BoothP[3]), .A1 (
             AdderResult[3]), .S0 (nx227)) ;
    mux21_ni ix31 (.Y (AdderBoothResult[3]), .A0 (BoothP[4]), .A1 (
             AdderResult[4]), .S0 (nx227)) ;
    mux21_ni ix39 (.Y (AdderBoothResult[4]), .A0 (BoothP[5]), .A1 (
             AdderResult[5]), .S0 (nx227)) ;
    mux21_ni ix49 (.Y (AdderBoothResult[5]), .A0 (BoothP[6]), .A1 (
             AdderResult[6]), .S0 (nx227)) ;
    mux21_ni ix55 (.Y (AdderBoothResult[6]), .A0 (BoothP[7]), .A1 (
             AdderResult[7]), .S0 (nx227)) ;
    mux21_ni ix63 (.Y (AdderBoothResult[7]), .A0 (BoothP[8]), .A1 (
             AdderResult_8_rename), .S0 (nx229)) ;
    mux21_ni ix71 (.Y (AdderBoothResult[8]), .A0 (BoothP[9]), .A1 (
             AdderResult_9_rename), .S0 (nx229)) ;
    mux21_ni ix79 (.Y (AdderBoothResult[9]), .A0 (BoothP[10]), .A1 (
             AdderResult_10_rename), .S0 (nx229)) ;
    mux21_ni ix87 (.Y (AdderBoothResult[10]), .A0 (BoothP[11]), .A1 (
             AdderResult_11_rename), .S0 (nx229)) ;
    mux21_ni ix95 (.Y (AdderBoothResult[11]), .A0 (BoothP[12]), .A1 (
             AdderResult_12_rename), .S0 (nx229)) ;
    mux21_ni ix103 (.Y (AdderBoothResult[12]), .A0 (BoothP[13]), .A1 (
             AdderResult_13_rename), .S0 (nx229)) ;
    mux21_ni ix111 (.Y (AdderBoothResult[13]), .A0 (BoothP[14]), .A1 (
             AdderResult_14_rename), .S0 (nx229)) ;
    mux21_ni ix119 (.Y (AdderBoothResult[14]), .A0 (BoothP[15]), .A1 (
             AdderResult_15_rename), .S0 (nx231)) ;
    mux21_ni ix127 (.Y (AdderBoothResult[15]), .A0 (BoothP[16]), .A1 (
             AdderResult_16_rename), .S0 (nx231)) ;
    and02 ix129 (.Y (SecondOperand_16), .A0 (nx243), .A1 (BoothP[16])) ;
    inv01 ix223 (.Y (nx224), .A (Operation)) ;
    inv02 ix226 (.Y (nx227), .A (nx224)) ;
    inv02 ix228 (.Y (nx229), .A (nx224)) ;
    inv02 ix230 (.Y (nx231), .A (nx224)) ;
    inv01 ix232 (.Y (nx233), .A (SelOperand)) ;
    inv02 ix234 (.Y (nx235), .A (nx233)) ;
    inv02 ix236 (.Y (nx237), .A (nx233)) ;
    inv02 ix238 (.Y (nx239), .A (nx233)) ;
    inv02 ix240 (.Y (nx241), .A (nx233)) ;
    inv02 ix242 (.Y (nx243), .A (nx233)) ;
endmodule


module booth_adder_17_unfolded16 ( AdderFirstOperand, AdderSecondOperand, 
                                   BoothOperand, BoothP, SelOperand, Operation, 
                                   AdderResult, AdderBoothResult ) ;

    input [16:0]AdderFirstOperand ;
    input [16:0]AdderSecondOperand ;
    input [16:0]BoothOperand ;
    input [16:0]BoothP ;
    input SelOperand ;
    input Operation ;
    output [16:0]AdderResult ;
    output [16:0]AdderBoothResult ;

    wire FirstOperand_16, FirstOperand_15, FirstOperand_14, FirstOperand_13, 
         FirstOperand_12, FirstOperand_11, FirstOperand_10, FirstOperand_9, 
         FirstOperand_8, FirstOperand_7, FirstOperand_6, FirstOperand_5, 
         FirstOperand_4, FirstOperand_3, FirstOperand_2, FirstOperand_1, 
         FirstOperand_0, SecondOperand_16, SecondOperand_15, SecondOperand_14, 
         SecondOperand_13, SecondOperand_12, SecondOperand_11, SecondOperand_10, 
         SecondOperand_9, SecondOperand_8, SecondOperand_7, SecondOperand_6, 
         SecondOperand_5, SecondOperand_4, SecondOperand_3, SecondOperand_2, 
         SecondOperand_1, SecondOperand_0, nx220, nx222, nx225, nx227, nx229, 
         nx231, nx233, nx235, nx237, nx239;
    wire [0:0] \$dummy ;




    adder_17 ADDER (.A ({FirstOperand_16,FirstOperand_15,FirstOperand_14,
             FirstOperand_13,FirstOperand_12,FirstOperand_11,FirstOperand_10,
             FirstOperand_9,FirstOperand_8,FirstOperand_7,FirstOperand_6,
             FirstOperand_5,FirstOperand_4,FirstOperand_3,FirstOperand_2,
             FirstOperand_1,FirstOperand_0}), .B ({SecondOperand_16,
             SecondOperand_15,SecondOperand_14,SecondOperand_13,SecondOperand_12
             ,SecondOperand_11,SecondOperand_10,SecondOperand_9,SecondOperand_8,
             SecondOperand_7,SecondOperand_6,SecondOperand_5,SecondOperand_4,
             SecondOperand_3,SecondOperand_2,SecondOperand_1,SecondOperand_0}), 
             .Cin (AdderBoothResult[16]), .Sum ({AdderResult[16],AdderResult[15]
             ,AdderResult[14],AdderResult[13],AdderResult[12],AdderResult[11],
             AdderResult[10],AdderResult[9],AdderResult[8],AdderResult[7],
             AdderResult[6],AdderResult[5],AdderResult[4],AdderResult[3],
             AdderResult[2],AdderResult[1],AdderResult[0]}), .Cout (\$dummy [0])
             ) ;
    fake_gnd ix45 (.Y (AdderBoothResult[16])) ;
    mux21_ni ix135 (.Y (SecondOperand_0), .A0 (AdderSecondOperand[0]), .A1 (
             BoothP[0]), .S0 (nx231)) ;
    mux21_ni ix143 (.Y (SecondOperand_1), .A0 (AdderSecondOperand[1]), .A1 (
             BoothP[1]), .S0 (nx231)) ;
    mux21_ni ix151 (.Y (SecondOperand_2), .A0 (AdderSecondOperand[2]), .A1 (
             BoothP[2]), .S0 (nx231)) ;
    mux21_ni ix159 (.Y (SecondOperand_3), .A0 (AdderSecondOperand[3]), .A1 (
             BoothP[3]), .S0 (nx231)) ;
    mux21_ni ix167 (.Y (SecondOperand_4), .A0 (AdderSecondOperand[4]), .A1 (
             BoothP[4]), .S0 (nx231)) ;
    mux21_ni ix175 (.Y (SecondOperand_5), .A0 (AdderSecondOperand[5]), .A1 (
             BoothP[5]), .S0 (nx231)) ;
    mux21_ni ix183 (.Y (SecondOperand_6), .A0 (AdderSecondOperand[6]), .A1 (
             BoothP[6]), .S0 (nx231)) ;
    mux21_ni ix191 (.Y (SecondOperand_7), .A0 (AdderSecondOperand[7]), .A1 (
             BoothP[7]), .S0 (nx233)) ;
    mux21_ni ix199 (.Y (SecondOperand_8), .A0 (AdderSecondOperand[8]), .A1 (
             BoothP[8]), .S0 (nx233)) ;
    mux21_ni ix207 (.Y (SecondOperand_9), .A0 (AdderSecondOperand[9]), .A1 (
             BoothP[9]), .S0 (nx233)) ;
    mux21_ni ix215 (.Y (SecondOperand_10), .A0 (AdderSecondOperand[10]), .A1 (
             BoothP[10]), .S0 (nx233)) ;
    mux21_ni ix223 (.Y (SecondOperand_11), .A0 (AdderSecondOperand[11]), .A1 (
             BoothP[11]), .S0 (nx233)) ;
    mux21_ni ix231 (.Y (SecondOperand_12), .A0 (AdderSecondOperand[12]), .A1 (
             BoothP[12]), .S0 (nx233)) ;
    mux21_ni ix239 (.Y (SecondOperand_13), .A0 (AdderSecondOperand[13]), .A1 (
             BoothP[13]), .S0 (nx233)) ;
    mux21_ni ix247 (.Y (SecondOperand_14), .A0 (AdderSecondOperand[14]), .A1 (
             BoothP[14]), .S0 (nx235)) ;
    mux21_ni ix255 (.Y (SecondOperand_15), .A0 (AdderSecondOperand[15]), .A1 (
             BoothP[15]), .S0 (nx235)) ;
    mux21_ni ix263 (.Y (SecondOperand_16), .A0 (AdderSecondOperand[16]), .A1 (
             BoothP[16]), .S0 (nx235)) ;
    nor02ii ix267 (.Y (FirstOperand_0), .A0 (nx235), .A1 (AdderFirstOperand[0])
            ) ;
    nor02ii ix271 (.Y (FirstOperand_1), .A0 (nx235), .A1 (AdderFirstOperand[1])
            ) ;
    nor02ii ix275 (.Y (FirstOperand_2), .A0 (nx235), .A1 (AdderFirstOperand[2])
            ) ;
    nor02ii ix279 (.Y (FirstOperand_3), .A0 (nx235), .A1 (AdderFirstOperand[3])
            ) ;
    nor02ii ix283 (.Y (FirstOperand_4), .A0 (nx237), .A1 (AdderFirstOperand[4])
            ) ;
    nor02ii ix287 (.Y (FirstOperand_5), .A0 (nx237), .A1 (AdderFirstOperand[5])
            ) ;
    nor02ii ix291 (.Y (FirstOperand_6), .A0 (nx237), .A1 (AdderFirstOperand[6])
            ) ;
    nor02ii ix295 (.Y (FirstOperand_7), .A0 (nx237), .A1 (AdderFirstOperand[7])
            ) ;
    nor02ii ix299 (.Y (FirstOperand_8), .A0 (nx237), .A1 (AdderFirstOperand[8])
            ) ;
    mux21_ni ix307 (.Y (FirstOperand_9), .A0 (AdderFirstOperand[9]), .A1 (
             BoothOperand[9]), .S0 (nx237)) ;
    mux21_ni ix315 (.Y (FirstOperand_10), .A0 (AdderFirstOperand[10]), .A1 (
             BoothOperand[10]), .S0 (nx237)) ;
    mux21_ni ix323 (.Y (FirstOperand_11), .A0 (AdderFirstOperand[11]), .A1 (
             BoothOperand[11]), .S0 (nx239)) ;
    mux21_ni ix331 (.Y (FirstOperand_12), .A0 (AdderFirstOperand[12]), .A1 (
             BoothOperand[12]), .S0 (nx239)) ;
    mux21_ni ix339 (.Y (FirstOperand_13), .A0 (AdderFirstOperand[13]), .A1 (
             BoothOperand[13]), .S0 (nx239)) ;
    mux21_ni ix347 (.Y (FirstOperand_14), .A0 (AdderFirstOperand[14]), .A1 (
             BoothOperand[14]), .S0 (nx239)) ;
    mux21_ni ix355 (.Y (FirstOperand_15), .A0 (AdderFirstOperand[15]), .A1 (
             BoothOperand[15]), .S0 (nx239)) ;
    mux21_ni ix363 (.Y (FirstOperand_16), .A0 (AdderFirstOperand[16]), .A1 (
             BoothOperand[16]), .S0 (nx239)) ;
    mux21_ni ix7 (.Y (AdderBoothResult[0]), .A0 (BoothP[1]), .A1 (AdderResult[1]
             ), .S0 (nx222)) ;
    mux21_ni ix15 (.Y (AdderBoothResult[1]), .A0 (BoothP[2]), .A1 (
             AdderResult[2]), .S0 (nx222)) ;
    mux21_ni ix23 (.Y (AdderBoothResult[2]), .A0 (BoothP[3]), .A1 (
             AdderResult[3]), .S0 (nx222)) ;
    mux21_ni ix31 (.Y (AdderBoothResult[3]), .A0 (BoothP[4]), .A1 (
             AdderResult[4]), .S0 (nx222)) ;
    mux21_ni ix39 (.Y (AdderBoothResult[4]), .A0 (BoothP[5]), .A1 (
             AdderResult[5]), .S0 (nx222)) ;
    mux21_ni ix48 (.Y (AdderBoothResult[5]), .A0 (BoothP[6]), .A1 (
             AdderResult[6]), .S0 (nx222)) ;
    mux21_ni ix55 (.Y (AdderBoothResult[6]), .A0 (BoothP[7]), .A1 (
             AdderResult[7]), .S0 (nx222)) ;
    mux21_ni ix63 (.Y (AdderBoothResult[7]), .A0 (BoothP[8]), .A1 (
             AdderResult[8]), .S0 (nx225)) ;
    mux21_ni ix71 (.Y (AdderBoothResult[8]), .A0 (BoothP[9]), .A1 (
             AdderResult[9]), .S0 (nx225)) ;
    mux21_ni ix79 (.Y (AdderBoothResult[9]), .A0 (BoothP[10]), .A1 (
             AdderResult[10]), .S0 (nx225)) ;
    mux21_ni ix87 (.Y (AdderBoothResult[10]), .A0 (BoothP[11]), .A1 (
             AdderResult[11]), .S0 (nx225)) ;
    mux21_ni ix95 (.Y (AdderBoothResult[11]), .A0 (BoothP[12]), .A1 (
             AdderResult[12]), .S0 (nx225)) ;
    mux21_ni ix103 (.Y (AdderBoothResult[12]), .A0 (BoothP[13]), .A1 (
             AdderResult[13]), .S0 (nx225)) ;
    mux21_ni ix111 (.Y (AdderBoothResult[13]), .A0 (BoothP[14]), .A1 (
             AdderResult[14]), .S0 (nx225)) ;
    mux21_ni ix119 (.Y (AdderBoothResult[14]), .A0 (BoothP[15]), .A1 (
             AdderResult[15]), .S0 (nx227)) ;
    mux21_ni ix127 (.Y (AdderBoothResult[15]), .A0 (BoothP[16]), .A1 (
             AdderResult[16]), .S0 (nx227)) ;
    inv01 ix219 (.Y (nx220), .A (Operation)) ;
    inv02 ix221 (.Y (nx222), .A (nx220)) ;
    inv02 ix224 (.Y (nx225), .A (nx220)) ;
    inv02 ix226 (.Y (nx227), .A (nx220)) ;
    inv01 ix228 (.Y (nx229), .A (SelOperand)) ;
    inv02 ix230 (.Y (nx231), .A (nx229)) ;
    inv02 ix232 (.Y (nx233), .A (nx229)) ;
    inv02 ix234 (.Y (nx235), .A (nx229)) ;
    inv02 ix236 (.Y (nx237), .A (nx229)) ;
    inv02 ix238 (.Y (nx239), .A (nx229)) ;
endmodule


module booth_unit_17_unfolded5 ( CLK, RST, Start, Instr, 
                                 LoopingAndResultNotReady, Filter, Window, 
                                 AdderBoothResult, BoothXORCheck, BoothResult, 
                                 BoothAddingOperand, BoothP, LargeWindowShifted
                                  ) ;

    input CLK ;
    input RST ;
    input Start ;
    input Instr ;
    input LoopingAndResultNotReady ;
    input [7:0]Filter ;
    input [7:0]Window ;
    input [16:0]AdderBoothResult ;
    output BoothXORCheck ;
    output [7:0]BoothResult ;
    output [16:0]BoothAddingOperand ;
    output [16:0]BoothP ;
    output [16:0]LargeWindowShifted ;

    wire BoothP_0_rename, RegisterPEN, RegisterPDin_16, RegisterPDin_15, 
         RegisterPDin_14, RegisterPDin_13, RegisterPDin_12, RegisterPDin_11, 
         RegisterPDin_10, RegisterPDin_9, RegisterPDin_8, RegisterPDin_7, 
         RegisterPDin_6, RegisterPDin_5, RegisterPDin_4, RegisterPDin_3, 
         RegisterPDin_2, RegisterPDin_1, RegisterPDin_0, RegisterSDout_10, nx12, 
         nx20, RegisterADout_10, RegisterSDout_11, nx52, nx60, RegisterADout_11, 
         RegisterSDout_12, nx92, nx100, RegisterADout_12, RegisterSDout_13, 
         nx132, nx140, RegisterADout_13, RegisterSDout_14, nx172, nx180, 
         RegisterADout_14, RegisterSDout_15, nx212, nx220, RegisterADout_15, 
         RegisterSDout_16, nx246, RegisterADout_16, nx69, nx79, nx89, nx99, 
         nx109, nx119, nx129, nx139, nx149, nx159, nx169, nx179, nx189, nx199, 
         nx209, nx224, nx226, nx235, nx249, nx261, nx273, nx286, nx299, nx315, 
         nx324, nx326, nx328;
    wire [14:0] \$dummy ;




    assign BoothResult[7] = LargeWindowShifted[16] ;
    assign BoothResult[6] = LargeWindowShifted[16] ;
    assign BoothResult[5] = LargeWindowShifted[16] ;
    assign BoothResult[4] = LargeWindowShifted[16] ;
    assign BoothResult[3] = LargeWindowShifted[16] ;
    assign BoothResult[2] = LargeWindowShifted[16] ;
    assign BoothResult[1] = LargeWindowShifted[16] ;
    assign BoothResult[0] = LargeWindowShifted[16] ;
    assign BoothAddingOperand[8] = LargeWindowShifted[16] ;
    assign BoothAddingOperand[7] = LargeWindowShifted[16] ;
    assign BoothAddingOperand[6] = LargeWindowShifted[16] ;
    assign BoothAddingOperand[5] = LargeWindowShifted[16] ;
    assign BoothAddingOperand[4] = LargeWindowShifted[16] ;
    assign BoothAddingOperand[3] = LargeWindowShifted[16] ;
    assign BoothAddingOperand[2] = LargeWindowShifted[16] ;
    assign BoothAddingOperand[1] = LargeWindowShifted[16] ;
    assign BoothAddingOperand[0] = LargeWindowShifted[16] ;
    assign BoothP[0] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[15] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[14] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[13] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[12] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[11] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[10] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[9] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[8] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[7] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[6] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[5] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[4] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[3] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[2] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[1] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[0] = LargeWindowShifted[16] ;
    register_edge_rising_17 REGISTER_P (.CLK (CLK), .RST (RST), .EN (RegisterPEN), .Din (
                     {RegisterPDin_16,RegisterPDin_15,RegisterPDin_14,
                     RegisterPDin_13,RegisterPDin_12,RegisterPDin_11,
                     RegisterPDin_10,RegisterPDin_9,RegisterPDin_8,
                     RegisterPDin_7,RegisterPDin_6,RegisterPDin_5,RegisterPDin_4
                     ,RegisterPDin_3,RegisterPDin_2,RegisterPDin_1,
                     RegisterPDin_0}), .Dout ({BoothP[16],BoothP[15],BoothP[14],
                     BoothP[13],BoothP[12],BoothP[11],BoothP[10],BoothP[9],
                     BoothP[8],BoothP[7],BoothP[6],BoothP[5],BoothP[4],BoothP[3]
                     ,BoothP[2],BoothP[1],BoothP_0_rename})) ;
    mux_4x1_17 P_INPUT_DATA_MUX (.A ({LargeWindowShifted[16],
               AdderBoothResult[15],AdderBoothResult[14],AdderBoothResult[13],
               AdderBoothResult[12],AdderBoothResult[11],AdderBoothResult[10],
               AdderBoothResult[9],AdderBoothResult[8],AdderBoothResult[7],
               AdderBoothResult[6],AdderBoothResult[5],AdderBoothResult[4],
               AdderBoothResult[3],AdderBoothResult[2],AdderBoothResult[1],
               AdderBoothResult[0]}), .B ({LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16]}), .C ({
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],Window[7],Window[6]
               ,Window[5],Window[4],Window[3],Window[2],Window[1],Window[0],
               LargeWindowShifted[16]}), .D ({LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16]}), .S ({Start,Instr
               }), .Dout ({RegisterPDin_16,RegisterPDin_15,RegisterPDin_14,
               RegisterPDin_13,RegisterPDin_12,RegisterPDin_11,RegisterPDin_10,
               RegisterPDin_9,RegisterPDin_8,RegisterPDin_7,RegisterPDin_6,
               RegisterPDin_5,RegisterPDin_4,RegisterPDin_3,RegisterPDin_2,
               RegisterPDin_1,RegisterPDin_0})) ;
    fake_gnd ix43 (.Y (LargeWindowShifted[16])) ;
    dff REGISTER_A_reg_Dout_9 (.Q (BoothAddingOperand[9]), .QB (\$dummy [0]), .D (
        nx209), .CLK (CLK)) ;
    ao32 ix210 (.Y (nx209), .A0 (nx324), .A1 (Filter[0]), .A2 (Start), .B0 (
         BoothAddingOperand[9]), .B1 (nx326)) ;
    inv01 ix225 (.Y (nx224), .A (RST)) ;
    nor02_2x ix227 (.Y (nx226), .A0 (Start), .A1 (RST)) ;
    or02 ix287 (.Y (RegisterPEN), .A0 (Start), .A1 (LoopingAndResultNotReady)) ;
    dff REGISTER_S_reg_Dout_10 (.Q (RegisterSDout_10), .QB (\$dummy [1]), .D (
        nx69), .CLK (CLK)) ;
    mux21_ni ix70 (.Y (nx69), .A0 (nx20), .A1 (RegisterSDout_10), .S0 (nx326)) ;
    aoi21 ix21 (.Y (nx20), .A0 (Filter[1]), .A1 (Filter[0]), .B0 (nx235)) ;
    or02 ix236 (.Y (nx235), .A0 (RST), .A1 (nx12)) ;
    nor02_2x ix13 (.Y (nx12), .A0 (Filter[0]), .A1 (Filter[1])) ;
    dff REGISTER_A_reg_Dout_10 (.Q (RegisterADout_10), .QB (\$dummy [2]), .D (
        nx79), .CLK (CLK)) ;
    ao32 ix80 (.Y (nx79), .A0 (nx324), .A1 (Filter[1]), .A2 (Start), .B0 (
         RegisterADout_10), .B1 (nx326)) ;
    dff REGISTER_S_reg_Dout_11 (.Q (RegisterSDout_11), .QB (\$dummy [3]), .D (
        nx89), .CLK (CLK)) ;
    mux21_ni ix90 (.Y (nx89), .A0 (nx60), .A1 (RegisterSDout_11), .S0 (nx326)) ;
    nor03_2x ix61 (.Y (nx60), .A0 (nx249), .A1 (RST), .A2 (nx52)) ;
    nor02ii ix250 (.Y (nx249), .A0 (nx12), .A1 (Filter[2])) ;
    nor03_2x ix53 (.Y (nx52), .A0 (Filter[2]), .A1 (Filter[0]), .A2 (Filter[1])
             ) ;
    dff REGISTER_A_reg_Dout_11 (.Q (RegisterADout_11), .QB (\$dummy [4]), .D (
        nx99), .CLK (CLK)) ;
    ao32 ix100 (.Y (nx99), .A0 (nx324), .A1 (Filter[2]), .A2 (Start), .B0 (
         RegisterADout_11), .B1 (nx326)) ;
    dff REGISTER_S_reg_Dout_12 (.Q (RegisterSDout_12), .QB (\$dummy [5]), .D (
        nx109), .CLK (CLK)) ;
    mux21_ni ix110 (.Y (nx109), .A0 (nx100), .A1 (RegisterSDout_12), .S0 (nx326)
             ) ;
    nor03_2x ix101 (.Y (nx100), .A0 (nx261), .A1 (RST), .A2 (nx92)) ;
    nor02ii ix262 (.Y (nx261), .A0 (nx52), .A1 (Filter[3])) ;
    nor04 ix93 (.Y (nx92), .A0 (Filter[3]), .A1 (Filter[2]), .A2 (Filter[0]), .A3 (
          Filter[1])) ;
    dff REGISTER_A_reg_Dout_12 (.Q (RegisterADout_12), .QB (\$dummy [6]), .D (
        nx119), .CLK (CLK)) ;
    ao32 ix120 (.Y (nx119), .A0 (nx324), .A1 (Filter[3]), .A2 (Start), .B0 (
         RegisterADout_12), .B1 (nx326)) ;
    dff REGISTER_S_reg_Dout_13 (.Q (RegisterSDout_13), .QB (\$dummy [7]), .D (
        nx129), .CLK (CLK)) ;
    mux21_ni ix130 (.Y (nx129), .A0 (nx140), .A1 (RegisterSDout_13), .S0 (nx328)
             ) ;
    nor03_2x ix141 (.Y (nx140), .A0 (nx273), .A1 (RST), .A2 (nx132)) ;
    nor02ii ix274 (.Y (nx273), .A0 (nx92), .A1 (Filter[4])) ;
    nor02ii ix133 (.Y (nx132), .A0 (Filter[4]), .A1 (nx92)) ;
    dff REGISTER_A_reg_Dout_13 (.Q (RegisterADout_13), .QB (\$dummy [8]), .D (
        nx139), .CLK (CLK)) ;
    ao32 ix140 (.Y (nx139), .A0 (nx324), .A1 (Filter[4]), .A2 (Start), .B0 (
         RegisterADout_13), .B1 (nx328)) ;
    dff REGISTER_S_reg_Dout_14 (.Q (RegisterSDout_14), .QB (\$dummy [9]), .D (
        nx149), .CLK (CLK)) ;
    mux21_ni ix150 (.Y (nx149), .A0 (nx180), .A1 (RegisterSDout_14), .S0 (nx328)
             ) ;
    nor03_2x ix181 (.Y (nx180), .A0 (nx286), .A1 (RST), .A2 (nx172)) ;
    nor02ii ix288 (.Y (nx286), .A0 (nx132), .A1 (Filter[5])) ;
    nor02ii ix173 (.Y (nx172), .A0 (Filter[5]), .A1 (nx132)) ;
    dff REGISTER_A_reg_Dout_14 (.Q (RegisterADout_14), .QB (\$dummy [10]), .D (
        nx159), .CLK (CLK)) ;
    ao32 ix160 (.Y (nx159), .A0 (nx324), .A1 (Filter[5]), .A2 (Start), .B0 (
         RegisterADout_14), .B1 (nx328)) ;
    dff REGISTER_S_reg_Dout_15 (.Q (RegisterSDout_15), .QB (\$dummy [11]), .D (
        nx169), .CLK (CLK)) ;
    mux21_ni ix170 (.Y (nx169), .A0 (nx220), .A1 (RegisterSDout_15), .S0 (nx328)
             ) ;
    nor03_2x ix221 (.Y (nx220), .A0 (nx299), .A1 (RST), .A2 (nx212)) ;
    nor02ii ix300 (.Y (nx299), .A0 (nx172), .A1 (Filter[6])) ;
    nor02ii ix213 (.Y (nx212), .A0 (Filter[6]), .A1 (nx172)) ;
    dff REGISTER_A_reg_Dout_15 (.Q (RegisterADout_15), .QB (\$dummy [12]), .D (
        nx179), .CLK (CLK)) ;
    ao32 ix180 (.Y (nx179), .A0 (nx324), .A1 (Filter[6]), .A2 (Start), .B0 (
         RegisterADout_15), .B1 (nx328)) ;
    dff REGISTER_S_reg_Dout_16 (.Q (RegisterSDout_16), .QB (\$dummy [13]), .D (
        nx189), .CLK (CLK)) ;
    ao32 ix190 (.Y (nx189), .A0 (nx224), .A1 (nx246), .A2 (Start), .B0 (
         RegisterSDout_16), .B1 (nx328)) ;
    xnor2 ix247 (.Y (nx246), .A0 (Filter[7]), .A1 (nx212)) ;
    dff REGISTER_A_reg_Dout_16 (.Q (RegisterADout_16), .QB (\$dummy [14]), .D (
        nx199), .CLK (CLK)) ;
    ao32 ix200 (.Y (nx199), .A0 (nx224), .A1 (Filter[7]), .A2 (Start), .B0 (
         RegisterADout_16), .B1 (nx226)) ;
    inv02 ix316 (.Y (nx315), .A (BoothP_0_rename)) ;
    inv01 ix323 (.Y (nx324), .A (RST)) ;
    nor02_2x ix325 (.Y (nx326), .A0 (Start), .A1 (RST)) ;
    nor02_2x ix327 (.Y (nx328), .A0 (Start), .A1 (RST)) ;
    mux21_ni ix46 (.Y (BoothAddingOperand[10]), .A0 (RegisterADout_10), .A1 (
             RegisterSDout_10), .S0 (nx315)) ;
    mux21_ni ix85 (.Y (BoothAddingOperand[11]), .A0 (RegisterADout_11), .A1 (
             RegisterSDout_11), .S0 (nx315)) ;
    mux21_ni ix125 (.Y (BoothAddingOperand[12]), .A0 (RegisterADout_12), .A1 (
             RegisterSDout_12), .S0 (nx315)) ;
    mux21_ni ix165 (.Y (BoothAddingOperand[13]), .A0 (RegisterADout_13), .A1 (
             RegisterSDout_13), .S0 (nx315)) ;
    mux21_ni ix205 (.Y (BoothAddingOperand[14]), .A0 (RegisterADout_14), .A1 (
             RegisterSDout_14), .S0 (nx315)) ;
    mux21_ni ix245 (.Y (BoothAddingOperand[15]), .A0 (RegisterADout_15), .A1 (
             RegisterSDout_15), .S0 (nx315)) ;
    mux21_ni ix275 (.Y (BoothAddingOperand[16]), .A0 (RegisterADout_16), .A1 (
             RegisterSDout_16), .S0 (nx315)) ;
    xor2 ix289 (.Y (BoothXORCheck), .A0 (BoothP[1]), .A1 (BoothP_0_rename)) ;
endmodule


module booth_adder_17_unfolded15 ( AdderFirstOperand, AdderSecondOperand, 
                                   BoothOperand, BoothP, SelOperand, Operation, 
                                   AdderResult, AdderBoothResult ) ;

    input [16:0]AdderFirstOperand ;
    input [16:0]AdderSecondOperand ;
    input [16:0]BoothOperand ;
    input [16:0]BoothP ;
    input SelOperand ;
    input Operation ;
    output [16:0]AdderResult ;
    output [16:0]AdderBoothResult ;

    wire AdderResult_16_rename, AdderResult_15_rename, AdderResult_14_rename, 
         AdderResult_13_rename, AdderResult_12_rename, AdderResult_11_rename, 
         AdderResult_10_rename, AdderResult_9_rename, FirstOperand_16, 
         FirstOperand_15, FirstOperand_14, FirstOperand_13, FirstOperand_12, 
         FirstOperand_11, FirstOperand_10, FirstOperand_9, SecondOperand_16, 
         SecondOperand_15, SecondOperand_14, SecondOperand_13, SecondOperand_12, 
         SecondOperand_11, SecondOperand_10, SecondOperand_9, SecondOperand_8, 
         SecondOperand_7, SecondOperand_6, SecondOperand_5, SecondOperand_4, 
         nx143, nx153, nx155, nx158, nx161, nx164, nx167, nx182, nx184, nx186, 
         nx188, nx190, nx192, nx194;
    wire [9:0] \$dummy ;




    assign AdderResult[16] = AdderBoothResult[16] ;
    assign AdderResult[15] = AdderBoothResult[16] ;
    assign AdderResult[14] = AdderBoothResult[16] ;
    assign AdderResult[13] = AdderBoothResult[16] ;
    assign AdderResult[12] = AdderBoothResult[16] ;
    assign AdderResult[11] = AdderBoothResult[16] ;
    assign AdderResult[10] = AdderBoothResult[16] ;
    assign AdderResult[9] = AdderBoothResult[16] ;
    assign AdderResult[8] = AdderBoothResult[16] ;
    assign AdderResult[7] = AdderBoothResult[16] ;
    assign AdderResult[6] = AdderBoothResult[16] ;
    assign AdderResult[5] = AdderBoothResult[16] ;
    assign AdderResult[4] = AdderBoothResult[16] ;
    assign AdderResult[3] = AdderBoothResult[16] ;
    assign AdderResult[2] = AdderBoothResult[16] ;
    assign AdderResult[1] = AdderBoothResult[16] ;
    assign AdderResult[0] = AdderBoothResult[16] ;
    adder_17_unfolded5 ADDER (.A ({FirstOperand_16,FirstOperand_15,
                       FirstOperand_14,FirstOperand_13,FirstOperand_12,
                       FirstOperand_11,FirstOperand_10,FirstOperand_9,
                       AdderBoothResult[16],AdderBoothResult[16],
                       AdderBoothResult[16],AdderBoothResult[16],
                       AdderBoothResult[16],AdderBoothResult[16],
                       AdderBoothResult[16],AdderBoothResult[16],
                       AdderBoothResult[16]}), .B ({SecondOperand_16,
                       SecondOperand_15,SecondOperand_14,SecondOperand_13,
                       SecondOperand_12,SecondOperand_11,SecondOperand_10,
                       SecondOperand_9,SecondOperand_8,SecondOperand_7,
                       SecondOperand_6,SecondOperand_5,SecondOperand_4,
                       AdderBoothResult[16],AdderBoothResult[16],
                       AdderBoothResult[16],AdderBoothResult[16]}), .Cin (
                       AdderBoothResult[16]), .Sum ({AdderResult_16_rename,
                       AdderResult_15_rename,AdderResult_14_rename,
                       AdderResult_13_rename,AdderResult_12_rename,
                       AdderResult_11_rename,AdderResult_10_rename,
                       AdderResult_9_rename,\$dummy [0],\$dummy [1],\$dummy [2],
                       \$dummy [3],\$dummy [4],\$dummy [5],\$dummy [6],
                       \$dummy [7],\$dummy [8]}), .Cout (\$dummy [9])) ;
    fake_gnd ix59 (.Y (AdderBoothResult[16])) ;
    and02 ix15 (.Y (SecondOperand_4), .A0 (BoothP[4]), .A1 (nx186)) ;
    and02 ix25 (.Y (SecondOperand_5), .A0 (BoothP[5]), .A1 (nx186)) ;
    and02 ix35 (.Y (SecondOperand_6), .A0 (BoothP[6]), .A1 (nx186)) ;
    and02 ix45 (.Y (SecondOperand_7), .A0 (BoothP[7]), .A1 (nx186)) ;
    and02 ix55 (.Y (SecondOperand_8), .A0 (BoothP[8]), .A1 (nx186)) ;
    and02 ix125 (.Y (SecondOperand_9), .A0 (BoothP[9]), .A1 (nx186)) ;
    and02 ix127 (.Y (SecondOperand_10), .A0 (BoothP[10]), .A1 (nx186)) ;
    and02 ix129 (.Y (SecondOperand_11), .A0 (BoothP[11]), .A1 (nx188)) ;
    and02 ix131 (.Y (SecondOperand_12), .A0 (BoothP[12]), .A1 (nx188)) ;
    and02 ix133 (.Y (SecondOperand_13), .A0 (BoothP[13]), .A1 (nx188)) ;
    and02 ix135 (.Y (SecondOperand_14), .A0 (BoothP[14]), .A1 (nx188)) ;
    and02 ix137 (.Y (SecondOperand_15), .A0 (BoothP[15]), .A1 (nx188)) ;
    and02 ix139 (.Y (SecondOperand_16), .A0 (BoothP[16]), .A1 (nx188)) ;
    and02 ix141 (.Y (FirstOperand_9), .A0 (BoothOperand[9]), .A1 (nx188)) ;
    and02 ix143 (.Y (FirstOperand_10), .A0 (BoothOperand[10]), .A1 (nx190)) ;
    and02 ix145 (.Y (FirstOperand_11), .A0 (BoothOperand[11]), .A1 (nx190)) ;
    and02 ix147 (.Y (FirstOperand_12), .A0 (BoothOperand[12]), .A1 (nx190)) ;
    and02 ix149 (.Y (FirstOperand_13), .A0 (BoothOperand[13]), .A1 (nx190)) ;
    and02 ix151 (.Y (FirstOperand_14), .A0 (BoothOperand[14]), .A1 (nx190)) ;
    and02 ix153 (.Y (FirstOperand_15), .A0 (BoothOperand[15]), .A1 (nx190)) ;
    and02 ix155 (.Y (FirstOperand_16), .A0 (nx190), .A1 (BoothOperand[16])) ;
    nor02ii ix5 (.Y (AdderBoothResult[0]), .A0 (nx143), .A1 (BoothP[1])) ;
    nor02ii ix7 (.Y (AdderBoothResult[1]), .A0 (nx143), .A1 (BoothP[2])) ;
    nor02ii ix9 (.Y (AdderBoothResult[2]), .A0 (nx143), .A1 (BoothP[3])) ;
    aoi21 ix19 (.Y (AdderBoothResult[3]), .A0 (nx182), .A1 (nx194), .B0 (nx155)
          ) ;
    inv01 ix154 (.Y (nx153), .A (SelOperand)) ;
    inv01 ix156 (.Y (nx155), .A (BoothP[4])) ;
    aoi21 ix29 (.Y (AdderBoothResult[4]), .A0 (nx182), .A1 (nx194), .B0 (nx158)
          ) ;
    inv01 ix159 (.Y (nx158), .A (BoothP[5])) ;
    aoi21 ix39 (.Y (AdderBoothResult[5]), .A0 (nx182), .A1 (nx194), .B0 (nx161)
          ) ;
    inv01 ix162 (.Y (nx161), .A (BoothP[6])) ;
    aoi21 ix49 (.Y (AdderBoothResult[6]), .A0 (nx182), .A1 (nx194), .B0 (nx164)
          ) ;
    inv01 ix165 (.Y (nx164), .A (BoothP[7])) ;
    aoi21 ix61 (.Y (AdderBoothResult[7]), .A0 (nx182), .A1 (nx194), .B0 (nx167)
          ) ;
    inv01 ix168 (.Y (nx167), .A (BoothP[8])) ;
    mux21_ni ix67 (.Y (AdderBoothResult[8]), .A0 (BoothP[9]), .A1 (
             AdderResult_9_rename), .S0 (nx182)) ;
    mux21_ni ix75 (.Y (AdderBoothResult[9]), .A0 (BoothP[10]), .A1 (
             AdderResult_10_rename), .S0 (nx182)) ;
    mux21_ni ix83 (.Y (AdderBoothResult[10]), .A0 (BoothP[11]), .A1 (
             AdderResult_11_rename), .S0 (nx184)) ;
    mux21_ni ix91 (.Y (AdderBoothResult[11]), .A0 (BoothP[12]), .A1 (
             AdderResult_12_rename), .S0 (nx184)) ;
    mux21_ni ix99 (.Y (AdderBoothResult[12]), .A0 (BoothP[13]), .A1 (
             AdderResult_13_rename), .S0 (nx184)) ;
    mux21_ni ix107 (.Y (AdderBoothResult[13]), .A0 (BoothP[14]), .A1 (
             AdderResult_14_rename), .S0 (nx184)) ;
    mux21_ni ix115 (.Y (AdderBoothResult[14]), .A0 (BoothP[15]), .A1 (
             AdderResult_15_rename), .S0 (nx184)) ;
    mux21_ni ix123 (.Y (AdderBoothResult[15]), .A0 (BoothP[16]), .A1 (
             AdderResult_16_rename), .S0 (nx184)) ;
    nor02ii ix144 (.Y (nx143), .A0 (nx192), .A1 (nx184)) ;
    buf02 ix181 (.Y (nx182), .A (Operation)) ;
    buf02 ix183 (.Y (nx184), .A (Operation)) ;
    inv02 ix185 (.Y (nx186), .A (nx194)) ;
    inv02 ix187 (.Y (nx188), .A (nx153)) ;
    inv02 ix189 (.Y (nx190), .A (nx153)) ;
    inv02 ix191 (.Y (nx192), .A (nx153)) ;
    inv01 ix193 (.Y (nx194), .A (SelOperand)) ;
endmodule


module adder_17_unfolded5 ( A, B, Cin, Sum, Cout ) ;

    input [16:0]A ;
    input [16:0]B ;
    input Cin ;
    output [16:0]Sum ;
    output Cout ;

    wire nx2, nx16, nx18, nx32, nx34, nx48, nx93, nx95, nx98, nx101, nx105, 
         nx107, nx110, nx113, nx117, nx119, nx122, nx125, nx129, nx131;



    assign Sum[8] = B[8] ;
    assign Sum[7] = B[7] ;
    assign Sum[6] = B[6] ;
    assign Sum[5] = B[5] ;
    assign Sum[4] = B[4] ;
    assign Sum[3] = Cout ;
    assign Sum[2] = Cout ;
    assign Sum[1] = Cout ;
    assign Sum[0] = Cout ;
    fake_gnd ix68 (.Y (Cout)) ;
    xor2 ix71 (.Y (Sum[9]), .A0 (B[9]), .A1 (A[9])) ;
    xor2 ix65 (.Y (Sum[10]), .A0 (nx93), .A1 (nx95)) ;
    nand02 ix94 (.Y (nx93), .A0 (B[9]), .A1 (A[9])) ;
    xnor2 ix96 (.Y (nx95), .A0 (A[10]), .A1 (B[10])) ;
    xor2 ix63 (.Y (Sum[11]), .A0 (nx98), .A1 (nx101)) ;
    aoi32 ix99 (.Y (nx98), .A0 (B[9]), .A1 (A[9]), .A2 (nx2), .B0 (B[10]), .B1 (
          A[10])) ;
    xnor2 ix102 (.Y (nx101), .A0 (A[11]), .A1 (B[11])) ;
    xnor2 ix61 (.Y (Sum[12]), .A0 (nx16), .A1 (nx107)) ;
    oai21 ix17 (.Y (nx16), .A0 (nx98), .A1 (nx101), .B0 (nx105)) ;
    nand02 ix106 (.Y (nx105), .A0 (B[11]), .A1 (A[11])) ;
    xnor2 ix108 (.Y (nx107), .A0 (A[12]), .A1 (B[12])) ;
    xor2 ix59 (.Y (Sum[13]), .A0 (nx110), .A1 (nx113)) ;
    aoi22 ix111 (.Y (nx110), .A0 (B[12]), .A1 (A[12]), .B0 (nx16), .B1 (nx18)) ;
    xnor2 ix114 (.Y (nx113), .A0 (A[13]), .A1 (B[13])) ;
    xnor2 ix57 (.Y (Sum[14]), .A0 (nx32), .A1 (nx119)) ;
    oai21 ix33 (.Y (nx32), .A0 (nx110), .A1 (nx113), .B0 (nx117)) ;
    nand02 ix118 (.Y (nx117), .A0 (B[13]), .A1 (A[13])) ;
    xnor2 ix120 (.Y (nx119), .A0 (A[14]), .A1 (B[14])) ;
    xor2 ix55 (.Y (Sum[15]), .A0 (nx122), .A1 (nx125)) ;
    aoi22 ix123 (.Y (nx122), .A0 (B[14]), .A1 (A[14]), .B0 (nx32), .B1 (nx34)) ;
    xnor2 ix126 (.Y (nx125), .A0 (A[15]), .A1 (B[15])) ;
    xnor2 ix53 (.Y (Sum[16]), .A0 (nx48), .A1 (nx131)) ;
    oai21 ix49 (.Y (nx48), .A0 (nx122), .A1 (nx125), .B0 (nx129)) ;
    nand02 ix130 (.Y (nx129), .A0 (B[15]), .A1 (A[15])) ;
    xnor2 ix132 (.Y (nx131), .A0 (A[16]), .A1 (B[16])) ;
    inv01 ix35 (.Y (nx34), .A (nx119)) ;
    inv01 ix19 (.Y (nx18), .A (nx107)) ;
    inv01 ix3 (.Y (nx2), .A (nx95)) ;
endmodule


module booth_unit_17 ( CLK, RST, Start, Instr, LoopingAndResultNotReady, Filter, 
                       Window, AdderBoothResult, BoothXORCheck, BoothResult, 
                       BoothAddingOperand, BoothP, LargeWindowShifted ) ;

    input CLK ;
    input RST ;
    input Start ;
    input Instr ;
    input LoopingAndResultNotReady ;
    input [7:0]Filter ;
    input [7:0]Window ;
    input [16:0]AdderBoothResult ;
    output BoothXORCheck ;
    output [7:0]BoothResult ;
    output [16:0]BoothAddingOperand ;
    output [16:0]BoothP ;
    output [16:0]LargeWindowShifted ;

    wire RegisterPEN, RegisterPDin_16, RegisterPDin_15, RegisterPDin_14, 
         RegisterPDin_13, RegisterPDin_12, RegisterPDin_11, RegisterPDin_10, 
         RegisterPDin_9, RegisterPDin_8, RegisterPDin_7, RegisterPDin_6, 
         RegisterPDin_5, RegisterPDin_4, RegisterPDin_3, RegisterPDin_2, 
         RegisterPDin_1, RegisterPDin_0, RegisterSDout_10, nx12, nx20, 
         RegisterADout_10, RegisterSDout_11, nx52, nx60, RegisterADout_11, 
         RegisterSDout_12, nx92, nx100, RegisterADout_12, RegisterSDout_13, 
         nx132, nx140, RegisterADout_13, RegisterSDout_14, nx172, nx180, 
         RegisterADout_14, RegisterSDout_15, nx212, nx220, RegisterADout_15, 
         RegisterSDout_16, nx246, RegisterADout_16, nx69, nx79, nx89, nx99, 
         nx109, nx119, nx129, nx139, nx149, nx159, nx169, nx179, nx189, nx199, 
         nx209, nx224, nx226, nx235, nx249, nx261, nx273, nx286, nx299, nx320, 
         nx322, nx324, nx326, nx328;
    wire [14:0] \$dummy ;




    assign BoothResult[7] = LargeWindowShifted[16] ;
    assign BoothResult[6] = LargeWindowShifted[16] ;
    assign BoothResult[5] = LargeWindowShifted[16] ;
    assign BoothResult[4] = LargeWindowShifted[16] ;
    assign BoothResult[3] = LargeWindowShifted[16] ;
    assign BoothResult[2] = LargeWindowShifted[16] ;
    assign BoothResult[1] = LargeWindowShifted[16] ;
    assign BoothResult[0] = LargeWindowShifted[16] ;
    assign BoothAddingOperand[8] = LargeWindowShifted[16] ;
    assign BoothAddingOperand[7] = LargeWindowShifted[16] ;
    assign BoothAddingOperand[6] = LargeWindowShifted[16] ;
    assign BoothAddingOperand[5] = LargeWindowShifted[16] ;
    assign BoothAddingOperand[4] = LargeWindowShifted[16] ;
    assign BoothAddingOperand[3] = LargeWindowShifted[16] ;
    assign BoothAddingOperand[2] = LargeWindowShifted[16] ;
    assign BoothAddingOperand[1] = LargeWindowShifted[16] ;
    assign BoothAddingOperand[0] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[15] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[14] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[13] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[12] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[11] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[10] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[9] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[8] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[7] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[6] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[5] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[4] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[3] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[2] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[1] = LargeWindowShifted[16] ;
    assign LargeWindowShifted[0] = LargeWindowShifted[16] ;
    register_edge_rising_17 REGISTER_P (.CLK (CLK), .RST (RST), .EN (RegisterPEN), .Din (
                     {RegisterPDin_16,RegisterPDin_15,RegisterPDin_14,
                     RegisterPDin_13,RegisterPDin_12,RegisterPDin_11,
                     RegisterPDin_10,RegisterPDin_9,RegisterPDin_8,
                     RegisterPDin_7,RegisterPDin_6,RegisterPDin_5,RegisterPDin_4
                     ,RegisterPDin_3,RegisterPDin_2,RegisterPDin_1,
                     RegisterPDin_0}), .Dout ({BoothP[16],BoothP[15],BoothP[14],
                     BoothP[13],BoothP[12],BoothP[11],BoothP[10],BoothP[9],
                     BoothP[8],BoothP[7],BoothP[6],BoothP[5],BoothP[4],BoothP[3]
                     ,BoothP[2],BoothP[1],BoothP[0]})) ;
    mux_4x1_17 P_INPUT_DATA_MUX (.A ({LargeWindowShifted[16],
               AdderBoothResult[15],AdderBoothResult[14],AdderBoothResult[13],
               AdderBoothResult[12],AdderBoothResult[11],AdderBoothResult[10],
               AdderBoothResult[9],AdderBoothResult[8],AdderBoothResult[7],
               AdderBoothResult[6],AdderBoothResult[5],AdderBoothResult[4],
               AdderBoothResult[3],AdderBoothResult[2],AdderBoothResult[1],
               AdderBoothResult[0]}), .B ({LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16]}), .C ({
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],Window[7],Window[6]
               ,Window[5],Window[4],Window[3],Window[2],Window[1],Window[0],
               LargeWindowShifted[16]}), .D ({LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16],
               LargeWindowShifted[16],LargeWindowShifted[16]}), .S ({Start,Instr
               }), .Dout ({RegisterPDin_16,RegisterPDin_15,RegisterPDin_14,
               RegisterPDin_13,RegisterPDin_12,RegisterPDin_11,RegisterPDin_10,
               RegisterPDin_9,RegisterPDin_8,RegisterPDin_7,RegisterPDin_6,
               RegisterPDin_5,RegisterPDin_4,RegisterPDin_3,RegisterPDin_2,
               RegisterPDin_1,RegisterPDin_0})) ;
    fake_gnd ix43 (.Y (LargeWindowShifted[16])) ;
    dff REGISTER_A_reg_Dout_9 (.Q (BoothAddingOperand[9]), .QB (\$dummy [0]), .D (
        nx209), .CLK (CLK)) ;
    ao32 ix210 (.Y (nx209), .A0 (nx324), .A1 (Filter[0]), .A2 (Start), .B0 (
         BoothAddingOperand[9]), .B1 (nx326)) ;
    inv01 ix225 (.Y (nx224), .A (RST)) ;
    nor02_2x ix227 (.Y (nx226), .A0 (Start), .A1 (RST)) ;
    or02 ix287 (.Y (RegisterPEN), .A0 (Start), .A1 (LoopingAndResultNotReady)) ;
    mux21_ni ix46 (.Y (BoothAddingOperand[10]), .A0 (RegisterSDout_10), .A1 (
             RegisterADout_10), .S0 (nx320)) ;
    dff REGISTER_S_reg_Dout_10 (.Q (RegisterSDout_10), .QB (\$dummy [1]), .D (
        nx69), .CLK (CLK)) ;
    mux21_ni ix70 (.Y (nx69), .A0 (nx20), .A1 (RegisterSDout_10), .S0 (nx326)) ;
    aoi21 ix21 (.Y (nx20), .A0 (Filter[1]), .A1 (Filter[0]), .B0 (nx235)) ;
    or02 ix236 (.Y (nx235), .A0 (RST), .A1 (nx12)) ;
    nor02_2x ix13 (.Y (nx12), .A0 (Filter[0]), .A1 (Filter[1])) ;
    dff REGISTER_A_reg_Dout_10 (.Q (RegisterADout_10), .QB (\$dummy [2]), .D (
        nx79), .CLK (CLK)) ;
    ao32 ix80 (.Y (nx79), .A0 (nx324), .A1 (Filter[1]), .A2 (Start), .B0 (
         RegisterADout_10), .B1 (nx326)) ;
    mux21_ni ix85 (.Y (BoothAddingOperand[11]), .A0 (RegisterSDout_11), .A1 (
             RegisterADout_11), .S0 (nx320)) ;
    dff REGISTER_S_reg_Dout_11 (.Q (RegisterSDout_11), .QB (\$dummy [3]), .D (
        nx89), .CLK (CLK)) ;
    mux21_ni ix90 (.Y (nx89), .A0 (nx60), .A1 (RegisterSDout_11), .S0 (nx326)) ;
    nor03_2x ix61 (.Y (nx60), .A0 (nx249), .A1 (RST), .A2 (nx52)) ;
    nor02ii ix250 (.Y (nx249), .A0 (nx12), .A1 (Filter[2])) ;
    nor03_2x ix53 (.Y (nx52), .A0 (Filter[2]), .A1 (Filter[0]), .A2 (Filter[1])
             ) ;
    dff REGISTER_A_reg_Dout_11 (.Q (RegisterADout_11), .QB (\$dummy [4]), .D (
        nx99), .CLK (CLK)) ;
    ao32 ix100 (.Y (nx99), .A0 (nx324), .A1 (Filter[2]), .A2 (Start), .B0 (
         RegisterADout_11), .B1 (nx326)) ;
    mux21_ni ix125 (.Y (BoothAddingOperand[12]), .A0 (RegisterSDout_12), .A1 (
             RegisterADout_12), .S0 (nx320)) ;
    dff REGISTER_S_reg_Dout_12 (.Q (RegisterSDout_12), .QB (\$dummy [5]), .D (
        nx109), .CLK (CLK)) ;
    mux21_ni ix110 (.Y (nx109), .A0 (nx100), .A1 (RegisterSDout_12), .S0 (nx326)
             ) ;
    nor03_2x ix101 (.Y (nx100), .A0 (nx261), .A1 (RST), .A2 (nx92)) ;
    nor02ii ix262 (.Y (nx261), .A0 (nx52), .A1 (Filter[3])) ;
    nor04 ix93 (.Y (nx92), .A0 (Filter[3]), .A1 (Filter[2]), .A2 (Filter[0]), .A3 (
          Filter[1])) ;
    dff REGISTER_A_reg_Dout_12 (.Q (RegisterADout_12), .QB (\$dummy [6]), .D (
        nx119), .CLK (CLK)) ;
    ao32 ix120 (.Y (nx119), .A0 (nx324), .A1 (Filter[3]), .A2 (Start), .B0 (
         RegisterADout_12), .B1 (nx326)) ;
    mux21_ni ix165 (.Y (BoothAddingOperand[13]), .A0 (RegisterSDout_13), .A1 (
             RegisterADout_13), .S0 (nx320)) ;
    dff REGISTER_S_reg_Dout_13 (.Q (RegisterSDout_13), .QB (\$dummy [7]), .D (
        nx129), .CLK (CLK)) ;
    mux21_ni ix130 (.Y (nx129), .A0 (nx140), .A1 (RegisterSDout_13), .S0 (nx328)
             ) ;
    nor03_2x ix141 (.Y (nx140), .A0 (nx273), .A1 (RST), .A2 (nx132)) ;
    nor02ii ix274 (.Y (nx273), .A0 (nx92), .A1 (Filter[4])) ;
    nor02ii ix133 (.Y (nx132), .A0 (Filter[4]), .A1 (nx92)) ;
    dff REGISTER_A_reg_Dout_13 (.Q (RegisterADout_13), .QB (\$dummy [8]), .D (
        nx139), .CLK (CLK)) ;
    ao32 ix140 (.Y (nx139), .A0 (nx324), .A1 (Filter[4]), .A2 (Start), .B0 (
         RegisterADout_13), .B1 (nx328)) ;
    mux21_ni ix205 (.Y (BoothAddingOperand[14]), .A0 (RegisterSDout_14), .A1 (
             RegisterADout_14), .S0 (nx320)) ;
    dff REGISTER_S_reg_Dout_14 (.Q (RegisterSDout_14), .QB (\$dummy [9]), .D (
        nx149), .CLK (CLK)) ;
    mux21_ni ix150 (.Y (nx149), .A0 (nx180), .A1 (RegisterSDout_14), .S0 (nx328)
             ) ;
    nor03_2x ix181 (.Y (nx180), .A0 (nx286), .A1 (RST), .A2 (nx172)) ;
    nor02ii ix288 (.Y (nx286), .A0 (nx132), .A1 (Filter[5])) ;
    nor02ii ix173 (.Y (nx172), .A0 (Filter[5]), .A1 (nx132)) ;
    dff REGISTER_A_reg_Dout_14 (.Q (RegisterADout_14), .QB (\$dummy [10]), .D (
        nx159), .CLK (CLK)) ;
    ao32 ix160 (.Y (nx159), .A0 (nx324), .A1 (Filter[5]), .A2 (Start), .B0 (
         RegisterADout_14), .B1 (nx328)) ;
    mux21_ni ix245 (.Y (BoothAddingOperand[15]), .A0 (RegisterSDout_15), .A1 (
             RegisterADout_15), .S0 (nx320)) ;
    dff REGISTER_S_reg_Dout_15 (.Q (RegisterSDout_15), .QB (\$dummy [11]), .D (
        nx169), .CLK (CLK)) ;
    mux21_ni ix170 (.Y (nx169), .A0 (nx220), .A1 (RegisterSDout_15), .S0 (nx328)
             ) ;
    nor03_2x ix221 (.Y (nx220), .A0 (nx299), .A1 (RST), .A2 (nx212)) ;
    nor02ii ix300 (.Y (nx299), .A0 (nx172), .A1 (Filter[6])) ;
    nor02ii ix213 (.Y (nx212), .A0 (Filter[6]), .A1 (nx172)) ;
    dff REGISTER_A_reg_Dout_15 (.Q (RegisterADout_15), .QB (\$dummy [12]), .D (
        nx179), .CLK (CLK)) ;
    ao32 ix180 (.Y (nx179), .A0 (nx324), .A1 (Filter[6]), .A2 (Start), .B0 (
         RegisterADout_15), .B1 (nx328)) ;
    mux21_ni ix275 (.Y (BoothAddingOperand[16]), .A0 (RegisterSDout_16), .A1 (
             RegisterADout_16), .S0 (nx320)) ;
    dff REGISTER_S_reg_Dout_16 (.Q (RegisterSDout_16), .QB (\$dummy [13]), .D (
        nx189), .CLK (CLK)) ;
    ao32 ix190 (.Y (nx189), .A0 (nx224), .A1 (nx246), .A2 (Start), .B0 (
         RegisterSDout_16), .B1 (nx328)) ;
    xnor2 ix247 (.Y (nx246), .A0 (Filter[7]), .A1 (nx212)) ;
    dff REGISTER_A_reg_Dout_16 (.Q (RegisterADout_16), .QB (\$dummy [14]), .D (
        nx199), .CLK (CLK)) ;
    ao32 ix200 (.Y (nx199), .A0 (nx224), .A1 (Filter[7]), .A2 (Start), .B0 (
         RegisterADout_16), .B1 (nx226)) ;
    xor2 ix289 (.Y (BoothXORCheck), .A0 (BoothP[1]), .A1 (nx322)) ;
    buf02 ix319 (.Y (nx320), .A (BoothP[0])) ;
    buf02 ix321 (.Y (nx322), .A (BoothP[0])) ;
    inv01 ix323 (.Y (nx324), .A (RST)) ;
    nor02_2x ix325 (.Y (nx326), .A0 (Start), .A1 (RST)) ;
    nor02_2x ix327 (.Y (nx328), .A0 (Start), .A1 (RST)) ;
endmodule


module mux_4x1_17 ( A, B, C, D, S, Dout ) ;

    input [16:0]A ;
    input [16:0]B ;
    input [16:0]C ;
    input [16:0]D ;
    input [1:0]S ;
    output [16:0]Dout ;

    wire nx28, nx46, nx131, nx136, nx139, nx142, nx145, nx148, nx151, nx166, 
         nx168, nx170, nx172, nx178, nx180;



    fake_gnd ix85 (.Y (Dout[16])) ;
    ao22 ix37 (.Y (Dout[0]), .A0 (A[0]), .A1 (nx170), .B0 (C[1]), .B1 (nx166)) ;
    and02 ix29 (.Y (nx28), .A0 (S[0]), .A1 (S[1])) ;
    inv01 ix53 (.Y (Dout[1]), .A (nx131)) ;
    aoi222 ix132 (.Y (nx131), .A0 (A[1]), .A1 (nx170), .B0 (C[1]), .B1 (nx178), 
           .C0 (C[2]), .C1 (nx166)) ;
    inv01 ix65 (.Y (Dout[2]), .A (nx136)) ;
    aoi222 ix137 (.Y (nx136), .A0 (A[2]), .A1 (nx170), .B0 (C[2]), .B1 (nx178), 
           .C0 (C[3]), .C1 (nx166)) ;
    inv01 ix77 (.Y (Dout[3]), .A (nx139)) ;
    aoi222 ix140 (.Y (nx139), .A0 (A[3]), .A1 (nx170), .B0 (C[3]), .B1 (nx178), 
           .C0 (C[4]), .C1 (nx166)) ;
    inv01 ix89 (.Y (Dout[4]), .A (nx142)) ;
    aoi222 ix143 (.Y (nx142), .A0 (A[4]), .A1 (nx170), .B0 (C[4]), .B1 (nx178), 
           .C0 (C[5]), .C1 (nx166)) ;
    inv01 ix101 (.Y (Dout[5]), .A (nx145)) ;
    aoi222 ix146 (.Y (nx145), .A0 (A[5]), .A1 (nx170), .B0 (C[5]), .B1 (nx178), 
           .C0 (C[6]), .C1 (nx166)) ;
    inv01 ix113 (.Y (Dout[6]), .A (nx148)) ;
    aoi222 ix149 (.Y (nx148), .A0 (A[6]), .A1 (nx172), .B0 (C[6]), .B1 (nx178), 
           .C0 (C[7]), .C1 (nx166)) ;
    inv01 ix125 (.Y (Dout[7]), .A (nx151)) ;
    aoi222 ix152 (.Y (nx151), .A0 (A[7]), .A1 (nx172), .B0 (C[7]), .B1 (nx178), 
           .C0 (C[8]), .C1 (nx168)) ;
    ao22 ix133 (.Y (Dout[8]), .A0 (nx172), .A1 (A[8]), .B0 (C[8]), .B1 (nx180)
         ) ;
    nor02ii ix3 (.Y (Dout[9]), .A0 (S[1]), .A1 (A[9])) ;
    nor02ii ix7 (.Y (Dout[10]), .A0 (S[1]), .A1 (A[10])) ;
    nor02ii ix11 (.Y (Dout[11]), .A0 (S[1]), .A1 (A[11])) ;
    nor02ii ix15 (.Y (Dout[12]), .A0 (S[1]), .A1 (A[12])) ;
    nor02ii ix19 (.Y (Dout[13]), .A0 (S[1]), .A1 (A[13])) ;
    nor02ii ix23 (.Y (Dout[14]), .A0 (S[1]), .A1 (A[14])) ;
    nor02ii ix27 (.Y (Dout[15]), .A0 (S[1]), .A1 (A[15])) ;
    buf02 ix165 (.Y (nx166), .A (nx28)) ;
    buf02 ix167 (.Y (nx168), .A (nx28)) ;
    inv02 ix169 (.Y (nx170), .A (S[1])) ;
    inv02 ix171 (.Y (nx172), .A (S[1])) ;
    nor02ii ix47 (.Y (nx46), .A0 (S[0]), .A1 (S[1])) ;
    buf02 ix177 (.Y (nx178), .A (nx46)) ;
    buf02 ix179 (.Y (nx180), .A (nx46)) ;
endmodule


module register_edge_rising_17 ( CLK, RST, EN, Din, Dout ) ;

    input CLK ;
    input RST ;
    input EN ;
    input [16:0]Din ;
    output [16:0]Dout ;

    wire nx402, nx412, nx422, nx432, nx442, nx452, nx462, nx472, nx482, nx492, 
         nx502, nx512, nx522, nx532, nx542, nx552, nx562, nx574, nx576, nx632, 
         nx634, nx636, nx638, nx644, nx646, nx648, nx650;
    wire [16:0] \$dummy ;




    dff reg_Dout_0 (.Q (Dout[0]), .QB (\$dummy [0]), .D (nx402), .CLK (CLK)) ;
    ao32 ix403 (.Y (nx402), .A0 (Din[0]), .A1 (nx632), .A2 (nx646), .B0 (Dout[0]
         ), .B1 (nx636)) ;
    inv01 ix575 (.Y (nx574), .A (RST)) ;
    nor02_2x ix577 (.Y (nx576), .A0 (RST), .A1 (nx646)) ;
    dff reg_Dout_1 (.Q (Dout[1]), .QB (\$dummy [1]), .D (nx412), .CLK (CLK)) ;
    ao32 ix413 (.Y (nx412), .A0 (Din[1]), .A1 (nx632), .A2 (nx646), .B0 (Dout[1]
         ), .B1 (nx636)) ;
    dff reg_Dout_2 (.Q (Dout[2]), .QB (\$dummy [2]), .D (nx422), .CLK (CLK)) ;
    ao32 ix423 (.Y (nx422), .A0 (Din[2]), .A1 (nx632), .A2 (nx646), .B0 (Dout[2]
         ), .B1 (nx636)) ;
    dff reg_Dout_3 (.Q (Dout[3]), .QB (\$dummy [3]), .D (nx432), .CLK (CLK)) ;
    ao32 ix433 (.Y (nx432), .A0 (Din[3]), .A1 (nx632), .A2 (nx646), .B0 (Dout[3]
         ), .B1 (nx636)) ;
    dff reg_Dout_4 (.Q (Dout[4]), .QB (\$dummy [4]), .D (nx442), .CLK (CLK)) ;
    ao32 ix443 (.Y (nx442), .A0 (Din[4]), .A1 (nx632), .A2 (nx646), .B0 (Dout[4]
         ), .B1 (nx636)) ;
    dff reg_Dout_5 (.Q (Dout[5]), .QB (\$dummy [5]), .D (nx452), .CLK (CLK)) ;
    ao32 ix453 (.Y (nx452), .A0 (Din[5]), .A1 (nx632), .A2 (nx646), .B0 (Dout[5]
         ), .B1 (nx636)) ;
    dff reg_Dout_6 (.Q (Dout[6]), .QB (\$dummy [6]), .D (nx462), .CLK (CLK)) ;
    ao32 ix463 (.Y (nx462), .A0 (Din[6]), .A1 (nx634), .A2 (nx648), .B0 (Dout[6]
         ), .B1 (nx636)) ;
    dff reg_Dout_7 (.Q (Dout[7]), .QB (\$dummy [7]), .D (nx472), .CLK (CLK)) ;
    ao32 ix473 (.Y (nx472), .A0 (Din[7]), .A1 (nx634), .A2 (nx648), .B0 (Dout[7]
         ), .B1 (nx638)) ;
    dff reg_Dout_8 (.Q (Dout[8]), .QB (\$dummy [8]), .D (nx482), .CLK (CLK)) ;
    ao32 ix483 (.Y (nx482), .A0 (Din[8]), .A1 (nx634), .A2 (nx648), .B0 (Dout[8]
         ), .B1 (nx638)) ;
    dff reg_Dout_9 (.Q (Dout[9]), .QB (\$dummy [9]), .D (nx492), .CLK (CLK)) ;
    ao32 ix493 (.Y (nx492), .A0 (Din[9]), .A1 (nx634), .A2 (nx648), .B0 (Dout[9]
         ), .B1 (nx638)) ;
    dff reg_Dout_10 (.Q (Dout[10]), .QB (\$dummy [10]), .D (nx502), .CLK (CLK)
        ) ;
    ao32 ix503 (.Y (nx502), .A0 (Din[10]), .A1 (nx634), .A2 (nx648), .B0 (
         Dout[10]), .B1 (nx638)) ;
    dff reg_Dout_11 (.Q (Dout[11]), .QB (\$dummy [11]), .D (nx512), .CLK (CLK)
        ) ;
    ao32 ix513 (.Y (nx512), .A0 (Din[11]), .A1 (nx634), .A2 (nx648), .B0 (
         Dout[11]), .B1 (nx638)) ;
    dff reg_Dout_12 (.Q (Dout[12]), .QB (\$dummy [12]), .D (nx522), .CLK (CLK)
        ) ;
    ao32 ix523 (.Y (nx522), .A0 (Din[12]), .A1 (nx574), .A2 (nx648), .B0 (
         Dout[12]), .B1 (nx638)) ;
    dff reg_Dout_13 (.Q (Dout[13]), .QB (\$dummy [13]), .D (nx532), .CLK (CLK)
        ) ;
    ao32 ix533 (.Y (nx532), .A0 (Din[13]), .A1 (nx574), .A2 (nx650), .B0 (
         Dout[13]), .B1 (nx638)) ;
    dff reg_Dout_14 (.Q (Dout[14]), .QB (\$dummy [14]), .D (nx542), .CLK (CLK)
        ) ;
    ao32 ix543 (.Y (nx542), .A0 (Din[14]), .A1 (nx574), .A2 (nx650), .B0 (
         Dout[14]), .B1 (nx576)) ;
    dff reg_Dout_15 (.Q (Dout[15]), .QB (\$dummy [15]), .D (nx552), .CLK (CLK)
        ) ;
    ao32 ix553 (.Y (nx552), .A0 (Din[15]), .A1 (nx574), .A2 (nx650), .B0 (
         Dout[15]), .B1 (nx576)) ;
    dff reg_Dout_16 (.Q (Dout[16]), .QB (\$dummy [16]), .D (nx562), .CLK (CLK)
        ) ;
    ao32 ix563 (.Y (nx562), .A0 (Din[16]), .A1 (nx574), .A2 (nx650), .B0 (
         Dout[16]), .B1 (nx576)) ;
    inv01 ix631 (.Y (nx632), .A (RST)) ;
    inv01 ix633 (.Y (nx634), .A (RST)) ;
    nor02_2x ix635 (.Y (nx636), .A0 (RST), .A1 (nx650)) ;
    nor02_2x ix637 (.Y (nx638), .A0 (RST), .A1 (nx650)) ;
    inv01 ix643 (.Y (nx644), .A (EN)) ;
    inv02 ix645 (.Y (nx646), .A (nx644)) ;
    inv02 ix647 (.Y (nx648), .A (nx644)) ;
    inv02 ix649 (.Y (nx650), .A (nx644)) ;
endmodule


module booth_adder_17 ( AdderFirstOperand, AdderSecondOperand, BoothOperand, 
                        BoothP, SelOperand, Operation, AdderResult, 
                        AdderBoothResult ) ;

    input [16:0]AdderFirstOperand ;
    input [16:0]AdderSecondOperand ;
    input [16:0]BoothOperand ;
    input [16:0]BoothP ;
    input SelOperand ;
    input Operation ;
    output [16:0]AdderResult ;
    output [16:0]AdderBoothResult ;

    wire FirstOperand_16, FirstOperand_15, FirstOperand_14, FirstOperand_13, 
         FirstOperand_12, FirstOperand_11, FirstOperand_10, FirstOperand_9, 
         FirstOperand_8, FirstOperand_7, FirstOperand_6, FirstOperand_5, 
         FirstOperand_4, FirstOperand_3, FirstOperand_2, FirstOperand_1, 
         FirstOperand_0, SecondOperand_16, SecondOperand_15, SecondOperand_14, 
         SecondOperand_13, SecondOperand_12, SecondOperand_11, SecondOperand_10, 
         SecondOperand_9, SecondOperand_8, SecondOperand_7, SecondOperand_6, 
         SecondOperand_5, SecondOperand_4, SecondOperand_3, SecondOperand_2, 
         SecondOperand_1, SecondOperand_0, nx224, nx227, nx229, nx231, nx233, 
         nx235, nx237, nx239, nx241, nx243;
    wire [0:0] \$dummy ;




    adder_17 ADDER (.A ({FirstOperand_16,FirstOperand_15,FirstOperand_14,
             FirstOperand_13,FirstOperand_12,FirstOperand_11,FirstOperand_10,
             FirstOperand_9,FirstOperand_8,FirstOperand_7,FirstOperand_6,
             FirstOperand_5,FirstOperand_4,FirstOperand_3,FirstOperand_2,
             FirstOperand_1,FirstOperand_0}), .B ({SecondOperand_16,
             SecondOperand_15,SecondOperand_14,SecondOperand_13,SecondOperand_12
             ,SecondOperand_11,SecondOperand_10,SecondOperand_9,SecondOperand_8,
             SecondOperand_7,SecondOperand_6,SecondOperand_5,SecondOperand_4,
             SecondOperand_3,SecondOperand_2,SecondOperand_1,SecondOperand_0}), 
             .Cin (AdderBoothResult[16]), .Sum ({AdderResult[16],AdderResult[15]
             ,AdderResult[14],AdderResult[13],AdderResult[12],AdderResult[11],
             AdderResult[10],AdderResult[9],AdderResult[8],AdderResult[7],
             AdderResult[6],AdderResult[5],AdderResult[4],AdderResult[3],
             AdderResult[2],AdderResult[1],AdderResult[0]}), .Cout (\$dummy [0])
             ) ;
    fake_gnd ix47 (.Y (AdderBoothResult[16])) ;
    mux21_ni ix137 (.Y (SecondOperand_0), .A0 (AdderSecondOperand[0]), .A1 (
             BoothP[0]), .S0 (nx235)) ;
    mux21_ni ix145 (.Y (SecondOperand_1), .A0 (AdderSecondOperand[1]), .A1 (
             BoothP[1]), .S0 (nx235)) ;
    mux21_ni ix153 (.Y (SecondOperand_2), .A0 (AdderSecondOperand[2]), .A1 (
             BoothP[2]), .S0 (nx235)) ;
    mux21_ni ix161 (.Y (SecondOperand_3), .A0 (AdderSecondOperand[3]), .A1 (
             BoothP[3]), .S0 (nx235)) ;
    mux21_ni ix169 (.Y (SecondOperand_4), .A0 (AdderSecondOperand[4]), .A1 (
             BoothP[4]), .S0 (nx235)) ;
    mux21_ni ix177 (.Y (SecondOperand_5), .A0 (AdderSecondOperand[5]), .A1 (
             BoothP[5]), .S0 (nx235)) ;
    mux21_ni ix185 (.Y (SecondOperand_6), .A0 (AdderSecondOperand[6]), .A1 (
             BoothP[6]), .S0 (nx235)) ;
    mux21_ni ix193 (.Y (SecondOperand_7), .A0 (AdderSecondOperand[7]), .A1 (
             BoothP[7]), .S0 (nx237)) ;
    mux21_ni ix201 (.Y (SecondOperand_8), .A0 (AdderSecondOperand[8]), .A1 (
             BoothP[8]), .S0 (nx237)) ;
    mux21_ni ix209 (.Y (SecondOperand_9), .A0 (AdderSecondOperand[9]), .A1 (
             BoothP[9]), .S0 (nx237)) ;
    mux21_ni ix217 (.Y (SecondOperand_10), .A0 (AdderSecondOperand[10]), .A1 (
             BoothP[10]), .S0 (nx237)) ;
    mux21_ni ix225 (.Y (SecondOperand_11), .A0 (AdderSecondOperand[11]), .A1 (
             BoothP[11]), .S0 (nx237)) ;
    mux21_ni ix233 (.Y (SecondOperand_12), .A0 (AdderSecondOperand[12]), .A1 (
             BoothP[12]), .S0 (nx237)) ;
    mux21_ni ix241 (.Y (SecondOperand_13), .A0 (AdderSecondOperand[13]), .A1 (
             BoothP[13]), .S0 (nx237)) ;
    mux21_ni ix249 (.Y (SecondOperand_14), .A0 (AdderSecondOperand[14]), .A1 (
             BoothP[14]), .S0 (nx239)) ;
    mux21_ni ix257 (.Y (SecondOperand_15), .A0 (AdderSecondOperand[15]), .A1 (
             BoothP[15]), .S0 (nx239)) ;
    nor02ii ix261 (.Y (FirstOperand_0), .A0 (nx239), .A1 (AdderFirstOperand[0])
            ) ;
    nor02ii ix265 (.Y (FirstOperand_1), .A0 (nx239), .A1 (AdderFirstOperand[1])
            ) ;
    nor02ii ix269 (.Y (FirstOperand_2), .A0 (nx239), .A1 (AdderFirstOperand[2])
            ) ;
    nor02ii ix273 (.Y (FirstOperand_3), .A0 (nx239), .A1 (AdderFirstOperand[3])
            ) ;
    nor02ii ix277 (.Y (FirstOperand_4), .A0 (nx239), .A1 (AdderFirstOperand[4])
            ) ;
    nor02ii ix281 (.Y (FirstOperand_5), .A0 (nx241), .A1 (AdderFirstOperand[5])
            ) ;
    nor02ii ix285 (.Y (FirstOperand_6), .A0 (nx241), .A1 (AdderFirstOperand[6])
            ) ;
    nor02ii ix289 (.Y (FirstOperand_7), .A0 (nx241), .A1 (AdderFirstOperand[7])
            ) ;
    nor02ii ix293 (.Y (FirstOperand_8), .A0 (nx241), .A1 (AdderFirstOperand[8])
            ) ;
    mux21_ni ix303 (.Y (FirstOperand_9), .A0 (AdderFirstOperand[9]), .A1 (
             BoothOperand[9]), .S0 (nx241)) ;
    mux21_ni ix311 (.Y (FirstOperand_10), .A0 (AdderFirstOperand[10]), .A1 (
             BoothOperand[10]), .S0 (nx241)) ;
    mux21_ni ix319 (.Y (FirstOperand_11), .A0 (AdderFirstOperand[11]), .A1 (
             BoothOperand[11]), .S0 (nx241)) ;
    mux21_ni ix327 (.Y (FirstOperand_12), .A0 (AdderFirstOperand[12]), .A1 (
             BoothOperand[12]), .S0 (nx243)) ;
    mux21_ni ix335 (.Y (FirstOperand_13), .A0 (AdderFirstOperand[13]), .A1 (
             BoothOperand[13]), .S0 (nx243)) ;
    mux21_ni ix343 (.Y (FirstOperand_14), .A0 (AdderFirstOperand[14]), .A1 (
             BoothOperand[14]), .S0 (nx243)) ;
    mux21_ni ix351 (.Y (FirstOperand_15), .A0 (AdderFirstOperand[15]), .A1 (
             BoothOperand[15]), .S0 (nx243)) ;
    mux21_ni ix7 (.Y (AdderBoothResult[0]), .A0 (BoothP[1]), .A1 (AdderResult[1]
             ), .S0 (nx227)) ;
    mux21_ni ix15 (.Y (AdderBoothResult[1]), .A0 (BoothP[2]), .A1 (
             AdderResult[2]), .S0 (nx227)) ;
    mux21_ni ix23 (.Y (AdderBoothResult[2]), .A0 (BoothP[3]), .A1 (
             AdderResult[3]), .S0 (nx227)) ;
    mux21_ni ix31 (.Y (AdderBoothResult[3]), .A0 (BoothP[4]), .A1 (
             AdderResult[4]), .S0 (nx227)) ;
    mux21_ni ix39 (.Y (AdderBoothResult[4]), .A0 (BoothP[5]), .A1 (
             AdderResult[5]), .S0 (nx227)) ;
    mux21_ni ix49 (.Y (AdderBoothResult[5]), .A0 (BoothP[6]), .A1 (
             AdderResult[6]), .S0 (nx227)) ;
    mux21_ni ix55 (.Y (AdderBoothResult[6]), .A0 (BoothP[7]), .A1 (
             AdderResult[7]), .S0 (nx227)) ;
    mux21_ni ix63 (.Y (AdderBoothResult[7]), .A0 (BoothP[8]), .A1 (
             AdderResult[8]), .S0 (nx229)) ;
    mux21_ni ix71 (.Y (AdderBoothResult[8]), .A0 (BoothP[9]), .A1 (
             AdderResult[9]), .S0 (nx229)) ;
    mux21_ni ix79 (.Y (AdderBoothResult[9]), .A0 (BoothP[10]), .A1 (
             AdderResult[10]), .S0 (nx229)) ;
    mux21_ni ix87 (.Y (AdderBoothResult[10]), .A0 (BoothP[11]), .A1 (
             AdderResult[11]), .S0 (nx229)) ;
    mux21_ni ix95 (.Y (AdderBoothResult[11]), .A0 (BoothP[12]), .A1 (
             AdderResult[12]), .S0 (nx229)) ;
    mux21_ni ix103 (.Y (AdderBoothResult[12]), .A0 (BoothP[13]), .A1 (
             AdderResult[13]), .S0 (nx229)) ;
    mux21_ni ix111 (.Y (AdderBoothResult[13]), .A0 (BoothP[14]), .A1 (
             AdderResult[14]), .S0 (nx229)) ;
    mux21_ni ix119 (.Y (AdderBoothResult[14]), .A0 (BoothP[15]), .A1 (
             AdderResult[15]), .S0 (nx231)) ;
    mux21_ni ix127 (.Y (AdderBoothResult[15]), .A0 (BoothP[16]), .A1 (
             AdderResult[16]), .S0 (nx231)) ;
    and02 ix129 (.Y (SecondOperand_16), .A0 (nx243), .A1 (BoothP[16])) ;
    and02 ix295 (.Y (FirstOperand_16), .A0 (nx243), .A1 (BoothOperand[16])) ;
    inv01 ix223 (.Y (nx224), .A (Operation)) ;
    inv02 ix226 (.Y (nx227), .A (nx224)) ;
    inv02 ix228 (.Y (nx229), .A (nx224)) ;
    inv02 ix230 (.Y (nx231), .A (nx224)) ;
    inv01 ix232 (.Y (nx233), .A (SelOperand)) ;
    inv02 ix234 (.Y (nx235), .A (nx233)) ;
    inv02 ix236 (.Y (nx237), .A (nx233)) ;
    inv02 ix238 (.Y (nx239), .A (nx233)) ;
    inv02 ix240 (.Y (nx241), .A (nx233)) ;
    inv02 ix242 (.Y (nx243), .A (nx233)) ;
endmodule


module adder_17 ( A, B, Cin, Sum, Cout ) ;

    input [16:0]A ;
    input [16:0]B ;
    input Cin ;
    output [16:0]Sum ;
    output Cout ;

    wire nx2, nx16, nx18, nx32, nx34, nx48, nx50, nx64, nx66, nx80, nx82, nx96, 
         nx98, nx112, nx114, nx122, nx105, nx107, nx111, nx115, nx121, nx123, 
         nx127, nx131, nx137, nx139, nx143, nx147, nx153, nx155, nx159, nx163, 
         nx167, nx169, nx172, nx175, nx179, nx181, nx184, nx187, nx191, nx193, 
         nx196, nx199, nx203, nx205, nx208;



    fake_gnd ix58 (.Y (Cout)) ;
    xor2 ix161 (.Y (Sum[0]), .A0 (B[0]), .A1 (A[0])) ;
    xor2 ix155 (.Y (Sum[1]), .A0 (nx105), .A1 (nx107)) ;
    nand02 ix106 (.Y (nx105), .A0 (B[0]), .A1 (A[0])) ;
    xnor2 ix108 (.Y (nx107), .A0 (A[1]), .A1 (B[1])) ;
    xor2 ix153 (.Y (Sum[2]), .A0 (nx111), .A1 (nx115)) ;
    aoi32 ix112 (.Y (nx111), .A0 (B[0]), .A1 (A[0]), .A2 (nx2), .B0 (B[1]), .B1 (
          A[1])) ;
    xnor2 ix116 (.Y (nx115), .A0 (A[2]), .A1 (B[2])) ;
    xnor2 ix151 (.Y (Sum[3]), .A0 (nx16), .A1 (nx123)) ;
    oai21 ix17 (.Y (nx16), .A0 (nx111), .A1 (nx115), .B0 (nx121)) ;
    nand02 ix122 (.Y (nx121), .A0 (B[2]), .A1 (A[2])) ;
    xnor2 ix124 (.Y (nx123), .A0 (A[3]), .A1 (B[3])) ;
    xor2 ix149 (.Y (Sum[4]), .A0 (nx127), .A1 (nx131)) ;
    aoi22 ix128 (.Y (nx127), .A0 (B[3]), .A1 (A[3]), .B0 (nx16), .B1 (nx18)) ;
    xnor2 ix132 (.Y (nx131), .A0 (A[4]), .A1 (B[4])) ;
    xnor2 ix147 (.Y (Sum[5]), .A0 (nx32), .A1 (nx139)) ;
    oai21 ix33 (.Y (nx32), .A0 (nx127), .A1 (nx131), .B0 (nx137)) ;
    nand02 ix138 (.Y (nx137), .A0 (B[4]), .A1 (A[4])) ;
    xnor2 ix140 (.Y (nx139), .A0 (A[5]), .A1 (B[5])) ;
    xor2 ix145 (.Y (Sum[6]), .A0 (nx143), .A1 (nx147)) ;
    aoi22 ix144 (.Y (nx143), .A0 (B[5]), .A1 (A[5]), .B0 (nx32), .B1 (nx34)) ;
    xnor2 ix148 (.Y (nx147), .A0 (A[6]), .A1 (B[6])) ;
    xnor2 ix143 (.Y (Sum[7]), .A0 (nx48), .A1 (nx155)) ;
    oai21 ix49 (.Y (nx48), .A0 (nx143), .A1 (nx147), .B0 (nx153)) ;
    nand02 ix154 (.Y (nx153), .A0 (B[6]), .A1 (A[6])) ;
    xnor2 ix156 (.Y (nx155), .A0 (A[7]), .A1 (B[7])) ;
    xor2 ix141 (.Y (Sum[8]), .A0 (nx159), .A1 (nx163)) ;
    aoi22 ix160 (.Y (nx159), .A0 (B[7]), .A1 (A[7]), .B0 (nx48), .B1 (nx50)) ;
    xnor2 ix164 (.Y (nx163), .A0 (A[8]), .A1 (B[8])) ;
    xnor2 ix139 (.Y (Sum[9]), .A0 (nx64), .A1 (nx169)) ;
    oai21 ix65 (.Y (nx64), .A0 (nx159), .A1 (nx163), .B0 (nx167)) ;
    nand02 ix168 (.Y (nx167), .A0 (B[8]), .A1 (A[8])) ;
    xnor2 ix170 (.Y (nx169), .A0 (A[9]), .A1 (B[9])) ;
    xor2 ix137 (.Y (Sum[10]), .A0 (nx172), .A1 (nx175)) ;
    aoi22 ix173 (.Y (nx172), .A0 (B[9]), .A1 (A[9]), .B0 (nx64), .B1 (nx66)) ;
    xnor2 ix176 (.Y (nx175), .A0 (A[10]), .A1 (B[10])) ;
    xnor2 ix135 (.Y (Sum[11]), .A0 (nx80), .A1 (nx181)) ;
    oai21 ix81 (.Y (nx80), .A0 (nx172), .A1 (nx175), .B0 (nx179)) ;
    nand02 ix180 (.Y (nx179), .A0 (B[10]), .A1 (A[10])) ;
    xnor2 ix182 (.Y (nx181), .A0 (A[11]), .A1 (B[11])) ;
    xor2 ix133 (.Y (Sum[12]), .A0 (nx184), .A1 (nx187)) ;
    aoi22 ix185 (.Y (nx184), .A0 (B[11]), .A1 (A[11]), .B0 (nx80), .B1 (nx82)) ;
    xnor2 ix188 (.Y (nx187), .A0 (A[12]), .A1 (B[12])) ;
    xnor2 ix131 (.Y (Sum[13]), .A0 (nx96), .A1 (nx193)) ;
    oai21 ix97 (.Y (nx96), .A0 (nx184), .A1 (nx187), .B0 (nx191)) ;
    nand02 ix192 (.Y (nx191), .A0 (B[12]), .A1 (A[12])) ;
    xnor2 ix194 (.Y (nx193), .A0 (A[13]), .A1 (B[13])) ;
    xor2 ix129 (.Y (Sum[14]), .A0 (nx196), .A1 (nx199)) ;
    aoi22 ix197 (.Y (nx196), .A0 (B[13]), .A1 (A[13]), .B0 (nx96), .B1 (nx98)) ;
    xnor2 ix200 (.Y (nx199), .A0 (A[14]), .A1 (B[14])) ;
    xnor2 ix127 (.Y (Sum[15]), .A0 (nx112), .A1 (nx205)) ;
    oai21 ix113 (.Y (nx112), .A0 (nx196), .A1 (nx199), .B0 (nx203)) ;
    nand02 ix204 (.Y (nx203), .A0 (B[14]), .A1 (A[14])) ;
    xnor2 ix206 (.Y (nx205), .A0 (A[15]), .A1 (B[15])) ;
    xnor2 ix125 (.Y (Sum[16]), .A0 (nx208), .A1 (nx122)) ;
    aoi22 ix209 (.Y (nx208), .A0 (B[15]), .A1 (A[15]), .B0 (nx112), .B1 (nx114)
          ) ;
    xor2 ix123 (.Y (nx122), .A0 (A[16]), .A1 (B[16])) ;
    inv01 ix115 (.Y (nx114), .A (nx205)) ;
    inv01 ix99 (.Y (nx98), .A (nx193)) ;
    inv01 ix83 (.Y (nx82), .A (nx181)) ;
    inv01 ix67 (.Y (nx66), .A (nx169)) ;
    inv01 ix51 (.Y (nx50), .A (nx155)) ;
    inv01 ix35 (.Y (nx34), .A (nx139)) ;
    inv01 ix19 (.Y (nx18), .A (nx123)) ;
    inv01 ix3 (.Y (nx2), .A (nx107)) ;
endmodule


module controller ( CLK, RST, Start, FilterSize, Stride, Instr, CalcFinished, 
                    Calc, MemRD, MemWR, MemAddr, CacheFilterWR, CacheWindowWR, 
                    FirstCycle, Done ) ;

    input CLK ;
    input RST ;
    input Start ;
    input FilterSize ;
    input Stride ;
    input Instr ;
    input CalcFinished ;
    output Calc ;
    output MemRD ;
    output MemWR ;
    output [17:0]MemAddr ;
    output CacheFilterWR ;
    output CacheWindowWR ;
    output FirstCycle ;
    output Done ;

    wire CurCol_5, nx483, CurRow_5, CurRow_4, CurRow_3, CurRow_2, CurRow_0, nx14, 
         nx34, nx46, nx491, nx82, nx102, CurRow_7, CurRow_6, nx118, nx138, nx162, 
         nx164, nx178, nx188, nx196, nx226, nx232, nx248, nx266, nx278, CurCol_4, 
         CurCol_3, CurCol_2, CurCol_1, CurCol_0, nx495, nx300, nx497, nx336, 
         nx501, nx362, nx372, nx392, nx400, CurCol_7, CurCol_6, nx414, nx426, 
         nx452, nx460, nx466, nx476, nx482, nx498, nx520, nx522, nx538, nx556, 
         nx558, nx574, nx592, nx594, nx610, nx626, nx644, nx660, nx666, nx688, 
         nx694, nx716, nx513, nx523, nx533, nx543, nx553, nx563, nx573, nx583, 
         nx593, nx603, nx613, nx623, nx633, nx643, nx653, nx663, nx681, nx693, 
         nx695, nx701, nx705, nx713, nx715, nx725, nx727, nx733, nx735, nx743, 
         nx745, nx748, nx752, nx754, nx758, nx761, nx764, nx768, nx770, nx773, 
         nx777, nx779, nx783, nx785, nx792, nx796, nx798, nx801, nx805, nx807, 
         nx810, nx814, nx817, nx822, nx825, nx828, nx831, nx835, nx837, nx845, 
         nx847, nx850, nx852, nx855, nx861, nx863, nx867, nx870, nx872, nx877, 
         nx880, nx882, nx884, nx900, nx904, nx913, nx916, nx923, nx926, nx929, 
         nx931, nx934, nx938, nx941, nx944, nx948, nx952, nx955, nx958, nx962, 
         nx968, nx975, nx979, nx981, nx987, nx989, nx992, nx1002, nx1004, nx1008, 
         nx1010, nx1012, nx1014, nx1016, nx1018, nx1020, nx1022, nx1024, nx1026, 
         nx1030, nx1032, nx1034, nx1036, nx1042, nx1044, nx1046, nx1048, nx1050, 
         nx1052, nx1054, nx1056, nx1058, nx1060, nx1062, nx1064, nx1066, nx1068, 
         nx1070, nx1072;
    wire [4:0] \$dummy ;




    assign MemAddr[16] = MemWR ;
    fake_gnd ix469 (.Y (MemRD)) ;
    and03 ix279 (.Y (nx278), .A0 (nx681), .A1 (CalcFinished), .A2 (Calc)) ;
    aoi21 ix682 (.Y (nx681), .A0 (Start), .A1 (nx483), .B0 (RST)) ;
    nor03_2x ix401 (.Y (nx400), .A0 (nx693), .A1 (nx1026), .A2 (nx392)) ;
    nand02 ix696 (.Y (nx695), .A0 (CurCol_4), .A1 (nx501)) ;
    oai21 ix634 (.Y (nx633), .A0 (nx701), .A1 (nx1020), .B0 (nx904)) ;
    dff COL_reg_Dout_4 (.Q (CurCol_4), .QB (nx701), .D (nx633), .CLK (CLK)) ;
    oai21 ix706 (.Y (nx705), .A0 (CacheFilterWR), .A1 (CacheWindowWR), .B0 (
          nx882)) ;
    aoi22 ix714 (.Y (nx713), .A0 (nx715), .A1 (FirstCycle), .B0 (CacheFilterWR)
          , .B1 (nx188)) ;
    inv01 ix716 (.Y (nx715), .A (Instr)) ;
    dff STATE_reg_Dout_3 (.Q (Calc), .QB (\$dummy [0]), .D (nx266), .CLK (CLK)
        ) ;
    aoi22 ix726 (.Y (nx725), .A0 (nx727), .A1 (Calc), .B0 (CacheWindowWR), .B1 (
          nx226)) ;
    inv01 ix728 (.Y (nx727), .A (CalcFinished)) ;
    dff STATE_reg_Dout_1 (.Q (CacheWindowWR), .QB (\$dummy [1]), .D (nx248), .CLK (
        CLK)) ;
    aoi221 ix734 (.Y (nx733), .A0 (CacheFilterWR), .A1 (nx735), .B0 (nx1002), .B1 (
           nx792), .C0 (nx232)) ;
    nand04 ix736 (.Y (nx735), .A0 (nx162), .A1 (nx178), .A2 (nx752), .A3 (nx758)
           ) ;
    oai21 ix564 (.Y (nx563), .A0 (nx743), .A1 (nx1014), .B0 (nx745)) ;
    dff ROW_reg_Dout_5 (.Q (CurRow_5), .QB (nx743), .D (nx563), .CLK (CLK)) ;
    nand02 ix749 (.Y (nx748), .A0 (CurRow_4), .A1 (nx491)) ;
    oai21 ix554 (.Y (nx553), .A0 (nx752), .A1 (nx1014), .B0 (nx754)) ;
    dff ROW_reg_Dout_4 (.Q (CurRow_4), .QB (nx752), .D (nx553), .CLK (CLK)) ;
    nand04 ix755 (.Y (nx754), .A0 (nx82), .A1 (nx748), .A2 (nx1032), .A3 (nx1020
           )) ;
    or02 ix83 (.Y (nx82), .A0 (nx491), .A1 (CurRow_4)) ;
    oai21 ix544 (.Y (nx543), .A0 (nx758), .A1 (nx1014), .B0 (nx761)) ;
    oai21 ix534 (.Y (nx533), .A0 (nx768), .A1 (nx1014), .B0 (nx770)) ;
    dff ROW_reg_Dout_2 (.Q (CurRow_2), .QB (nx768), .D (nx533), .CLK (CLK)) ;
    nand04 ix771 (.Y (nx770), .A0 (nx46), .A1 (nx764), .A2 (nx1030), .A3 (nx1018
           )) ;
    nand02 ix47 (.Y (nx46), .A0 (nx773), .A1 (nx768)) ;
    dff ROW_reg_Dout_1 (.Q (\$dummy [2]), .QB (nx777), .D (nx523), .CLK (CLK)) ;
    oai21 ix780 (.Y (nx779), .A0 (CurRow_0), .A1 (nx1022), .B0 (nx34)) ;
    oai21 ix514 (.Y (nx513), .A0 (nx783), .A1 (nx1014), .B0 (nx785)) ;
    dff ROW_reg_Dout_0 (.Q (CurRow_0), .QB (nx783), .D (nx513), .CLK (CLK)) ;
    nand04 ix793 (.Y (nx792), .A0 (CurCol_5), .A1 (CurCol_7), .A2 (CurCol_6), .A3 (
           nx460)) ;
    oai21 ix664 (.Y (nx663), .A0 (nx796), .A1 (nx1014), .B0 (nx798)) ;
    dff COL_reg_Dout_7 (.Q (CurCol_7), .QB (nx796), .D (nx663), .CLK (CLK)) ;
    nand03 ix799 (.Y (nx798), .A0 (nx1030), .A1 (nx426), .A2 (nx1016)) ;
    nand02 ix802 (.Y (nx801), .A0 (CurCol_6), .A1 (nx392)) ;
    dff COL_reg_Dout_6 (.Q (CurCol_6), .QB (nx805), .D (nx653), .CLK (CLK)) ;
    oai21 ix808 (.Y (nx807), .A0 (nx392), .A1 (CurCol_6), .B0 (nx414)) ;
    dff COL_reg_Dout_5 (.Q (CurCol_5), .QB (nx810), .D (nx643), .CLK (CLK)) ;
    aoi21 ix415 (.Y (nx414), .A0 (CurCol_6), .A1 (nx392), .B0 (nx1026)) ;
    oai21 ix15 (.Y (nx14), .A0 (nx814), .A1 (nx733), .B0 (nx681)) ;
    dff STATE_reg_Dout_0 (.Q (CacheFilterWR), .QB (nx814), .D (nx196), .CLK (CLK
        )) ;
    nor03_2x ix461 (.Y (nx460), .A0 (nx817), .A1 (nx701), .A2 (nx872)) ;
    aoi32 ix818 (.Y (nx817), .A0 (CurCol_0), .A1 (FilterSize), .A2 (CurCol_1), .B0 (
          CurCol_2), .B1 (nx452)) ;
    dff COL_reg_Dout_0 (.Q (CurCol_0), .QB (nx847), .D (nx593), .CLK (CLK)) ;
    xnor2 ix823 (.Y (nx822), .A0 (nx138), .A1 (nx495)) ;
    oai21 ix584 (.Y (nx583), .A0 (nx825), .A1 (nx1016), .B0 (nx828)) ;
    nand02 ix832 (.Y (nx831), .A0 (CurRow_6), .A1 (nx102)) ;
    oai21 ix574 (.Y (nx573), .A0 (nx835), .A1 (nx1016), .B0 (nx837)) ;
    dff ROW_reg_Dout_6 (.Q (CurRow_6), .QB (nx835), .D (nx573), .CLK (CLK)) ;
    nand04 ix838 (.Y (nx837), .A0 (nx118), .A1 (nx831), .A2 (nx1030), .A3 (
           nx1016)) ;
    or02 ix119 (.Y (nx118), .A0 (nx102), .A1 (CurRow_6)) ;
    dff ROW_reg_Dout_7 (.Q (CurRow_7), .QB (nx825), .D (nx583), .CLK (CLK)) ;
    nand02 ix846 (.Y (nx845), .A0 (Stride), .A1 (nx138)) ;
    oai21 ix604 (.Y (nx603), .A0 (nx850), .A1 (nx1016), .B0 (nx852)) ;
    dff COL_reg_Dout_1 (.Q (CurCol_1), .QB (nx850), .D (nx603), .CLK (CLK)) ;
    oai21 ix856 (.Y (nx855), .A0 (CurCol_0), .A1 (Stride), .B0 (nx138)) ;
    oai21 ix614 (.Y (nx613), .A0 (nx861), .A1 (nx1018), .B0 (nx863)) ;
    dff COL_reg_Dout_2 (.Q (CurCol_2), .QB (nx861), .D (nx613), .CLK (CLK)) ;
    nand04 ix864 (.Y (nx863), .A0 (nx336), .A1 (nx1030), .A2 (nx867), .A3 (
           nx1018)) ;
    or02 ix337 (.Y (nx336), .A0 (nx497), .A1 (CurCol_2)) ;
    nand02 ix868 (.Y (nx867), .A0 (CurCol_2), .A1 (nx497)) ;
    inv01 ix871 (.Y (nx870), .A (FilterSize)) ;
    dff COL_reg_Dout_3 (.Q (CurCol_3), .QB (nx872), .D (nx623), .CLK (CLK)) ;
    nor03_2x ix363 (.Y (nx362), .A0 (nx877), .A1 (nx1026), .A2 (nx501)) ;
    aoi22 ix881 (.Y (nx880), .A0 (Instr), .A1 (FirstCycle), .B0 (CacheWindowWR)
          , .B1 (nx882)) ;
    oai21 ix883 (.Y (nx882), .A0 (nx783), .A1 (nx884), .B0 (nx735)) ;
    inv01 ix885 (.Y (nx884), .A (Stride)) ;
    aoi21 ix35 (.Y (nx34), .A0 (nx1022), .A1 (CurRow_0), .B0 (nx1026)) ;
    dff ROW_reg_Dout_3 (.Q (CurRow_3), .QB (nx758), .D (nx543), .CLK (CLK)) ;
    aoi21 ix179 (.Y (nx178), .A0 (nx870), .A1 (nx1022), .B0 (CurRow_2)) ;
    dff STATE_reg_Dout_2 (.Q (MemWR), .QB (\$dummy [3]), .D (nx278), .CLK (CLK)
        ) ;
    nand04 ix905 (.Y (nx904), .A0 (nx372), .A1 (nx1032), .A2 (nx695), .A3 (
           nx1020)) ;
    or02 ix373 (.Y (nx372), .A0 (nx501), .A1 (CurCol_4)) ;
    dff STATE_reg_Dout_4 (.Q (Done), .QB (\$dummy [4]), .D (nx466), .CLK (CLK)
        ) ;
    nor03_2x ix470 (.Y (nx466), .A0 (nx792), .A1 (Start), .A2 (RST)) ;
    oai21 ix495 (.Y (MemAddr[0]), .A0 (nx847), .A1 (nx1034), .B0 (nx913)) ;
    aoi32 ix914 (.Y (nx913), .A0 (nx482), .A1 (nx1002), .A2 (nx916), .B0 (
          CurRow_0), .B1 (nx1008)) ;
    nand02 ix483 (.Y (nx482), .A0 (nx847), .A1 (FilterSize)) ;
    xor2 ix499 (.Y (nx498), .A0 (nx916), .A1 (nx923)) ;
    oai21 ix535 (.Y (MemAddr[2]), .A0 (nx861), .A1 (nx1034), .B0 (nx926)) ;
    aoi32 ix927 (.Y (nx926), .A0 (nx520), .A1 (nx1002), .A2 (nx931), .B0 (
          CurRow_2), .B1 (nx1008)) ;
    nand02 ix521 (.Y (nx520), .A0 (nx929), .A1 (nx861)) ;
    oai21 ix930 (.Y (nx929), .A0 (FilterSize), .A1 (CurCol_0), .B0 (CurCol_1)) ;
    oai21 ix553 (.Y (MemAddr[3]), .A0 (nx872), .A1 (nx1034), .B0 (nx934)) ;
    aoi32 ix935 (.Y (nx934), .A0 (nx538), .A1 (nx1002), .A2 (nx938), .B0 (
          CurRow_3), .B1 (nx1008)) ;
    or02 ix539 (.Y (nx538), .A0 (nx522), .A1 (CurCol_3)) ;
    nand02 ix939 (.Y (nx938), .A0 (CurCol_3), .A1 (nx522)) ;
    oai21 ix571 (.Y (MemAddr[4]), .A0 (nx701), .A1 (nx1034), .B0 (nx941)) ;
    aoi32 ix942 (.Y (nx941), .A0 (nx556), .A1 (nx1004), .A2 (nx944), .B0 (
          CurRow_4), .B1 (nx1008)) ;
    nand02 ix557 (.Y (nx556), .A0 (nx938), .A1 (nx701)) ;
    oai21 ix589 (.Y (MemAddr[5]), .A0 (nx810), .A1 (nx1034), .B0 (nx948)) ;
    aoi32 ix949 (.Y (nx948), .A0 (nx574), .A1 (nx1004), .A2 (nx952), .B0 (
          CurRow_5), .B1 (nx1008)) ;
    or02 ix575 (.Y (nx574), .A0 (nx558), .A1 (CurCol_5)) ;
    nand02 ix953 (.Y (nx952), .A0 (CurCol_5), .A1 (nx558)) ;
    oai21 ix607 (.Y (MemAddr[6]), .A0 (nx805), .A1 (nx1034), .B0 (nx955)) ;
    aoi32 ix956 (.Y (nx955), .A0 (nx592), .A1 (nx1004), .A2 (nx958), .B0 (
          CurRow_6), .B1 (nx1010)) ;
    nand02 ix593 (.Y (nx592), .A0 (nx952), .A1 (nx805)) ;
    oai21 ix623 (.Y (MemAddr[7]), .A0 (nx796), .A1 (nx1034), .B0 (nx962)) ;
    aoi32 ix963 (.Y (nx962), .A0 (nx610), .A1 (nx884), .A2 (nx1004), .B0 (
          CurRow_7), .B1 (nx1010)) ;
    ao32 ix641 (.Y (MemAddr[8]), .A0 (nx626), .A1 (CurRow_0), .A2 (nx900), .B0 (
         nx1004), .B1 (nx968)) ;
    xnor2 ix645 (.Y (nx644), .A0 (nx968), .A1 (nx164)) ;
    oai21 ix667 (.Y (nx666), .A0 (nx768), .A1 (nx975), .B0 (nx660)) ;
    aoi21 ix976 (.Y (nx975), .A0 (CurRow_0), .A1 (nx870), .B0 (nx1024)) ;
    nand02 ix661 (.Y (nx660), .A0 (nx975), .A1 (nx768)) ;
    oai22 ix687 (.Y (MemAddr[11]), .A0 (nx1066), .A1 (nx979), .B0 (nx758), .B1 (
          nx1036)) ;
    aoi21 ix980 (.Y (nx979), .A0 (CurRow_3), .A1 (nx660), .B0 (nx981)) ;
    oai21 ix695 (.Y (nx694), .A0 (nx752), .A1 (nx981), .B0 (nx688)) ;
    nand02 ix689 (.Y (nx688), .A0 (nx981), .A1 (nx752)) ;
    oai22 ix715 (.Y (MemAddr[13]), .A0 (nx1066), .A1 (nx987), .B0 (nx743), .B1 (
          nx1036)) ;
    aoi21 ix988 (.Y (nx987), .A0 (CurRow_5), .A1 (nx688), .B0 (nx989)) ;
    oai22 ix729 (.Y (MemAddr[14]), .A0 (nx1066), .A1 (nx992), .B0 (nx835), .B1 (
          nx1036)) ;
    nand02 ix717 (.Y (nx716), .A0 (nx989), .A1 (nx835)) ;
    inv01 ix959 (.Y (nx958), .A (nx594)) ;
    inv01 ix945 (.Y (nx944), .A (nx558)) ;
    inv01 ix932 (.Y (nx931), .A (nx522)) ;
    inv01 ix233 (.Y (nx232), .A (nx880)) ;
    inv01 ix227 (.Y (nx226), .A (nx882)) ;
    inv01 ix189 (.Y (nx188), .A (nx735)) ;
    inv01 ix463 (.Y (nx483), .A (nx792)) ;
    inv01 ix901 (.Y (nx900), .A (MemAddr[17])) ;
    inv02 ix1001 (.Y (nx1002), .A (nx1066)) ;
    inv02 ix1003 (.Y (nx1004), .A (nx1066)) ;
    inv01 ix1007 (.Y (nx1008), .A (nx900)) ;
    inv01 ix1009 (.Y (nx1010), .A (nx900)) ;
    inv02 ix1013 (.Y (nx1014), .A (nx1012)) ;
    inv02 ix1015 (.Y (nx1016), .A (nx1070)) ;
    inv02 ix1017 (.Y (nx1018), .A (nx1070)) ;
    inv02 ix1019 (.Y (nx1020), .A (nx1070)) ;
    inv02 ix1021 (.Y (nx1022), .A (nx777)) ;
    inv02 ix1023 (.Y (nx1024), .A (nx777)) ;
    inv02 ix1025 (.Y (nx1026), .A (nx1032)) ;
    inv02 ix1029 (.Y (nx1030), .A (nx14)) ;
    inv02 ix1031 (.Y (nx1032), .A (nx1064)) ;
    inv02 ix1033 (.Y (nx1034), .A (nx476)) ;
    inv02 ix1035 (.Y (nx1036), .A (nx476)) ;
    nor02ii ix209 (.Y (MemAddr[17]), .A0 (CacheWindowWR), .A1 (nx1066)) ;
    mux21_ni ix644 (.Y (nx643), .A0 (nx400), .A1 (CurCol_5), .S0 (nx1070)) ;
    and02 ix694 (.Y (nx693), .A0 (nx810), .A1 (nx695)) ;
    nor03_2x ix295 (.Y (nx1012), .A0 (nx1042), .A1 (nx1064), .A2 (MemWR)) ;
    inv01 ix1041 (.Y (nx1042), .A (nx705)) ;
    nor02ii ix197 (.Y (nx196), .A0 (nx713), .A1 (nx681)) ;
    and04 ix215 (.Y (FirstCycle), .A0 (Start), .A1 (nx1044), .A2 (nx814), .A3 (
          MemAddr[17])) ;
    inv01 ix1043 (.Y (nx1044), .A (Calc)) ;
    nor02ii ix267 (.Y (nx266), .A0 (nx725), .A1 (nx681)) ;
    nor02ii ix249 (.Y (nx248), .A0 (nx733), .A1 (nx681)) ;
    and03 ix163 (.Y (nx162), .A0 (nx743), .A1 (nx825), .A2 (nx835)) ;
    or04 ix746 (.Y (nx745), .A0 (nx1046), .A1 (nx102), .A2 (nx1064), .A3 (nx1070
         )) ;
    nor02ii ix101 (.Y (nx1046), .A0 (CurRow_5), .A1 (nx748)) ;
    nor02ii ix81 (.Y (nx491), .A0 (nx764), .A1 (CurRow_3)) ;
    or04 ix762 (.Y (nx761), .A0 (nx1048), .A1 (nx491), .A2 (nx1064), .A3 (nx1070
         )) ;
    nor02ii ix65 (.Y (nx1048), .A0 (CurRow_3), .A1 (nx764)) ;
    or03 ix765 (.Y (nx764), .A0 (nx768), .A1 (nx777), .A2 (nx783)) ;
    or02 ix774 (.Y (nx773), .A0 (nx777), .A1 (nx783)) ;
    mux21 ix524 (.Y (nx523), .A0 (nx779), .A1 (nx777), .S0 (nx1070)) ;
    or03 ix786 (.Y (nx785), .A0 (CurRow_0), .A1 (nx1064), .A2 (nx1072)) ;
    xor2 ix427 (.Y (nx426), .A0 (nx796), .A1 (nx801)) ;
    mux21 ix654 (.Y (nx653), .A0 (nx807), .A1 (nx805), .S0 (nx1072)) ;
    nor02ii ix393 (.Y (nx392), .A0 (nx695), .A1 (CurCol_5)) ;
    mux21_ni ix594 (.Y (nx593), .A0 (nx300), .A1 (CurCol_0), .S0 (nx1072)) ;
    nor02ii ix301 (.Y (nx300), .A0 (nx822), .A1 (nx1032)) ;
    nor02ii ix139 (.Y (nx138), .A0 (nx831), .A1 (CurRow_7)) ;
    or04 ix829 (.Y (nx828), .A0 (nx1050), .A1 (nx1064), .A2 (nx138), .A3 (nx1072
         )) ;
    nor02ii ix137 (.Y (nx1050), .A0 (CurRow_7), .A1 (nx831)) ;
    nor02ii ix103 (.Y (nx102), .A0 (nx748), .A1 (CurRow_5)) ;
    xor2 ix311 (.Y (nx495), .A0 (nx847), .A1 (nx845)) ;
    or04 ix853 (.Y (nx852), .A0 (nx1052), .A1 (nx1064), .A2 (nx497), .A3 (nx1072
         )) ;
    nor02ii ix319 (.Y (nx1052), .A0 (CurCol_1), .A1 (nx855)) ;
    nor02ii ix335 (.Y (nx497), .A0 (nx855), .A1 (CurCol_1)) ;
    or03 ix453 (.Y (nx452), .A0 (CurCol_1), .A1 (FilterSize), .A2 (CurCol_0)) ;
    mux21_ni ix624 (.Y (nx623), .A0 (nx362), .A1 (CurCol_3), .S0 (nx1072)) ;
    and02 ix878 (.Y (nx877), .A0 (nx872), .A1 (nx867)) ;
    nor02ii ix371 (.Y (nx501), .A0 (nx867), .A1 (CurCol_3)) ;
    or02 ix917 (.Y (nx916), .A0 (FilterSize), .A1 (nx847)) ;
    oai222 ix920 (.Y (MemAddr[1]), .A0 (nx1066), .A1 (nx1054), .B0 (nx850), .B1 (
           nx1036), .C0 (nx777), .C1 (nx900)) ;
    inv01 ix1053 (.Y (nx1054), .A (nx498)) ;
    and02 ix477 (.Y (nx476), .A0 (nx1068), .A1 (CacheWindowWR)) ;
    xor2 ix924 (.Y (nx923), .A0 (FilterSize), .A1 (nx850)) ;
    nor02ii ix523 (.Y (nx522), .A0 (nx929), .A1 (CurCol_2)) ;
    nor02ii ix559 (.Y (nx558), .A0 (nx938), .A1 (CurCol_4)) ;
    xor2 ix611 (.Y (nx610), .A0 (nx594), .A1 (CurCol_7)) ;
    nor02ii ix595 (.Y (nx594), .A0 (nx952), .A1 (CurCol_6)) ;
    or02 ix627 (.Y (nx626), .A0 (nx1068), .A1 (FilterSize)) ;
    nor02ii ix969 (.Y (nx968), .A0 (FilterSize), .A1 (nx783)) ;
    oai22 ix649 (.Y (MemAddr[9]), .A0 (nx1068), .A1 (nx1056), .B0 (nx777), .B1 (
          nx1036)) ;
    inv01 ix1055 (.Y (nx1056), .A (nx644)) ;
    xor2 ix165 (.Y (nx164), .A0 (FilterSize), .A1 (nx777)) ;
    oai22 ix673 (.Y (MemAddr[10]), .A0 (nx1068), .A1 (nx1058), .B0 (nx768), .B1 (
          nx1036)) ;
    inv01 ix1057 (.Y (nx1058), .A (nx666)) ;
    nor02ii ix982 (.Y (nx981), .A0 (nx660), .A1 (nx758)) ;
    oai22 ix701 (.Y (MemAddr[12]), .A0 (nx1068), .A1 (nx1060), .B0 (nx752), .B1 (
          nx1036)) ;
    inv01 ix1059 (.Y (nx1060), .A (nx694)) ;
    nor02ii ix990 (.Y (nx989), .A0 (nx688), .A1 (nx743)) ;
    xor2 ix993 (.Y (nx992), .A0 (nx835), .A1 (nx989)) ;
    oai32 ix741 (.Y (MemAddr[15]), .A0 (nx1062), .A1 (Stride), .A2 (nx1068), .B0 (
          nx825), .B1 (nx1036)) ;
    xnor2 ix731 (.Y (nx1062), .A0 (nx825), .A1 (nx716)) ;
    inv02 ix1063 (.Y (nx1064), .A (nx1030)) ;
    inv02 ix1065 (.Y (nx1066), .A (MemWR)) ;
    inv02 ix1067 (.Y (nx1068), .A (MemWR)) ;
    inv02 ix1069 (.Y (nx1070), .A (nx1014)) ;
    inv02 ix1071 (.Y (nx1072), .A (nx1014)) ;
endmodule

